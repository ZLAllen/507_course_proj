
module memory_WIDTH8_SIZE9_LOGSIZE4 ( clk, data_in, data_out, addr, wr_en );
  input [7:0] data_in;
  output [7:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] ,
         \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] ,
         \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] ,
         \mem[6][0] , \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] ,
         \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] ,
         \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] ,
         \mem[4][1] , \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] ,
         \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] ,
         \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] ,
         \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] ,
         \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] ,
         \mem[1][0] , N40, N41, N42, N43, N44, N45, N46, N47, n1, n2, n3, n4,
         n5, n6, n7, n8, n65, n66, n67, n68, n69, n70, n71, n72, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93;

  DFF_X1 \mem_reg[8][7]  ( .D(n216), .CK(clk), .QN(n1) );
  DFF_X1 \mem_reg[8][6]  ( .D(n215), .CK(clk), .QN(n2) );
  DFF_X1 \mem_reg[8][5]  ( .D(n214), .CK(clk), .QN(n3) );
  DFF_X1 \mem_reg[8][4]  ( .D(n213), .CK(clk), .QN(n4) );
  DFF_X1 \mem_reg[8][3]  ( .D(n212), .CK(clk), .QN(n5) );
  DFF_X1 \mem_reg[8][2]  ( .D(n211), .CK(clk), .QN(n6) );
  DFF_X1 \mem_reg[8][1]  ( .D(n210), .CK(clk), .QN(n7) );
  DFF_X1 \mem_reg[8][0]  ( .D(n209), .CK(clk), .QN(n8) );
  DFF_X1 \mem_reg[7][7]  ( .D(n9), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n10), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n11), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n12), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n13), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n14), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n15), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n16), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n17), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n18), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n19), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n20), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n21), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n22), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n23), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n24), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n25), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n26), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n27), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n28), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n29), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n30), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n31), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n32), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n33), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n34), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n35), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n36), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n37), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n38), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n39), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n40), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n41), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n42), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n43), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n44), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n45), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n46), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n47), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n48), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n49), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n50), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n51), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n52), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n53), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n54), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n55), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n56), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n57), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n58), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n59), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n60), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n61), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n62), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n63), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n64), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n208), .CK(clk), .QN(n65) );
  DFF_X1 \data_out_reg[7]  ( .D(N40), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n207), .CK(clk), .QN(n66) );
  DFF_X1 \data_out_reg[6]  ( .D(N41), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n206), .CK(clk), .QN(n67) );
  DFF_X1 \data_out_reg[5]  ( .D(N42), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n205), .CK(clk), .QN(n68) );
  DFF_X1 \data_out_reg[4]  ( .D(N43), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n204), .CK(clk), .QN(n69) );
  DFF_X1 \data_out_reg[3]  ( .D(N44), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n203), .CK(clk), .QN(n70) );
  DFF_X1 \data_out_reg[2]  ( .D(N45), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n202), .CK(clk), .QN(n71) );
  DFF_X1 \data_out_reg[1]  ( .D(N46), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n201), .CK(clk), .QN(n72) );
  DFF_X1 \data_out_reg[0]  ( .D(N47), .CK(clk), .Q(data_out[0]) );
  NAND3_X1 U202 ( .A1(n169), .A2(n170), .A3(n171), .ZN(N47) );
  NAND3_X1 U203 ( .A1(n173), .A2(n174), .A3(n175), .ZN(N46) );
  NAND3_X1 U204 ( .A1(n177), .A2(n178), .A3(n179), .ZN(N45) );
  NAND3_X1 U205 ( .A1(n181), .A2(n182), .A3(n183), .ZN(N44) );
  NAND3_X1 U206 ( .A1(n185), .A2(n186), .A3(n187), .ZN(N43) );
  NAND3_X1 U207 ( .A1(n189), .A2(n190), .A3(n191), .ZN(N42) );
  NAND3_X1 U208 ( .A1(n193), .A2(n194), .A3(n195), .ZN(N41) );
  NAND3_X1 U209 ( .A1(n197), .A2(n198), .A3(n199), .ZN(N40) );
  NAND3_X1 U210 ( .A1(n91), .A2(n93), .A3(n168), .ZN(n95) );
  NOR2_X1 U3 ( .A1(n81), .A2(addr[3]), .ZN(n106) );
  INV_X1 U4 ( .A(n94), .ZN(n73) );
  NOR2_X1 U5 ( .A1(n81), .A2(n95), .ZN(n94) );
  INV_X1 U6 ( .A(n118), .ZN(n78) );
  INV_X1 U7 ( .A(n108), .ZN(n79) );
  INV_X1 U8 ( .A(n97), .ZN(n80) );
  INV_X1 U9 ( .A(n128), .ZN(n77) );
  INV_X1 U10 ( .A(n138), .ZN(n76) );
  INV_X1 U11 ( .A(n148), .ZN(n75) );
  INV_X1 U12 ( .A(n158), .ZN(n74) );
  INV_X1 U13 ( .A(wr_en), .ZN(n81) );
  NAND2_X1 U14 ( .A1(n105), .A2(n106), .ZN(n97) );
  NAND2_X1 U15 ( .A1(n116), .A2(n106), .ZN(n108) );
  NAND2_X1 U16 ( .A1(n126), .A2(n106), .ZN(n118) );
  NAND2_X1 U17 ( .A1(n136), .A2(n106), .ZN(n128) );
  NAND2_X1 U18 ( .A1(n146), .A2(n106), .ZN(n138) );
  NAND2_X1 U19 ( .A1(n156), .A2(n106), .ZN(n148) );
  NAND2_X1 U20 ( .A1(n166), .A2(n106), .ZN(n158) );
  INV_X1 U21 ( .A(n167), .ZN(n82) );
  NOR3_X2 U22 ( .A1(n91), .A2(addr[2]), .A3(n92), .ZN(n126) );
  NOR3_X2 U23 ( .A1(addr[0]), .A2(addr[2]), .A3(n92), .ZN(n116) );
  AND3_X1 U24 ( .A1(n91), .A2(n92), .A3(addr[2]), .ZN(n136) );
  AND3_X1 U25 ( .A1(addr[1]), .A2(addr[0]), .A3(addr[2]), .ZN(n166) );
  AND3_X1 U26 ( .A1(addr[1]), .A2(n91), .A3(addr[2]), .ZN(n156) );
  AND3_X1 U27 ( .A1(addr[0]), .A2(n92), .A3(addr[2]), .ZN(n146) );
  OAI22_X1 U28 ( .A1(n93), .A2(n8), .B1(n95), .B2(n72), .ZN(n172) );
  OAI22_X1 U29 ( .A1(n93), .A2(n7), .B1(n95), .B2(n71), .ZN(n176) );
  OAI22_X1 U30 ( .A1(n93), .A2(n6), .B1(n95), .B2(n70), .ZN(n180) );
  OAI22_X1 U31 ( .A1(n93), .A2(n5), .B1(n95), .B2(n69), .ZN(n184) );
  OAI22_X1 U32 ( .A1(n93), .A2(n4), .B1(n95), .B2(n68), .ZN(n188) );
  OAI22_X1 U33 ( .A1(n93), .A2(n3), .B1(n95), .B2(n67), .ZN(n192) );
  OAI22_X1 U34 ( .A1(n93), .A2(n2), .B1(n95), .B2(n66), .ZN(n196) );
  OAI22_X1 U35 ( .A1(n93), .A2(n1), .B1(n95), .B2(n65), .ZN(n200) );
  NAND4_X1 U36 ( .A1(addr[3]), .A2(wr_en), .A3(n168), .A4(n91), .ZN(n167) );
  INV_X1 U37 ( .A(addr[3]), .ZN(n93) );
  NOR2_X1 U38 ( .A1(addr[1]), .A2(addr[2]), .ZN(n168) );
  OAI22_X1 U39 ( .A1(n73), .A2(n90), .B1(n94), .B2(n72), .ZN(n201) );
  OAI22_X1 U40 ( .A1(n73), .A2(n89), .B1(n94), .B2(n71), .ZN(n202) );
  OAI22_X1 U41 ( .A1(n73), .A2(n88), .B1(n94), .B2(n70), .ZN(n203) );
  OAI22_X1 U42 ( .A1(n73), .A2(n87), .B1(n94), .B2(n69), .ZN(n204) );
  OAI22_X1 U43 ( .A1(n73), .A2(n86), .B1(n94), .B2(n68), .ZN(n205) );
  OAI22_X1 U44 ( .A1(n73), .A2(n85), .B1(n94), .B2(n67), .ZN(n206) );
  OAI22_X1 U45 ( .A1(n73), .A2(n84), .B1(n94), .B2(n66), .ZN(n207) );
  OAI22_X1 U46 ( .A1(n73), .A2(n83), .B1(n94), .B2(n65), .ZN(n208) );
  INV_X1 U47 ( .A(addr[0]), .ZN(n91) );
  OAI22_X1 U48 ( .A1(n90), .A2(n167), .B1(n82), .B2(n8), .ZN(n209) );
  OAI22_X1 U49 ( .A1(n89), .A2(n167), .B1(n82), .B2(n7), .ZN(n210) );
  OAI22_X1 U50 ( .A1(n88), .A2(n167), .B1(n82), .B2(n6), .ZN(n211) );
  OAI22_X1 U51 ( .A1(n87), .A2(n167), .B1(n82), .B2(n5), .ZN(n212) );
  OAI22_X1 U52 ( .A1(n86), .A2(n167), .B1(n82), .B2(n4), .ZN(n213) );
  OAI22_X1 U53 ( .A1(n85), .A2(n167), .B1(n82), .B2(n3), .ZN(n214) );
  OAI22_X1 U54 ( .A1(n84), .A2(n167), .B1(n82), .B2(n2), .ZN(n215) );
  OAI22_X1 U55 ( .A1(n83), .A2(n167), .B1(n82), .B2(n1), .ZN(n216) );
  AND2_X1 U56 ( .A1(addr[0]), .A2(n168), .ZN(n105) );
  INV_X1 U57 ( .A(addr[1]), .ZN(n92) );
  AOI22_X1 U58 ( .A1(\mem[4][0] ), .A2(n136), .B1(\mem[3][0] ), .B2(n126), 
        .ZN(n169) );
  AOI222_X1 U59 ( .A1(\mem[5][0] ), .A2(n146), .B1(\mem[7][0] ), .B2(n166), 
        .C1(\mem[6][0] ), .C2(n156), .ZN(n170) );
  AOI221_X1 U60 ( .B1(\mem[2][0] ), .B2(n116), .C1(\mem[1][0] ), .C2(n105), 
        .A(n172), .ZN(n171) );
  AOI22_X1 U61 ( .A1(\mem[4][1] ), .A2(n136), .B1(\mem[3][1] ), .B2(n126), 
        .ZN(n173) );
  AOI222_X1 U62 ( .A1(\mem[5][1] ), .A2(n146), .B1(\mem[7][1] ), .B2(n166), 
        .C1(\mem[6][1] ), .C2(n156), .ZN(n174) );
  AOI221_X1 U63 ( .B1(\mem[2][1] ), .B2(n116), .C1(\mem[1][1] ), .C2(n105), 
        .A(n176), .ZN(n175) );
  AOI22_X1 U64 ( .A1(\mem[4][2] ), .A2(n136), .B1(\mem[3][2] ), .B2(n126), 
        .ZN(n177) );
  AOI222_X1 U65 ( .A1(\mem[5][2] ), .A2(n146), .B1(\mem[7][2] ), .B2(n166), 
        .C1(\mem[6][2] ), .C2(n156), .ZN(n178) );
  AOI221_X1 U66 ( .B1(\mem[2][2] ), .B2(n116), .C1(\mem[1][2] ), .C2(n105), 
        .A(n180), .ZN(n179) );
  AOI22_X1 U67 ( .A1(\mem[4][3] ), .A2(n136), .B1(\mem[3][3] ), .B2(n126), 
        .ZN(n181) );
  AOI222_X1 U68 ( .A1(\mem[5][3] ), .A2(n146), .B1(\mem[7][3] ), .B2(n166), 
        .C1(\mem[6][3] ), .C2(n156), .ZN(n182) );
  AOI221_X1 U69 ( .B1(\mem[2][3] ), .B2(n116), .C1(\mem[1][3] ), .C2(n105), 
        .A(n184), .ZN(n183) );
  AOI22_X1 U70 ( .A1(\mem[4][4] ), .A2(n136), .B1(\mem[3][4] ), .B2(n126), 
        .ZN(n185) );
  AOI222_X1 U71 ( .A1(\mem[5][4] ), .A2(n146), .B1(\mem[7][4] ), .B2(n166), 
        .C1(\mem[6][4] ), .C2(n156), .ZN(n186) );
  AOI221_X1 U72 ( .B1(\mem[2][4] ), .B2(n116), .C1(\mem[1][4] ), .C2(n105), 
        .A(n188), .ZN(n187) );
  AOI22_X1 U73 ( .A1(\mem[4][5] ), .A2(n136), .B1(\mem[3][5] ), .B2(n126), 
        .ZN(n189) );
  AOI222_X1 U74 ( .A1(\mem[5][5] ), .A2(n146), .B1(\mem[7][5] ), .B2(n166), 
        .C1(\mem[6][5] ), .C2(n156), .ZN(n190) );
  AOI221_X1 U75 ( .B1(\mem[2][5] ), .B2(n116), .C1(\mem[1][5] ), .C2(n105), 
        .A(n192), .ZN(n191) );
  AOI22_X1 U76 ( .A1(\mem[4][6] ), .A2(n136), .B1(\mem[3][6] ), .B2(n126), 
        .ZN(n193) );
  AOI222_X1 U77 ( .A1(\mem[5][6] ), .A2(n146), .B1(\mem[7][6] ), .B2(n166), 
        .C1(\mem[6][6] ), .C2(n156), .ZN(n194) );
  AOI221_X1 U78 ( .B1(\mem[2][6] ), .B2(n116), .C1(\mem[1][6] ), .C2(n105), 
        .A(n196), .ZN(n195) );
  AOI22_X1 U79 ( .A1(\mem[4][7] ), .A2(n136), .B1(\mem[3][7] ), .B2(n126), 
        .ZN(n197) );
  AOI222_X1 U80 ( .A1(\mem[5][7] ), .A2(n146), .B1(\mem[7][7] ), .B2(n166), 
        .C1(\mem[6][7] ), .C2(n156), .ZN(n198) );
  AOI221_X1 U81 ( .B1(\mem[2][7] ), .B2(n116), .C1(\mem[1][7] ), .C2(n105), 
        .A(n200), .ZN(n199) );
  INV_X1 U82 ( .A(data_in[0]), .ZN(n90) );
  INV_X1 U83 ( .A(data_in[1]), .ZN(n89) );
  INV_X1 U84 ( .A(data_in[2]), .ZN(n88) );
  INV_X1 U85 ( .A(data_in[3]), .ZN(n87) );
  INV_X1 U86 ( .A(data_in[4]), .ZN(n86) );
  INV_X1 U87 ( .A(data_in[5]), .ZN(n85) );
  INV_X1 U88 ( .A(data_in[6]), .ZN(n84) );
  INV_X1 U89 ( .A(data_in[7]), .ZN(n83) );
  INV_X1 U90 ( .A(n96), .ZN(n64) );
  AOI22_X1 U91 ( .A1(data_in[0]), .A2(n80), .B1(n97), .B2(\mem[1][0] ), .ZN(
        n96) );
  INV_X1 U92 ( .A(n98), .ZN(n63) );
  AOI22_X1 U93 ( .A1(data_in[1]), .A2(n80), .B1(n97), .B2(\mem[1][1] ), .ZN(
        n98) );
  INV_X1 U94 ( .A(n99), .ZN(n62) );
  AOI22_X1 U95 ( .A1(data_in[2]), .A2(n80), .B1(n97), .B2(\mem[1][2] ), .ZN(
        n99) );
  INV_X1 U96 ( .A(n100), .ZN(n61) );
  AOI22_X1 U97 ( .A1(data_in[3]), .A2(n80), .B1(n97), .B2(\mem[1][3] ), .ZN(
        n100) );
  INV_X1 U98 ( .A(n101), .ZN(n60) );
  AOI22_X1 U99 ( .A1(data_in[4]), .A2(n80), .B1(n97), .B2(\mem[1][4] ), .ZN(
        n101) );
  INV_X1 U100 ( .A(n102), .ZN(n59) );
  AOI22_X1 U101 ( .A1(data_in[5]), .A2(n80), .B1(n97), .B2(\mem[1][5] ), .ZN(
        n102) );
  INV_X1 U102 ( .A(n103), .ZN(n58) );
  AOI22_X1 U103 ( .A1(data_in[6]), .A2(n80), .B1(n97), .B2(\mem[1][6] ), .ZN(
        n103) );
  INV_X1 U104 ( .A(n104), .ZN(n57) );
  AOI22_X1 U105 ( .A1(data_in[7]), .A2(n80), .B1(n97), .B2(\mem[1][7] ), .ZN(
        n104) );
  INV_X1 U106 ( .A(n107), .ZN(n56) );
  AOI22_X1 U107 ( .A1(data_in[0]), .A2(n79), .B1(n108), .B2(\mem[2][0] ), .ZN(
        n107) );
  INV_X1 U108 ( .A(n109), .ZN(n55) );
  AOI22_X1 U109 ( .A1(data_in[1]), .A2(n79), .B1(n108), .B2(\mem[2][1] ), .ZN(
        n109) );
  INV_X1 U110 ( .A(n110), .ZN(n54) );
  AOI22_X1 U111 ( .A1(data_in[2]), .A2(n79), .B1(n108), .B2(\mem[2][2] ), .ZN(
        n110) );
  INV_X1 U112 ( .A(n111), .ZN(n53) );
  AOI22_X1 U113 ( .A1(data_in[3]), .A2(n79), .B1(n108), .B2(\mem[2][3] ), .ZN(
        n111) );
  INV_X1 U114 ( .A(n112), .ZN(n52) );
  AOI22_X1 U115 ( .A1(data_in[4]), .A2(n79), .B1(n108), .B2(\mem[2][4] ), .ZN(
        n112) );
  INV_X1 U116 ( .A(n113), .ZN(n51) );
  AOI22_X1 U117 ( .A1(data_in[5]), .A2(n79), .B1(n108), .B2(\mem[2][5] ), .ZN(
        n113) );
  INV_X1 U118 ( .A(n114), .ZN(n50) );
  AOI22_X1 U119 ( .A1(data_in[6]), .A2(n79), .B1(n108), .B2(\mem[2][6] ), .ZN(
        n114) );
  INV_X1 U120 ( .A(n115), .ZN(n49) );
  AOI22_X1 U121 ( .A1(data_in[7]), .A2(n79), .B1(n108), .B2(\mem[2][7] ), .ZN(
        n115) );
  INV_X1 U122 ( .A(n117), .ZN(n48) );
  AOI22_X1 U123 ( .A1(data_in[0]), .A2(n78), .B1(n118), .B2(\mem[3][0] ), .ZN(
        n117) );
  INV_X1 U124 ( .A(n119), .ZN(n47) );
  AOI22_X1 U125 ( .A1(data_in[1]), .A2(n78), .B1(n118), .B2(\mem[3][1] ), .ZN(
        n119) );
  INV_X1 U126 ( .A(n120), .ZN(n46) );
  AOI22_X1 U127 ( .A1(data_in[2]), .A2(n78), .B1(n118), .B2(\mem[3][2] ), .ZN(
        n120) );
  INV_X1 U128 ( .A(n121), .ZN(n45) );
  AOI22_X1 U129 ( .A1(data_in[3]), .A2(n78), .B1(n118), .B2(\mem[3][3] ), .ZN(
        n121) );
  INV_X1 U130 ( .A(n122), .ZN(n44) );
  AOI22_X1 U131 ( .A1(data_in[4]), .A2(n78), .B1(n118), .B2(\mem[3][4] ), .ZN(
        n122) );
  INV_X1 U132 ( .A(n123), .ZN(n43) );
  AOI22_X1 U133 ( .A1(data_in[5]), .A2(n78), .B1(n118), .B2(\mem[3][5] ), .ZN(
        n123) );
  INV_X1 U134 ( .A(n124), .ZN(n42) );
  AOI22_X1 U135 ( .A1(data_in[6]), .A2(n78), .B1(n118), .B2(\mem[3][6] ), .ZN(
        n124) );
  INV_X1 U136 ( .A(n125), .ZN(n41) );
  AOI22_X1 U137 ( .A1(data_in[7]), .A2(n78), .B1(n118), .B2(\mem[3][7] ), .ZN(
        n125) );
  INV_X1 U138 ( .A(n127), .ZN(n40) );
  AOI22_X1 U139 ( .A1(data_in[0]), .A2(n77), .B1(n128), .B2(\mem[4][0] ), .ZN(
        n127) );
  INV_X1 U140 ( .A(n129), .ZN(n39) );
  AOI22_X1 U141 ( .A1(data_in[1]), .A2(n77), .B1(n128), .B2(\mem[4][1] ), .ZN(
        n129) );
  INV_X1 U142 ( .A(n130), .ZN(n38) );
  AOI22_X1 U143 ( .A1(data_in[2]), .A2(n77), .B1(n128), .B2(\mem[4][2] ), .ZN(
        n130) );
  INV_X1 U144 ( .A(n131), .ZN(n37) );
  AOI22_X1 U145 ( .A1(data_in[3]), .A2(n77), .B1(n128), .B2(\mem[4][3] ), .ZN(
        n131) );
  INV_X1 U146 ( .A(n132), .ZN(n36) );
  AOI22_X1 U147 ( .A1(data_in[4]), .A2(n77), .B1(n128), .B2(\mem[4][4] ), .ZN(
        n132) );
  INV_X1 U148 ( .A(n133), .ZN(n35) );
  AOI22_X1 U149 ( .A1(data_in[5]), .A2(n77), .B1(n128), .B2(\mem[4][5] ), .ZN(
        n133) );
  INV_X1 U150 ( .A(n134), .ZN(n34) );
  AOI22_X1 U151 ( .A1(data_in[6]), .A2(n77), .B1(n128), .B2(\mem[4][6] ), .ZN(
        n134) );
  INV_X1 U152 ( .A(n135), .ZN(n33) );
  AOI22_X1 U153 ( .A1(data_in[7]), .A2(n77), .B1(n128), .B2(\mem[4][7] ), .ZN(
        n135) );
  INV_X1 U154 ( .A(n137), .ZN(n32) );
  AOI22_X1 U155 ( .A1(data_in[0]), .A2(n76), .B1(n138), .B2(\mem[5][0] ), .ZN(
        n137) );
  INV_X1 U156 ( .A(n139), .ZN(n31) );
  AOI22_X1 U157 ( .A1(data_in[1]), .A2(n76), .B1(n138), .B2(\mem[5][1] ), .ZN(
        n139) );
  INV_X1 U158 ( .A(n140), .ZN(n30) );
  AOI22_X1 U159 ( .A1(data_in[2]), .A2(n76), .B1(n138), .B2(\mem[5][2] ), .ZN(
        n140) );
  INV_X1 U160 ( .A(n141), .ZN(n29) );
  AOI22_X1 U161 ( .A1(data_in[3]), .A2(n76), .B1(n138), .B2(\mem[5][3] ), .ZN(
        n141) );
  INV_X1 U162 ( .A(n142), .ZN(n28) );
  AOI22_X1 U163 ( .A1(data_in[4]), .A2(n76), .B1(n138), .B2(\mem[5][4] ), .ZN(
        n142) );
  INV_X1 U164 ( .A(n143), .ZN(n27) );
  AOI22_X1 U165 ( .A1(data_in[5]), .A2(n76), .B1(n138), .B2(\mem[5][5] ), .ZN(
        n143) );
  INV_X1 U166 ( .A(n144), .ZN(n26) );
  AOI22_X1 U167 ( .A1(data_in[6]), .A2(n76), .B1(n138), .B2(\mem[5][6] ), .ZN(
        n144) );
  INV_X1 U168 ( .A(n145), .ZN(n25) );
  AOI22_X1 U169 ( .A1(data_in[7]), .A2(n76), .B1(n138), .B2(\mem[5][7] ), .ZN(
        n145) );
  INV_X1 U170 ( .A(n147), .ZN(n24) );
  AOI22_X1 U171 ( .A1(data_in[0]), .A2(n75), .B1(n148), .B2(\mem[6][0] ), .ZN(
        n147) );
  INV_X1 U172 ( .A(n149), .ZN(n23) );
  AOI22_X1 U173 ( .A1(data_in[1]), .A2(n75), .B1(n148), .B2(\mem[6][1] ), .ZN(
        n149) );
  INV_X1 U174 ( .A(n150), .ZN(n22) );
  AOI22_X1 U175 ( .A1(data_in[2]), .A2(n75), .B1(n148), .B2(\mem[6][2] ), .ZN(
        n150) );
  INV_X1 U176 ( .A(n151), .ZN(n21) );
  AOI22_X1 U177 ( .A1(data_in[3]), .A2(n75), .B1(n148), .B2(\mem[6][3] ), .ZN(
        n151) );
  INV_X1 U178 ( .A(n152), .ZN(n20) );
  AOI22_X1 U179 ( .A1(data_in[4]), .A2(n75), .B1(n148), .B2(\mem[6][4] ), .ZN(
        n152) );
  INV_X1 U180 ( .A(n153), .ZN(n19) );
  AOI22_X1 U181 ( .A1(data_in[5]), .A2(n75), .B1(n148), .B2(\mem[6][5] ), .ZN(
        n153) );
  INV_X1 U182 ( .A(n154), .ZN(n18) );
  AOI22_X1 U183 ( .A1(data_in[6]), .A2(n75), .B1(n148), .B2(\mem[6][6] ), .ZN(
        n154) );
  INV_X1 U184 ( .A(n155), .ZN(n17) );
  AOI22_X1 U185 ( .A1(data_in[7]), .A2(n75), .B1(n148), .B2(\mem[6][7] ), .ZN(
        n155) );
  INV_X1 U186 ( .A(n157), .ZN(n16) );
  AOI22_X1 U187 ( .A1(data_in[0]), .A2(n74), .B1(n158), .B2(\mem[7][0] ), .ZN(
        n157) );
  INV_X1 U188 ( .A(n159), .ZN(n15) );
  AOI22_X1 U189 ( .A1(data_in[1]), .A2(n74), .B1(n158), .B2(\mem[7][1] ), .ZN(
        n159) );
  INV_X1 U190 ( .A(n160), .ZN(n14) );
  AOI22_X1 U191 ( .A1(data_in[2]), .A2(n74), .B1(n158), .B2(\mem[7][2] ), .ZN(
        n160) );
  INV_X1 U192 ( .A(n161), .ZN(n13) );
  AOI22_X1 U193 ( .A1(data_in[3]), .A2(n74), .B1(n158), .B2(\mem[7][3] ), .ZN(
        n161) );
  INV_X1 U194 ( .A(n162), .ZN(n12) );
  AOI22_X1 U195 ( .A1(data_in[4]), .A2(n74), .B1(n158), .B2(\mem[7][4] ), .ZN(
        n162) );
  INV_X1 U196 ( .A(n163), .ZN(n11) );
  AOI22_X1 U197 ( .A1(data_in[5]), .A2(n74), .B1(n158), .B2(\mem[7][5] ), .ZN(
        n163) );
  INV_X1 U198 ( .A(n164), .ZN(n10) );
  AOI22_X1 U199 ( .A1(data_in[6]), .A2(n74), .B1(n158), .B2(\mem[7][6] ), .ZN(
        n164) );
  INV_X1 U200 ( .A(n165), .ZN(n9) );
  AOI22_X1 U201 ( .A1(data_in[7]), .A2(n74), .B1(n158), .B2(\mem[7][7] ), .ZN(
        n165) );
endmodule


module memory_WIDTH8_SIZE3_LOGSIZE2_0 ( clk, data_in, data_out, addr, wr_en );
  input [7:0] data_in;
  output [7:0] data_out;
  input [1:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, N15, N16, N17, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38;

  DFF_X1 \mem_reg[2][7]  ( .D(n66), .CK(clk), .QN(n1) );
  DFF_X1 \mem_reg[2][6]  ( .D(n65), .CK(clk), .QN(n2) );
  DFF_X1 \mem_reg[2][5]  ( .D(n64), .CK(clk), .QN(n3) );
  DFF_X1 \mem_reg[2][4]  ( .D(n63), .CK(clk), .QN(n4) );
  DFF_X1 \mem_reg[2][3]  ( .D(n62), .CK(clk), .QN(n5) );
  DFF_X1 \mem_reg[2][2]  ( .D(n61), .CK(clk), .QN(n6) );
  DFF_X1 \mem_reg[2][1]  ( .D(n60), .CK(clk), .QN(n7) );
  DFF_X1 \mem_reg[2][0]  ( .D(n59), .CK(clk), .QN(n8) );
  DFF_X1 \mem_reg[1][7]  ( .D(n58), .CK(clk), .QN(n9) );
  DFF_X1 \mem_reg[1][6]  ( .D(n57), .CK(clk), .QN(n10) );
  DFF_X1 \mem_reg[1][5]  ( .D(n56), .CK(clk), .QN(n11) );
  DFF_X1 \mem_reg[1][4]  ( .D(n55), .CK(clk), .QN(n12) );
  DFF_X1 \mem_reg[1][3]  ( .D(n54), .CK(clk), .QN(n13) );
  DFF_X1 \mem_reg[1][2]  ( .D(n53), .CK(clk), .QN(n14) );
  DFF_X1 \mem_reg[1][1]  ( .D(n52), .CK(clk), .QN(n15) );
  DFF_X1 \mem_reg[1][0]  ( .D(n51), .CK(clk), .QN(n16) );
  DFF_X1 \mem_reg[0][7]  ( .D(n50), .CK(clk), .QN(n17) );
  DFF_X1 \data_out_reg[7]  ( .D(N10), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n49), .CK(clk), .QN(n18) );
  DFF_X1 \data_out_reg[6]  ( .D(N11), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n48), .CK(clk), .QN(n19) );
  DFF_X1 \data_out_reg[5]  ( .D(N12), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n47), .CK(clk), .QN(n20) );
  DFF_X1 \data_out_reg[4]  ( .D(N13), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n46), .CK(clk), .QN(n21) );
  DFF_X1 \data_out_reg[3]  ( .D(N14), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n45), .CK(clk), .QN(n22) );
  DFF_X1 \data_out_reg[2]  ( .D(N15), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n44), .CK(clk), .QN(n23) );
  DFF_X1 \data_out_reg[1]  ( .D(N16), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n43), .CK(clk), .QN(n24) );
  DFF_X1 \data_out_reg[0]  ( .D(N17), .CK(clk), .Q(data_out[0]) );
  NOR3_X2 U20 ( .A1(n28), .A2(addr[1]), .A3(n37), .ZN(n41) );
  NOR3_X2 U29 ( .A1(n28), .A2(addr[0]), .A3(n38), .ZN(n42) );
  INV_X1 U3 ( .A(n39), .ZN(n25) );
  NOR2_X1 U4 ( .A1(n28), .A2(n40), .ZN(n39) );
  INV_X1 U5 ( .A(wr_en), .ZN(n28) );
  NAND2_X1 U6 ( .A1(n37), .A2(n38), .ZN(n40) );
  INV_X1 U7 ( .A(n41), .ZN(n26) );
  INV_X1 U8 ( .A(n42), .ZN(n27) );
  INV_X1 U9 ( .A(addr[1]), .ZN(n38) );
  INV_X1 U10 ( .A(addr[0]), .ZN(n37) );
  OAI222_X1 U11 ( .A1(n37), .A2(n16), .B1(n40), .B2(n24), .C1(n38), .C2(n8), 
        .ZN(N17) );
  OAI222_X1 U12 ( .A1(n37), .A2(n15), .B1(n40), .B2(n23), .C1(n38), .C2(n7), 
        .ZN(N16) );
  OAI222_X1 U13 ( .A1(n37), .A2(n14), .B1(n40), .B2(n22), .C1(n38), .C2(n6), 
        .ZN(N15) );
  OAI222_X1 U14 ( .A1(n37), .A2(n13), .B1(n40), .B2(n21), .C1(n38), .C2(n5), 
        .ZN(N14) );
  OAI222_X1 U15 ( .A1(n37), .A2(n12), .B1(n40), .B2(n20), .C1(n38), .C2(n4), 
        .ZN(N13) );
  OAI222_X1 U16 ( .A1(n37), .A2(n11), .B1(n40), .B2(n19), .C1(n38), .C2(n3), 
        .ZN(N12) );
  OAI222_X1 U17 ( .A1(n37), .A2(n10), .B1(n40), .B2(n18), .C1(n38), .C2(n2), 
        .ZN(N11) );
  OAI222_X1 U18 ( .A1(n37), .A2(n9), .B1(n40), .B2(n17), .C1(n38), .C2(n1), 
        .ZN(N10) );
  OAI22_X1 U19 ( .A1(n36), .A2(n27), .B1(n42), .B2(n8), .ZN(n59) );
  OAI22_X1 U21 ( .A1(n35), .A2(n27), .B1(n42), .B2(n7), .ZN(n60) );
  OAI22_X1 U22 ( .A1(n34), .A2(n27), .B1(n42), .B2(n6), .ZN(n61) );
  OAI22_X1 U23 ( .A1(n33), .A2(n27), .B1(n42), .B2(n5), .ZN(n62) );
  OAI22_X1 U24 ( .A1(n32), .A2(n27), .B1(n42), .B2(n4), .ZN(n63) );
  OAI22_X1 U25 ( .A1(n31), .A2(n27), .B1(n42), .B2(n3), .ZN(n64) );
  OAI22_X1 U26 ( .A1(n30), .A2(n27), .B1(n42), .B2(n2), .ZN(n65) );
  OAI22_X1 U27 ( .A1(n29), .A2(n27), .B1(n42), .B2(n1), .ZN(n66) );
  OAI22_X1 U28 ( .A1(n36), .A2(n26), .B1(n41), .B2(n16), .ZN(n51) );
  OAI22_X1 U30 ( .A1(n35), .A2(n26), .B1(n41), .B2(n15), .ZN(n52) );
  OAI22_X1 U31 ( .A1(n34), .A2(n26), .B1(n41), .B2(n14), .ZN(n53) );
  OAI22_X1 U32 ( .A1(n33), .A2(n26), .B1(n41), .B2(n13), .ZN(n54) );
  OAI22_X1 U33 ( .A1(n32), .A2(n26), .B1(n41), .B2(n12), .ZN(n55) );
  OAI22_X1 U34 ( .A1(n31), .A2(n26), .B1(n41), .B2(n11), .ZN(n56) );
  OAI22_X1 U35 ( .A1(n30), .A2(n26), .B1(n41), .B2(n10), .ZN(n57) );
  OAI22_X1 U36 ( .A1(n29), .A2(n26), .B1(n41), .B2(n9), .ZN(n58) );
  OAI22_X1 U37 ( .A1(n25), .A2(n36), .B1(n39), .B2(n24), .ZN(n43) );
  OAI22_X1 U38 ( .A1(n25), .A2(n35), .B1(n39), .B2(n23), .ZN(n44) );
  OAI22_X1 U39 ( .A1(n25), .A2(n34), .B1(n39), .B2(n22), .ZN(n45) );
  OAI22_X1 U40 ( .A1(n25), .A2(n33), .B1(n39), .B2(n21), .ZN(n46) );
  OAI22_X1 U41 ( .A1(n25), .A2(n32), .B1(n39), .B2(n20), .ZN(n47) );
  OAI22_X1 U42 ( .A1(n25), .A2(n31), .B1(n39), .B2(n19), .ZN(n48) );
  OAI22_X1 U43 ( .A1(n25), .A2(n30), .B1(n39), .B2(n18), .ZN(n49) );
  OAI22_X1 U44 ( .A1(n25), .A2(n29), .B1(n39), .B2(n17), .ZN(n50) );
  INV_X1 U45 ( .A(data_in[0]), .ZN(n36) );
  INV_X1 U46 ( .A(data_in[1]), .ZN(n35) );
  INV_X1 U47 ( .A(data_in[2]), .ZN(n34) );
  INV_X1 U48 ( .A(data_in[3]), .ZN(n33) );
  INV_X1 U49 ( .A(data_in[4]), .ZN(n32) );
  INV_X1 U50 ( .A(data_in[5]), .ZN(n31) );
  INV_X1 U51 ( .A(data_in[6]), .ZN(n30) );
  INV_X1 U52 ( .A(data_in[7]), .ZN(n29) );
endmodule


module memory_WIDTH8_SIZE3_LOGSIZE2_1 ( clk, data_in, data_out, addr, wr_en );
  input [7:0] data_in;
  output [7:0] data_out;
  input [1:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, N15, N16, N17, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118;

  DFF_X1 \mem_reg[2][7]  ( .D(n67), .CK(clk), .QN(n118) );
  DFF_X1 \mem_reg[2][6]  ( .D(n68), .CK(clk), .QN(n117) );
  DFF_X1 \mem_reg[2][5]  ( .D(n69), .CK(clk), .QN(n116) );
  DFF_X1 \mem_reg[2][4]  ( .D(n70), .CK(clk), .QN(n115) );
  DFF_X1 \mem_reg[2][3]  ( .D(n71), .CK(clk), .QN(n114) );
  DFF_X1 \mem_reg[2][2]  ( .D(n72), .CK(clk), .QN(n113) );
  DFF_X1 \mem_reg[2][1]  ( .D(n73), .CK(clk), .QN(n112) );
  DFF_X1 \mem_reg[2][0]  ( .D(n74), .CK(clk), .QN(n111) );
  DFF_X1 \mem_reg[1][7]  ( .D(n75), .CK(clk), .QN(n110) );
  DFF_X1 \mem_reg[1][6]  ( .D(n76), .CK(clk), .QN(n109) );
  DFF_X1 \mem_reg[1][5]  ( .D(n77), .CK(clk), .QN(n108) );
  DFF_X1 \mem_reg[1][4]  ( .D(n78), .CK(clk), .QN(n107) );
  DFF_X1 \mem_reg[1][3]  ( .D(n79), .CK(clk), .QN(n106) );
  DFF_X1 \mem_reg[1][2]  ( .D(n80), .CK(clk), .QN(n105) );
  DFF_X1 \mem_reg[1][1]  ( .D(n81), .CK(clk), .QN(n104) );
  DFF_X1 \mem_reg[1][0]  ( .D(n82), .CK(clk), .QN(n103) );
  DFF_X1 \mem_reg[0][7]  ( .D(n83), .CK(clk), .QN(n102) );
  DFF_X1 \data_out_reg[7]  ( .D(N10), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n84), .CK(clk), .QN(n101) );
  DFF_X1 \data_out_reg[6]  ( .D(N11), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n85), .CK(clk), .QN(n100) );
  DFF_X1 \data_out_reg[5]  ( .D(N12), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n86), .CK(clk), .QN(n99) );
  DFF_X1 \data_out_reg[4]  ( .D(N13), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n87), .CK(clk), .QN(n98) );
  DFF_X1 \data_out_reg[3]  ( .D(N14), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n88), .CK(clk), .QN(n97) );
  DFF_X1 \data_out_reg[2]  ( .D(N15), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n89), .CK(clk), .QN(n96) );
  DFF_X1 \data_out_reg[1]  ( .D(N16), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n90), .CK(clk), .QN(n95) );
  DFF_X1 \data_out_reg[0]  ( .D(N17), .CK(clk), .Q(data_out[0]) );
  NOR3_X2 U20 ( .A1(n28), .A2(addr[1]), .A3(n37), .ZN(n92) );
  NOR3_X2 U29 ( .A1(n28), .A2(addr[0]), .A3(n38), .ZN(n91) );
  INV_X1 U3 ( .A(n94), .ZN(n25) );
  NOR2_X1 U4 ( .A1(n28), .A2(n93), .ZN(n94) );
  NAND2_X1 U5 ( .A1(n37), .A2(n38), .ZN(n93) );
  INV_X1 U6 ( .A(n92), .ZN(n26) );
  INV_X1 U7 ( .A(n91), .ZN(n27) );
  INV_X1 U8 ( .A(wr_en), .ZN(n28) );
  INV_X1 U9 ( .A(addr[1]), .ZN(n38) );
  INV_X1 U10 ( .A(addr[0]), .ZN(n37) );
  OAI222_X1 U11 ( .A1(n37), .A2(n103), .B1(n93), .B2(n95), .C1(n38), .C2(n111), 
        .ZN(N17) );
  OAI222_X1 U12 ( .A1(n37), .A2(n104), .B1(n93), .B2(n96), .C1(n38), .C2(n112), 
        .ZN(N16) );
  OAI222_X1 U13 ( .A1(n37), .A2(n105), .B1(n93), .B2(n97), .C1(n38), .C2(n113), 
        .ZN(N15) );
  OAI222_X1 U14 ( .A1(n37), .A2(n106), .B1(n93), .B2(n98), .C1(n38), .C2(n114), 
        .ZN(N14) );
  OAI222_X1 U15 ( .A1(n37), .A2(n107), .B1(n93), .B2(n99), .C1(n38), .C2(n115), 
        .ZN(N13) );
  OAI222_X1 U16 ( .A1(n37), .A2(n108), .B1(n93), .B2(n100), .C1(n38), .C2(n116), .ZN(N12) );
  OAI222_X1 U17 ( .A1(n37), .A2(n109), .B1(n93), .B2(n101), .C1(n38), .C2(n117), .ZN(N11) );
  OAI222_X1 U18 ( .A1(n37), .A2(n110), .B1(n93), .B2(n102), .C1(n38), .C2(n118), .ZN(N10) );
  OAI22_X1 U19 ( .A1(n36), .A2(n27), .B1(n91), .B2(n111), .ZN(n74) );
  OAI22_X1 U21 ( .A1(n35), .A2(n27), .B1(n91), .B2(n112), .ZN(n73) );
  OAI22_X1 U22 ( .A1(n34), .A2(n27), .B1(n91), .B2(n113), .ZN(n72) );
  OAI22_X1 U23 ( .A1(n33), .A2(n27), .B1(n91), .B2(n114), .ZN(n71) );
  OAI22_X1 U24 ( .A1(n32), .A2(n27), .B1(n91), .B2(n115), .ZN(n70) );
  OAI22_X1 U25 ( .A1(n31), .A2(n27), .B1(n91), .B2(n116), .ZN(n69) );
  OAI22_X1 U26 ( .A1(n30), .A2(n27), .B1(n91), .B2(n117), .ZN(n68) );
  OAI22_X1 U27 ( .A1(n29), .A2(n27), .B1(n91), .B2(n118), .ZN(n67) );
  OAI22_X1 U28 ( .A1(n36), .A2(n26), .B1(n92), .B2(n103), .ZN(n82) );
  OAI22_X1 U30 ( .A1(n35), .A2(n26), .B1(n92), .B2(n104), .ZN(n81) );
  OAI22_X1 U31 ( .A1(n34), .A2(n26), .B1(n92), .B2(n105), .ZN(n80) );
  OAI22_X1 U32 ( .A1(n33), .A2(n26), .B1(n92), .B2(n106), .ZN(n79) );
  OAI22_X1 U33 ( .A1(n32), .A2(n26), .B1(n92), .B2(n107), .ZN(n78) );
  OAI22_X1 U34 ( .A1(n31), .A2(n26), .B1(n92), .B2(n108), .ZN(n77) );
  OAI22_X1 U35 ( .A1(n30), .A2(n26), .B1(n92), .B2(n109), .ZN(n76) );
  OAI22_X1 U36 ( .A1(n29), .A2(n26), .B1(n92), .B2(n110), .ZN(n75) );
  OAI22_X1 U37 ( .A1(n25), .A2(n36), .B1(n94), .B2(n95), .ZN(n90) );
  OAI22_X1 U38 ( .A1(n25), .A2(n35), .B1(n94), .B2(n96), .ZN(n89) );
  OAI22_X1 U39 ( .A1(n25), .A2(n34), .B1(n94), .B2(n97), .ZN(n88) );
  OAI22_X1 U40 ( .A1(n25), .A2(n33), .B1(n94), .B2(n98), .ZN(n87) );
  OAI22_X1 U41 ( .A1(n25), .A2(n32), .B1(n94), .B2(n99), .ZN(n86) );
  OAI22_X1 U42 ( .A1(n25), .A2(n31), .B1(n94), .B2(n100), .ZN(n85) );
  OAI22_X1 U43 ( .A1(n25), .A2(n30), .B1(n94), .B2(n101), .ZN(n84) );
  OAI22_X1 U44 ( .A1(n25), .A2(n29), .B1(n94), .B2(n102), .ZN(n83) );
  INV_X1 U45 ( .A(data_in[0]), .ZN(n36) );
  INV_X1 U46 ( .A(data_in[1]), .ZN(n35) );
  INV_X1 U47 ( .A(data_in[2]), .ZN(n34) );
  INV_X1 U48 ( .A(data_in[3]), .ZN(n33) );
  INV_X1 U49 ( .A(data_in[4]), .ZN(n32) );
  INV_X1 U50 ( .A(data_in[5]), .ZN(n31) );
  INV_X1 U51 ( .A(data_in[6]), .ZN(n30) );
  INV_X1 U52 ( .A(data_in[7]), .ZN(n29) );
endmodule


module part2_mac_DW_mult_tc_2 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n16, n18, n20,
         n21, n22, n23, n24, n25, n27, n29, n30, n31, n32, n33, n34, n35, n36,
         n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n72, n74, n75, n76, n77, n78, n79, n80, n81, n82, n84,
         n86, n87, n89, n91, n92, n93, n94, n95, n96, n97, n100, n101, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n152, n153, n154, n155, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n238, n239, n240, n241, n246, n247, n248, n249, n251,
         n253, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324;
  assign product[15] = n16;

  FA_X1 U120 ( .A(n163), .B(n110), .CI(n168), .CO(n106), .S(n107) );
  FA_X1 U121 ( .A(n111), .B(n169), .CI(n114), .CO(n108), .S(n109) );
  FA_X1 U123 ( .A(n118), .B(n164), .CI(n115), .CO(n112), .S(n113) );
  FA_X1 U124 ( .A(n170), .B(n120), .CI(n177), .CO(n114), .S(n115) );
  FA_X1 U125 ( .A(n124), .B(n126), .CI(n119), .CO(n116), .S(n117) );
  FA_X1 U126 ( .A(n171), .B(n178), .CI(n121), .CO(n118), .S(n119) );
  FA_X1 U129 ( .A(n186), .B(n172), .CI(n132), .CO(n124), .S(n125) );
  FA_X1 U132 ( .A(n136), .B(n133), .CI(n131), .CO(n128), .S(n129) );
  FA_X1 U133 ( .A(n173), .B(n180), .CI(n187), .CO(n130), .S(n131) );
  HA_X1 U134 ( .A(n158), .B(n166), .CO(n132), .S(n133) );
  FA_X1 U136 ( .A(n181), .B(n167), .CI(n174), .CO(n136), .S(n137) );
  HA_X1 U138 ( .A(n159), .B(n182), .CO(n140), .S(n141) );
  FA_X1 U139 ( .A(n183), .B(n176), .CI(n190), .CO(n142), .S(n143) );
  HA_X1 U140 ( .A(n184), .B(n160), .CO(n144), .S(n145) );
  XNOR2_X1 U260 ( .A(n179), .B(n165), .ZN(n127) );
  OAI22_X1 U261 ( .A1(n261), .A2(n224), .B1(n223), .B2(n249), .ZN(n189) );
  AND2_X1 U262 ( .A1(n322), .A2(n89), .ZN(product[1]) );
  XOR2_X1 U263 ( .A(n175), .B(n189), .Z(n296) );
  XOR2_X1 U264 ( .A(n141), .B(n296), .Z(n139) );
  NAND2_X1 U265 ( .A1(n141), .A2(n175), .ZN(n297) );
  NAND2_X1 U266 ( .A1(n141), .A2(n189), .ZN(n298) );
  NAND2_X1 U267 ( .A1(n175), .A2(n189), .ZN(n299) );
  NAND3_X1 U268 ( .A1(n297), .A2(n298), .A3(n299), .ZN(n138) );
  CLKBUF_X1 U269 ( .A(n255), .Z(n300) );
  BUF_X2 U270 ( .A(a[5]), .Z(n255) );
  XOR2_X1 U271 ( .A(n140), .B(n188), .Z(n301) );
  XOR2_X1 U272 ( .A(n137), .B(n301), .Z(n135) );
  NAND2_X1 U273 ( .A1(n137), .A2(n140), .ZN(n302) );
  NAND2_X1 U274 ( .A1(n137), .A2(n188), .ZN(n303) );
  NAND2_X1 U275 ( .A1(n140), .A2(n188), .ZN(n304) );
  NAND3_X1 U276 ( .A1(n302), .A2(n303), .A3(n304), .ZN(n134) );
  NOR2_X2 U277 ( .A1(n129), .A2(n134), .ZN(n64) );
  INV_X1 U278 ( .A(n251), .ZN(n305) );
  NAND2_X2 U279 ( .A1(n239), .A2(n263), .ZN(n259) );
  BUF_X2 U280 ( .A(n263), .Z(n247) );
  XOR2_X1 U281 ( .A(n130), .B(n127), .Z(n306) );
  XOR2_X1 U282 ( .A(n125), .B(n306), .Z(n123) );
  NAND2_X1 U283 ( .A1(n125), .A2(n130), .ZN(n307) );
  NAND2_X1 U284 ( .A1(n125), .A2(n127), .ZN(n308) );
  NAND2_X1 U285 ( .A1(n130), .A2(n127), .ZN(n309) );
  NAND3_X1 U286 ( .A1(n307), .A2(n308), .A3(n309), .ZN(n122) );
  BUF_X2 U287 ( .A(n262), .Z(n246) );
  CLKBUF_X3 U288 ( .A(a[3]), .Z(n256) );
  OR2_X1 U289 ( .A1(n135), .A2(n138), .ZN(n310) );
  NOR2_X1 U290 ( .A1(n123), .A2(n128), .ZN(n311) );
  NAND2_X1 U291 ( .A1(n240), .A2(n264), .ZN(n312) );
  AOI21_X1 U292 ( .B1(n320), .B2(n75), .A(n72), .ZN(n313) );
  NAND2_X1 U293 ( .A1(n59), .A2(n67), .ZN(n314) );
  INV_X1 U294 ( .A(n60), .ZN(n315) );
  AND2_X2 U295 ( .A1(n314), .A2(n315), .ZN(n58) );
  CLKBUF_X1 U296 ( .A(n258), .Z(n316) );
  OR2_X1 U297 ( .A1(n39), .A2(n30), .ZN(n317) );
  NOR2_X1 U298 ( .A1(n123), .A2(n128), .ZN(n61) );
  OR2_X1 U299 ( .A1(n162), .A2(n104), .ZN(n318) );
  XNOR2_X1 U300 ( .A(n319), .B(n78), .ZN(product[4]) );
  AND2_X1 U301 ( .A1(n100), .A2(n77), .ZN(n319) );
  OR2_X1 U302 ( .A1(n139), .A2(n142), .ZN(n320) );
  OR2_X1 U303 ( .A1(n192), .A2(n185), .ZN(n321) );
  OR2_X1 U304 ( .A1(n193), .A2(n161), .ZN(n322) );
  NAND2_X1 U305 ( .A1(n241), .A2(n265), .ZN(n261) );
  NAND2_X1 U306 ( .A1(n240), .A2(n264), .ZN(n260) );
  INV_X1 U307 ( .A(n146), .ZN(n162) );
  NAND2_X1 U308 ( .A1(n318), .A2(n20), .ZN(n2) );
  INV_X1 U309 ( .A(n20), .ZN(n18) );
  NAND2_X1 U310 ( .A1(n162), .A2(n104), .ZN(n20) );
  NAND2_X1 U311 ( .A1(n91), .A2(n31), .ZN(n3) );
  NAND2_X1 U312 ( .A1(n106), .A2(n105), .ZN(n31) );
  NOR2_X1 U313 ( .A1(n109), .A2(n112), .ZN(n46) );
  NAND2_X1 U314 ( .A1(n93), .A2(n47), .ZN(n5) );
  INV_X1 U315 ( .A(n47), .ZN(n45) );
  NAND2_X1 U316 ( .A1(n109), .A2(n112), .ZN(n47) );
  BUF_X2 U317 ( .A(n265), .Z(n249) );
  INV_X1 U318 ( .A(n30), .ZN(n91) );
  NOR2_X1 U319 ( .A1(n106), .A2(n105), .ZN(n30) );
  INV_X1 U320 ( .A(n29), .ZN(n27) );
  CLKBUF_X1 U321 ( .A(a[7]), .Z(n323) );
  OAI22_X1 U322 ( .A1(n261), .A2(n227), .B1(n226), .B2(n249), .ZN(n192) );
  OAI21_X1 U323 ( .B1(n53), .B2(n57), .A(n54), .ZN(n52) );
  NOR2_X1 U324 ( .A1(n113), .A2(n116), .ZN(n53) );
  OAI22_X1 U325 ( .A1(n261), .A2(n253), .B1(n229), .B2(n249), .ZN(n161) );
  OAI22_X1 U326 ( .A1(n261), .A2(n228), .B1(n227), .B2(n249), .ZN(n193) );
  INV_X1 U327 ( .A(n56), .ZN(n95) );
  OR2_X1 U328 ( .A1(b[0]), .A2(n157), .ZN(n229) );
  OR2_X1 U329 ( .A1(b[0]), .A2(n154), .ZN(n220) );
  NOR2_X1 U330 ( .A1(n56), .A2(n53), .ZN(n51) );
  NAND2_X1 U331 ( .A1(n238), .A2(n262), .ZN(n258) );
  NOR2_X1 U332 ( .A1(n145), .A2(n191), .ZN(n80) );
  OAI21_X1 U333 ( .B1(n317), .B2(n47), .A(n27), .ZN(n25) );
  NAND2_X1 U334 ( .A1(n143), .A2(n144), .ZN(n77) );
  NAND2_X1 U335 ( .A1(n108), .A2(n107), .ZN(n40) );
  NAND2_X1 U336 ( .A1(n97), .A2(n65), .ZN(n9) );
  INV_X1 U337 ( .A(n89), .ZN(n87) );
  CLKBUF_X3 U338 ( .A(a[1]), .Z(n257) );
  XNOR2_X1 U339 ( .A(b[5]), .B(n323), .ZN(n196) );
  XNOR2_X1 U340 ( .A(n323), .B(b[0]), .ZN(n201) );
  XNOR2_X1 U341 ( .A(b[3]), .B(n323), .ZN(n198) );
  INV_X1 U342 ( .A(n86), .ZN(n84) );
  AND2_X1 U343 ( .A1(b[0]), .A2(n153), .ZN(n185) );
  NAND2_X1 U344 ( .A1(n92), .A2(n40), .ZN(n4) );
  OAI21_X1 U345 ( .B1(n47), .B2(n39), .A(n40), .ZN(n36) );
  XNOR2_X1 U346 ( .A(b[7]), .B(n324), .ZN(n194) );
  OR2_X1 U347 ( .A1(b[0]), .A2(n148), .ZN(n202) );
  NAND2_X1 U348 ( .A1(n129), .A2(n134), .ZN(n65) );
  NAND2_X1 U349 ( .A1(n135), .A2(n138), .ZN(n69) );
  NOR2_X1 U350 ( .A1(n135), .A2(n138), .ZN(n68) );
  NOR2_X1 U351 ( .A1(n143), .A2(n144), .ZN(n76) );
  AND2_X1 U352 ( .A1(b[0]), .A2(n147), .ZN(n167) );
  INV_X1 U353 ( .A(n76), .ZN(n100) );
  AOI21_X1 U354 ( .B1(n321), .B2(n87), .A(n84), .ZN(n82) );
  OAI21_X1 U355 ( .B1(n61), .B2(n65), .A(n62), .ZN(n60) );
  INV_X1 U356 ( .A(n74), .ZN(n72) );
  OR2_X1 U357 ( .A1(b[0]), .A2(n251), .ZN(n211) );
  AOI21_X1 U358 ( .B1(n320), .B2(n75), .A(n72), .ZN(n70) );
  NAND2_X1 U359 ( .A1(n123), .A2(n128), .ZN(n62) );
  INV_X1 U360 ( .A(n80), .ZN(n101) );
  OAI21_X1 U361 ( .B1(n76), .B2(n78), .A(n77), .ZN(n75) );
  OAI21_X1 U362 ( .B1(n58), .B2(n22), .A(n23), .ZN(n21) );
  INV_X1 U363 ( .A(n53), .ZN(n94) );
  NAND2_X1 U364 ( .A1(n94), .A2(n54), .ZN(n6) );
  INV_X1 U365 ( .A(n51), .ZN(n49) );
  NAND2_X1 U366 ( .A1(n51), .A2(n93), .ZN(n42) );
  NAND2_X1 U367 ( .A1(n51), .A2(n35), .ZN(n33) );
  NAND2_X1 U368 ( .A1(n51), .A2(n24), .ZN(n22) );
  INV_X1 U369 ( .A(n52), .ZN(n50) );
  AOI21_X1 U370 ( .B1(n52), .B2(n93), .A(n45), .ZN(n43) );
  AOI21_X1 U371 ( .B1(n52), .B2(n35), .A(n36), .ZN(n34) );
  AOI21_X1 U372 ( .B1(n52), .B2(n24), .A(n25), .ZN(n23) );
  NAND2_X1 U373 ( .A1(n113), .A2(n116), .ZN(n54) );
  INV_X1 U374 ( .A(n247), .ZN(n150) );
  OAI22_X1 U375 ( .A1(n259), .A2(n210), .B1(n209), .B2(n247), .ZN(n175) );
  OAI22_X1 U376 ( .A1(n259), .A2(n209), .B1(n208), .B2(n247), .ZN(n174) );
  OAI22_X1 U377 ( .A1(n259), .A2(n208), .B1(n207), .B2(n247), .ZN(n173) );
  OAI22_X1 U378 ( .A1(n259), .A2(n207), .B1(n206), .B2(n247), .ZN(n172) );
  OAI22_X1 U379 ( .A1(n259), .A2(n206), .B1(n205), .B2(n247), .ZN(n171) );
  OAI22_X1 U380 ( .A1(n259), .A2(n205), .B1(n204), .B2(n247), .ZN(n170) );
  OAI22_X1 U381 ( .A1(n259), .A2(n204), .B1(n203), .B2(n247), .ZN(n169) );
  AOI21_X1 U382 ( .B1(n259), .B2(n247), .A(n203), .ZN(n149) );
  OAI22_X1 U383 ( .A1(n259), .A2(n251), .B1(n211), .B2(n247), .ZN(n159) );
  AND2_X1 U384 ( .A1(b[0]), .A2(n150), .ZN(n176) );
  INV_X1 U385 ( .A(n149), .ZN(n168) );
  INV_X1 U386 ( .A(n311), .ZN(n96) );
  NAND2_X1 U387 ( .A1(n95), .A2(n57), .ZN(n7) );
  NOR2_X1 U388 ( .A1(n117), .A2(n122), .ZN(n56) );
  OAI22_X1 U389 ( .A1(n316), .A2(n195), .B1(n246), .B2(n194), .ZN(n104) );
  OAI22_X1 U390 ( .A1(n258), .A2(n197), .B1(n246), .B2(n196), .ZN(n110) );
  INV_X1 U391 ( .A(n246), .ZN(n147) );
  XOR2_X1 U392 ( .A(a[6]), .B(a[7]), .Z(n238) );
  XNOR2_X1 U393 ( .A(a[3]), .B(a[4]), .ZN(n263) );
  OAI22_X1 U394 ( .A1(n261), .A2(n226), .B1(n225), .B2(n249), .ZN(n191) );
  OAI22_X1 U395 ( .A1(n261), .A2(n225), .B1(n224), .B2(n249), .ZN(n190) );
  OAI22_X1 U396 ( .A1(n261), .A2(n223), .B1(n222), .B2(n249), .ZN(n188) );
  OAI22_X1 U397 ( .A1(n261), .A2(n222), .B1(n221), .B2(n249), .ZN(n187) );
  AOI21_X1 U398 ( .B1(n261), .B2(n249), .A(n221), .ZN(n155) );
  NAND2_X1 U399 ( .A1(n193), .A2(n161), .ZN(n89) );
  NAND2_X1 U400 ( .A1(n192), .A2(n185), .ZN(n86) );
  NAND2_X1 U401 ( .A1(n145), .A2(n191), .ZN(n81) );
  INV_X1 U402 ( .A(n155), .ZN(n186) );
  INV_X1 U403 ( .A(n104), .ZN(n105) );
  NAND2_X1 U404 ( .A1(n139), .A2(n142), .ZN(n74) );
  INV_X1 U405 ( .A(n110), .ZN(n111) );
  XOR2_X1 U406 ( .A(a[0]), .B(a[1]), .Z(n241) );
  NAND2_X1 U407 ( .A1(n117), .A2(n122), .ZN(n57) );
  XNOR2_X1 U408 ( .A(b[6]), .B(n324), .ZN(n195) );
  XNOR2_X1 U409 ( .A(b[1]), .B(n323), .ZN(n200) );
  BUF_X2 U410 ( .A(a[7]), .Z(n324) );
  XOR2_X1 U411 ( .A(a[5]), .B(a[4]), .Z(n239) );
  INV_X1 U412 ( .A(n79), .ZN(n78) );
  OAI21_X1 U413 ( .B1(n80), .B2(n82), .A(n81), .ZN(n79) );
  INV_X1 U414 ( .A(n39), .ZN(n92) );
  NOR2_X1 U415 ( .A1(n108), .A2(n107), .ZN(n39) );
  XNOR2_X1 U416 ( .A(b[4]), .B(n324), .ZN(n197) );
  XNOR2_X1 U417 ( .A(b[2]), .B(n324), .ZN(n199) );
  INV_X1 U418 ( .A(n324), .ZN(n148) );
  INV_X1 U419 ( .A(n248), .ZN(n153) );
  OAI22_X1 U420 ( .A1(n260), .A2(n219), .B1(n218), .B2(n248), .ZN(n184) );
  OAI22_X1 U421 ( .A1(n312), .A2(n218), .B1(n217), .B2(n248), .ZN(n183) );
  OAI22_X1 U422 ( .A1(n260), .A2(n217), .B1(n216), .B2(n248), .ZN(n182) );
  OAI22_X1 U423 ( .A1(n260), .A2(n216), .B1(n215), .B2(n248), .ZN(n181) );
  OAI22_X1 U424 ( .A1(n312), .A2(n215), .B1(n214), .B2(n248), .ZN(n180) );
  OAI22_X1 U425 ( .A1(n260), .A2(n214), .B1(n213), .B2(n248), .ZN(n179) );
  OAI22_X1 U426 ( .A1(n312), .A2(n213), .B1(n212), .B2(n248), .ZN(n178) );
  AOI21_X1 U427 ( .B1(n260), .B2(n248), .A(n212), .ZN(n152) );
  OAI22_X1 U428 ( .A1(n312), .A2(n154), .B1(n220), .B2(n248), .ZN(n160) );
  BUF_X2 U429 ( .A(n264), .Z(n248) );
  OR2_X1 U430 ( .A1(n179), .A2(n165), .ZN(n126) );
  INV_X1 U431 ( .A(n152), .ZN(n177) );
  OAI21_X1 U432 ( .B1(n40), .B2(n30), .A(n31), .ZN(n29) );
  INV_X1 U433 ( .A(n64), .ZN(n97) );
  NOR2_X1 U434 ( .A1(n311), .A2(n64), .ZN(n59) );
  XNOR2_X1 U435 ( .A(a[1]), .B(a[2]), .ZN(n264) );
  XOR2_X1 U436 ( .A(a[3]), .B(a[2]), .Z(n240) );
  INV_X1 U437 ( .A(n46), .ZN(n93) );
  NOR2_X1 U438 ( .A1(n46), .A2(n39), .ZN(n35) );
  NOR2_X1 U439 ( .A1(n46), .A2(n317), .ZN(n24) );
  AOI21_X1 U440 ( .B1(n316), .B2(n246), .A(n194), .ZN(n146) );
  OAI22_X1 U441 ( .A1(n316), .A2(n198), .B1(n246), .B2(n197), .ZN(n164) );
  OAI22_X1 U442 ( .A1(n316), .A2(n196), .B1(n246), .B2(n195), .ZN(n163) );
  OAI22_X1 U443 ( .A1(n258), .A2(n200), .B1(n246), .B2(n199), .ZN(n165) );
  OAI22_X1 U444 ( .A1(n258), .A2(n201), .B1(n246), .B2(n200), .ZN(n166) );
  OAI21_X1 U445 ( .B1(n68), .B2(n70), .A(n69), .ZN(n67) );
  XNOR2_X1 U446 ( .A(n305), .B(b[0]), .ZN(n210) );
  XNOR2_X1 U447 ( .A(n305), .B(b[7]), .ZN(n203) );
  XNOR2_X1 U448 ( .A(n300), .B(b[6]), .ZN(n204) );
  INV_X1 U449 ( .A(n255), .ZN(n251) );
  XNOR2_X1 U450 ( .A(n300), .B(b[5]), .ZN(n205) );
  XNOR2_X1 U451 ( .A(n300), .B(b[4]), .ZN(n206) );
  XNOR2_X1 U452 ( .A(n255), .B(b[1]), .ZN(n209) );
  XNOR2_X1 U453 ( .A(n255), .B(b[3]), .ZN(n207) );
  XNOR2_X1 U454 ( .A(n255), .B(b[2]), .ZN(n208) );
  OAI22_X1 U455 ( .A1(n258), .A2(n148), .B1(n202), .B2(n246), .ZN(n158) );
  XNOR2_X1 U456 ( .A(n256), .B(b[6]), .ZN(n213) );
  XNOR2_X1 U457 ( .A(n256), .B(b[2]), .ZN(n217) );
  XNOR2_X1 U458 ( .A(n256), .B(b[3]), .ZN(n216) );
  XNOR2_X1 U459 ( .A(n256), .B(b[7]), .ZN(n212) );
  XNOR2_X1 U460 ( .A(n256), .B(b[0]), .ZN(n219) );
  XNOR2_X1 U461 ( .A(n256), .B(b[5]), .ZN(n214) );
  XNOR2_X1 U462 ( .A(n256), .B(b[4]), .ZN(n215) );
  XNOR2_X1 U463 ( .A(n256), .B(b[1]), .ZN(n218) );
  INV_X1 U464 ( .A(a[3]), .ZN(n154) );
  XNOR2_X1 U465 ( .A(n257), .B(b[5]), .ZN(n223) );
  XNOR2_X1 U466 ( .A(n257), .B(b[3]), .ZN(n225) );
  XNOR2_X1 U467 ( .A(n257), .B(b[4]), .ZN(n224) );
  INV_X1 U468 ( .A(n257), .ZN(n253) );
  XNOR2_X1 U469 ( .A(n257), .B(b[6]), .ZN(n222) );
  XNOR2_X1 U470 ( .A(n257), .B(b[7]), .ZN(n221) );
  XNOR2_X1 U471 ( .A(n257), .B(b[0]), .ZN(n228) );
  XNOR2_X1 U472 ( .A(n257), .B(b[2]), .ZN(n226) );
  XNOR2_X1 U473 ( .A(n257), .B(b[1]), .ZN(n227) );
  INV_X1 U474 ( .A(n257), .ZN(n157) );
  INV_X1 U475 ( .A(n120), .ZN(n121) );
  OAI22_X1 U476 ( .A1(n258), .A2(n199), .B1(n246), .B2(n198), .ZN(n120) );
  INV_X1 U477 ( .A(a[0]), .ZN(n265) );
  XNOR2_X1 U478 ( .A(a[5]), .B(a[6]), .ZN(n262) );
  AND2_X1 U479 ( .A1(b[0]), .A2(a[0]), .ZN(product[0]) );
  XNOR2_X1 U480 ( .A(n14), .B(n87), .ZN(product[2]) );
  NAND2_X1 U481 ( .A1(n321), .A2(n86), .ZN(n14) );
  NAND2_X1 U482 ( .A1(n310), .A2(n69), .ZN(n10) );
  XOR2_X1 U483 ( .A(n10), .B(n313), .Z(product[6]) );
  XOR2_X1 U484 ( .A(n13), .B(n82), .Z(product[3]) );
  NAND2_X1 U485 ( .A1(n101), .A2(n81), .ZN(n13) );
  XNOR2_X1 U486 ( .A(n11), .B(n75), .ZN(product[5]) );
  NAND2_X1 U487 ( .A1(n320), .A2(n74), .ZN(n11) );
  NAND2_X1 U488 ( .A1(n96), .A2(n62), .ZN(n8) );
  AOI21_X1 U489 ( .B1(n21), .B2(n318), .A(n18), .ZN(n16) );
  XNOR2_X1 U490 ( .A(n63), .B(n8), .ZN(product[8]) );
  OAI21_X1 U491 ( .B1(n66), .B2(n64), .A(n65), .ZN(n63) );
  XOR2_X1 U492 ( .A(n66), .B(n9), .Z(product[7]) );
  INV_X1 U493 ( .A(n67), .ZN(n66) );
  XOR2_X1 U494 ( .A(n58), .B(n7), .Z(product[9]) );
  XNOR2_X1 U495 ( .A(n41), .B(n4), .ZN(product[12]) );
  OAI21_X1 U496 ( .B1(n58), .B2(n42), .A(n43), .ZN(n41) );
  XNOR2_X1 U497 ( .A(n32), .B(n3), .ZN(product[13]) );
  OAI21_X1 U498 ( .B1(n58), .B2(n33), .A(n34), .ZN(n32) );
  XNOR2_X1 U499 ( .A(n21), .B(n2), .ZN(product[14]) );
  XNOR2_X1 U500 ( .A(n55), .B(n6), .ZN(product[10]) );
  OAI21_X1 U501 ( .B1(n58), .B2(n56), .A(n57), .ZN(n55) );
  XNOR2_X1 U502 ( .A(n48), .B(n5), .ZN(product[11]) );
  OAI21_X1 U503 ( .B1(n58), .B2(n49), .A(n50), .ZN(n48) );
endmodule


module part2_mac_DW01_add_2 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n19, n20, n21, n22, n24, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n46, n47, n48, n50,
         n52, n53, n54, n55, n56, n58, n60, n61, n62, n63, n64, n66, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n78, n80, n81, n83, n86, n87, n88,
         n89, n90, n94, n96, n97, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n170, n171;

  NOR2_X2 U119 ( .A1(B[9]), .A2(A[9]), .ZN(n46) );
  OR2_X1 U120 ( .A1(B[7]), .A2(A[7]), .ZN(n154) );
  OAI21_X1 U121 ( .B1(n48), .B2(n46), .A(n47), .ZN(n155) );
  CLKBUF_X1 U122 ( .A(n61), .Z(n156) );
  AOI21_X1 U123 ( .B1(n53), .B2(n165), .A(n50), .ZN(n157) );
  AOI21_X1 U124 ( .B1(n53), .B2(n165), .A(n50), .ZN(n48) );
  NOR2_X1 U125 ( .A1(B[11]), .A2(A[11]), .ZN(n158) );
  CLKBUF_X1 U126 ( .A(n53), .Z(n159) );
  OAI21_X1 U127 ( .B1(n48), .B2(n46), .A(n47), .ZN(n160) );
  OAI21_X1 U128 ( .B1(n157), .B2(n46), .A(n47), .ZN(n161) );
  AOI21_X1 U129 ( .B1(n166), .B2(n156), .A(n58), .ZN(n162) );
  AOI21_X1 U130 ( .B1(n155), .B2(n37), .A(n38), .ZN(n163) );
  OR2_X1 U131 ( .A1(B[14]), .A2(A[14]), .ZN(n164) );
  OR2_X1 U132 ( .A1(B[8]), .A2(A[8]), .ZN(n165) );
  OR2_X1 U133 ( .A1(B[6]), .A2(A[6]), .ZN(n166) );
  OR2_X1 U134 ( .A1(B[4]), .A2(A[4]), .ZN(n167) );
  OR2_X1 U135 ( .A1(B[1]), .A2(A[1]), .ZN(n168) );
  AND2_X1 U136 ( .A1(n171), .A2(n83), .ZN(SUM[0]) );
  OR2_X1 U137 ( .A1(B[15]), .A2(A[15]), .ZN(n170) );
  OR2_X1 U138 ( .A1(B[0]), .A2(A[0]), .ZN(n171) );
  INV_X1 U139 ( .A(n83), .ZN(n81) );
  NAND2_X1 U140 ( .A1(B[0]), .A2(A[0]), .ZN(n83) );
  NOR2_X1 U141 ( .A1(B[11]), .A2(A[11]), .ZN(n39) );
  NAND2_X1 U142 ( .A1(B[15]), .A2(A[15]), .ZN(n19) );
  NAND2_X1 U143 ( .A1(n170), .A2(n19), .ZN(n2) );
  NAND2_X1 U144 ( .A1(B[2]), .A2(A[2]), .ZN(n75) );
  NAND2_X1 U145 ( .A1(n164), .A2(n26), .ZN(n3) );
  NAND2_X1 U146 ( .A1(n86), .A2(n33), .ZN(n4) );
  NAND2_X1 U147 ( .A1(B[13]), .A2(A[13]), .ZN(n33) );
  NAND2_X1 U148 ( .A1(B[9]), .A2(A[9]), .ZN(n47) );
  NAND2_X1 U149 ( .A1(B[14]), .A2(A[14]), .ZN(n26) );
  NAND2_X1 U150 ( .A1(n87), .A2(n36), .ZN(n5) );
  NAND2_X1 U151 ( .A1(B[12]), .A2(A[12]), .ZN(n36) );
  NOR2_X1 U152 ( .A1(A[10]), .A2(B[10]), .ZN(n42) );
  INV_X1 U153 ( .A(n74), .ZN(n97) );
  NOR2_X1 U154 ( .A1(B[2]), .A2(A[2]), .ZN(n74) );
  NAND2_X1 U155 ( .A1(B[3]), .A2(A[3]), .ZN(n71) );
  INV_X1 U156 ( .A(n30), .ZN(n28) );
  NOR2_X1 U157 ( .A1(n35), .A2(n32), .ZN(n30) );
  NAND2_X1 U158 ( .A1(n88), .A2(n40), .ZN(n6) );
  NOR2_X1 U159 ( .A1(B[13]), .A2(A[13]), .ZN(n32) );
  NAND2_X1 U160 ( .A1(B[5]), .A2(A[5]), .ZN(n63) );
  NAND2_X1 U161 ( .A1(n89), .A2(n43), .ZN(n7) );
  INV_X1 U162 ( .A(n26), .ZN(n24) );
  NAND2_X1 U163 ( .A1(B[7]), .A2(A[7]), .ZN(n55) );
  NAND2_X1 U164 ( .A1(n30), .A2(n164), .ZN(n21) );
  NAND2_X1 U165 ( .A1(B[11]), .A2(A[11]), .ZN(n40) );
  NAND2_X1 U166 ( .A1(B[10]), .A2(A[10]), .ZN(n43) );
  INV_X1 U167 ( .A(n80), .ZN(n78) );
  NAND2_X1 U168 ( .A1(B[1]), .A2(A[1]), .ZN(n80) );
  INV_X1 U169 ( .A(n31), .ZN(n29) );
  AOI21_X1 U170 ( .B1(n31), .B2(n164), .A(n24), .ZN(n22) );
  OAI21_X1 U171 ( .B1(n32), .B2(n36), .A(n33), .ZN(n31) );
  INV_X1 U172 ( .A(n70), .ZN(n96) );
  NOR2_X1 U173 ( .A1(B[3]), .A2(A[3]), .ZN(n70) );
  INV_X1 U174 ( .A(n62), .ZN(n94) );
  NOR2_X1 U175 ( .A1(B[5]), .A2(A[5]), .ZN(n62) );
  INV_X1 U176 ( .A(n73), .ZN(n72) );
  NOR2_X1 U177 ( .A1(B[7]), .A2(A[7]), .ZN(n54) );
  AOI21_X1 U178 ( .B1(n168), .B2(n81), .A(n78), .ZN(n76) );
  INV_X1 U179 ( .A(n52), .ZN(n50) );
  NAND2_X1 U180 ( .A1(B[8]), .A2(A[8]), .ZN(n52) );
  INV_X1 U181 ( .A(n60), .ZN(n58) );
  NAND2_X1 U182 ( .A1(B[6]), .A2(A[6]), .ZN(n60) );
  INV_X1 U183 ( .A(n68), .ZN(n66) );
  NAND2_X1 U184 ( .A1(B[4]), .A2(A[4]), .ZN(n68) );
  INV_X1 U185 ( .A(n46), .ZN(n90) );
  AOI21_X1 U186 ( .B1(n69), .B2(n167), .A(n66), .ZN(n64) );
  AOI21_X1 U187 ( .B1(n37), .B2(n160), .A(n38), .ZN(n1) );
  AOI21_X1 U188 ( .B1(n166), .B2(n61), .A(n58), .ZN(n56) );
  OAI21_X1 U189 ( .B1(n62), .B2(n64), .A(n63), .ZN(n61) );
  INV_X1 U190 ( .A(n158), .ZN(n88) );
  OAI21_X1 U191 ( .B1(n39), .B2(n43), .A(n40), .ZN(n38) );
  NOR2_X1 U192 ( .A1(n42), .A2(n158), .ZN(n37) );
  INV_X1 U193 ( .A(n32), .ZN(n86) );
  INV_X1 U194 ( .A(n42), .ZN(n89) );
  INV_X1 U195 ( .A(n35), .ZN(n87) );
  NOR2_X1 U196 ( .A1(B[12]), .A2(A[12]), .ZN(n35) );
  OAI21_X1 U197 ( .B1(n70), .B2(n72), .A(n71), .ZN(n69) );
  OAI21_X1 U198 ( .B1(n74), .B2(n76), .A(n75), .ZN(n73) );
  XNOR2_X1 U199 ( .A(n16), .B(n81), .ZN(SUM[1]) );
  NAND2_X1 U200 ( .A1(n168), .A2(n80), .ZN(n16) );
  XOR2_X1 U201 ( .A(n15), .B(n76), .Z(SUM[2]) );
  NAND2_X1 U202 ( .A1(n97), .A2(n75), .ZN(n15) );
  XOR2_X1 U203 ( .A(n14), .B(n72), .Z(SUM[3]) );
  NAND2_X1 U204 ( .A1(n96), .A2(n71), .ZN(n14) );
  XNOR2_X1 U205 ( .A(n13), .B(n69), .ZN(SUM[4]) );
  NAND2_X1 U206 ( .A1(n167), .A2(n68), .ZN(n13) );
  XOR2_X1 U207 ( .A(n12), .B(n64), .Z(SUM[5]) );
  NAND2_X1 U208 ( .A1(n94), .A2(n63), .ZN(n12) );
  XNOR2_X1 U209 ( .A(n11), .B(n156), .ZN(SUM[6]) );
  NAND2_X1 U210 ( .A1(n166), .A2(n60), .ZN(n11) );
  OAI21_X1 U211 ( .B1(n56), .B2(n54), .A(n55), .ZN(n53) );
  XNOR2_X1 U212 ( .A(n9), .B(n159), .ZN(SUM[8]) );
  NAND2_X1 U213 ( .A1(n165), .A2(n52), .ZN(n9) );
  XOR2_X1 U214 ( .A(n10), .B(n162), .Z(SUM[7]) );
  NAND2_X1 U215 ( .A1(n154), .A2(n55), .ZN(n10) );
  NAND2_X1 U216 ( .A1(n90), .A2(n47), .ZN(n8) );
  XOR2_X1 U217 ( .A(n8), .B(n157), .Z(SUM[9]) );
  XOR2_X1 U218 ( .A(n44), .B(n7), .Z(SUM[10]) );
  INV_X1 U219 ( .A(n161), .ZN(n44) );
  XOR2_X1 U220 ( .A(n163), .B(n5), .Z(SUM[12]) );
  XNOR2_X1 U221 ( .A(n41), .B(n6), .ZN(SUM[11]) );
  OAI21_X1 U222 ( .B1(n44), .B2(n42), .A(n43), .ZN(n41) );
  XNOR2_X1 U223 ( .A(n20), .B(n2), .ZN(SUM[15]) );
  OAI21_X1 U224 ( .B1(n1), .B2(n21), .A(n22), .ZN(n20) );
  XNOR2_X1 U225 ( .A(n27), .B(n3), .ZN(SUM[14]) );
  OAI21_X1 U226 ( .B1(n163), .B2(n28), .A(n29), .ZN(n27) );
  XNOR2_X1 U227 ( .A(n34), .B(n4), .ZN(SUM[13]) );
  OAI21_X1 U228 ( .B1(n1), .B2(n35), .A(n36), .ZN(n34) );
endmodule


module part2_mac ( clk, reset, a, b, valid_in, f, valid_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] f;
  input clk, reset, valid_in;
  output valid_out;
  wire   en_f, N53, N54, n34, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43,
         N42, N41, N40, N39, N38, N37, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77;
  wire   [7:0] ffAOut;
  wire   [7:0] ffBOut;
  wire   [15:0] adderOut;

  DFF_X1 \ffAOut_reg[7]  ( .D(n62), .CK(clk), .Q(ffAOut[7]) );
  DFF_X1 \ffAOut_reg[6]  ( .D(n63), .CK(clk), .Q(ffAOut[6]) );
  DFF_X1 \ffAOut_reg[5]  ( .D(n64), .CK(clk), .Q(ffAOut[5]) );
  DFF_X1 \ffAOut_reg[4]  ( .D(n65), .CK(clk), .Q(ffAOut[4]) );
  DFF_X1 \ffAOut_reg[3]  ( .D(n66), .CK(clk), .Q(ffAOut[3]), .QN(n1) );
  DFF_X1 \ffAOut_reg[2]  ( .D(n67), .CK(clk), .Q(ffAOut[2]) );
  DFF_X1 \ffAOut_reg[1]  ( .D(n68), .CK(clk), .Q(ffAOut[1]), .QN(n5) );
  DFF_X1 \ffAOut_reg[0]  ( .D(n69), .CK(clk), .Q(ffAOut[0]) );
  DFF_X1 \ffBOut_reg[7]  ( .D(n70), .CK(clk), .Q(ffBOut[7]) );
  DFF_X1 \ffBOut_reg[6]  ( .D(n71), .CK(clk), .Q(ffBOut[6]) );
  DFF_X1 \ffBOut_reg[5]  ( .D(n72), .CK(clk), .Q(ffBOut[5]) );
  DFF_X1 \ffBOut_reg[4]  ( .D(n73), .CK(clk), .Q(ffBOut[4]) );
  DFF_X1 \ffBOut_reg[3]  ( .D(n74), .CK(clk), .Q(ffBOut[3]) );
  DFF_X1 \ffBOut_reg[2]  ( .D(n75), .CK(clk), .Q(ffBOut[2]) );
  DFF_X1 \ffBOut_reg[1]  ( .D(n76), .CK(clk), .Q(ffBOut[1]) );
  DFF_X1 \ffBOut_reg[0]  ( .D(n77), .CK(clk), .Q(ffBOut[0]) );
  DFF_X1 en_f_reg ( .D(N53), .CK(clk), .Q(en_f), .QN(n34) );
  DFF_X1 valid_out_reg ( .D(N54), .CK(clk), .Q(valid_out) );
  DFF_X1 \f_reg[15]  ( .D(n46), .CK(clk), .Q(f[15]) );
  DFF_X1 \f_reg[14]  ( .D(n47), .CK(clk), .Q(f[14]) );
  DFF_X1 \f_reg[13]  ( .D(n48), .CK(clk), .Q(f[13]) );
  DFF_X1 \f_reg[12]  ( .D(n49), .CK(clk), .Q(f[12]) );
  DFF_X1 \f_reg[11]  ( .D(n50), .CK(clk), .Q(f[11]) );
  DFF_X1 \f_reg[10]  ( .D(n51), .CK(clk), .Q(f[10]) );
  DFF_X1 \f_reg[9]  ( .D(n52), .CK(clk), .Q(f[9]) );
  DFF_X1 \f_reg[8]  ( .D(n53), .CK(clk), .Q(f[8]) );
  DFF_X1 \f_reg[7]  ( .D(n54), .CK(clk), .Q(f[7]) );
  DFF_X1 \f_reg[6]  ( .D(n55), .CK(clk), .Q(f[6]) );
  DFF_X1 \f_reg[5]  ( .D(n56), .CK(clk), .Q(f[5]) );
  DFF_X1 \f_reg[4]  ( .D(n57), .CK(clk), .Q(f[4]) );
  DFF_X1 \f_reg[3]  ( .D(n58), .CK(clk), .Q(f[3]) );
  DFF_X1 \f_reg[2]  ( .D(n59), .CK(clk), .Q(f[2]) );
  DFF_X1 \f_reg[1]  ( .D(n60), .CK(clk), .Q(f[1]) );
  DFF_X1 \f_reg[0]  ( .D(n61), .CK(clk), .Q(f[0]) );
  part2_mac_DW_mult_tc_2 mult_35 ( .a(ffAOut), .b(ffBOut), .product({N52, N51, 
        N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37})
         );
  part2_mac_DW01_add_2 add_35 ( .A(f), .B({N52, N51, N50, N49, N48, N47, N46, 
        N45, N44, N43, N42, N41, N40, N39, N38, N37}), .CI(1'b0), .SUM(
        adderOut) );
  INV_X1 U3 ( .A(n1), .ZN(n2) );
  INV_X1 U4 ( .A(n7), .ZN(n44) );
  INV_X1 U5 ( .A(n25), .ZN(n42) );
  AND2_X1 U6 ( .A1(n7), .A2(n24), .ZN(n3) );
  AND2_X1 U7 ( .A1(n25), .A2(n24), .ZN(n4) );
  NOR2_X1 U8 ( .A1(reset), .A2(n34), .ZN(N54) );
  NOR2_X1 U9 ( .A1(reset), .A2(n23), .ZN(N53) );
  INV_X1 U10 ( .A(n5), .ZN(n6) );
  OR2_X1 U11 ( .A1(en_f), .A2(reset), .ZN(n7) );
  INV_X1 U12 ( .A(reset), .ZN(n24) );
  AOI22_X1 U13 ( .A1(f[15]), .A2(n44), .B1(adderOut[15]), .B2(n3), .ZN(n8) );
  INV_X1 U14 ( .A(n8), .ZN(n46) );
  AOI22_X1 U15 ( .A1(f[14]), .A2(n44), .B1(adderOut[14]), .B2(n3), .ZN(n9) );
  INV_X1 U16 ( .A(n9), .ZN(n47) );
  AOI22_X1 U17 ( .A1(f[13]), .A2(n44), .B1(adderOut[13]), .B2(n3), .ZN(n10) );
  INV_X1 U18 ( .A(n10), .ZN(n48) );
  AOI22_X1 U19 ( .A1(f[12]), .A2(n44), .B1(adderOut[12]), .B2(n3), .ZN(n11) );
  INV_X1 U20 ( .A(n11), .ZN(n49) );
  AOI22_X1 U21 ( .A1(f[11]), .A2(n44), .B1(adderOut[11]), .B2(n3), .ZN(n12) );
  INV_X1 U22 ( .A(n12), .ZN(n50) );
  AOI22_X1 U23 ( .A1(f[10]), .A2(n44), .B1(adderOut[10]), .B2(n3), .ZN(n13) );
  INV_X1 U24 ( .A(n13), .ZN(n51) );
  AOI22_X1 U25 ( .A1(f[9]), .A2(n44), .B1(adderOut[9]), .B2(n3), .ZN(n14) );
  INV_X1 U26 ( .A(n14), .ZN(n52) );
  AOI22_X1 U27 ( .A1(f[8]), .A2(n44), .B1(adderOut[8]), .B2(n3), .ZN(n15) );
  INV_X1 U28 ( .A(n15), .ZN(n53) );
  AOI22_X1 U29 ( .A1(f[7]), .A2(n44), .B1(adderOut[7]), .B2(n3), .ZN(n16) );
  INV_X1 U30 ( .A(n16), .ZN(n54) );
  AOI22_X1 U31 ( .A1(f[6]), .A2(n44), .B1(adderOut[6]), .B2(n3), .ZN(n17) );
  INV_X1 U32 ( .A(n17), .ZN(n55) );
  AOI22_X1 U33 ( .A1(f[5]), .A2(n44), .B1(adderOut[5]), .B2(n3), .ZN(n18) );
  INV_X1 U34 ( .A(n18), .ZN(n56) );
  AOI22_X1 U35 ( .A1(f[4]), .A2(n44), .B1(adderOut[4]), .B2(n3), .ZN(n19) );
  INV_X1 U36 ( .A(n19), .ZN(n57) );
  AOI22_X1 U37 ( .A1(f[3]), .A2(n44), .B1(adderOut[3]), .B2(n3), .ZN(n20) );
  INV_X1 U38 ( .A(n20), .ZN(n58) );
  AOI22_X1 U39 ( .A1(f[2]), .A2(n44), .B1(adderOut[2]), .B2(n3), .ZN(n21) );
  INV_X1 U40 ( .A(n21), .ZN(n59) );
  AOI22_X1 U41 ( .A1(f[1]), .A2(n44), .B1(adderOut[1]), .B2(n3), .ZN(n22) );
  INV_X1 U42 ( .A(n22), .ZN(n60) );
  INV_X1 U43 ( .A(valid_in), .ZN(n23) );
  NAND2_X1 U44 ( .A1(n24), .A2(n23), .ZN(n25) );
  AOI22_X1 U45 ( .A1(ffAOut[7]), .A2(n42), .B1(a[7]), .B2(n4), .ZN(n26) );
  INV_X1 U46 ( .A(n26), .ZN(n62) );
  AOI22_X1 U47 ( .A1(ffAOut[6]), .A2(n42), .B1(a[6]), .B2(n4), .ZN(n27) );
  INV_X1 U48 ( .A(n27), .ZN(n63) );
  AOI22_X1 U49 ( .A1(ffAOut[5]), .A2(n42), .B1(a[5]), .B2(n4), .ZN(n28) );
  INV_X1 U50 ( .A(n28), .ZN(n64) );
  AOI22_X1 U51 ( .A1(ffAOut[4]), .A2(n42), .B1(a[4]), .B2(n4), .ZN(n29) );
  INV_X1 U52 ( .A(n29), .ZN(n65) );
  AOI22_X1 U53 ( .A1(n2), .A2(n42), .B1(a[3]), .B2(n4), .ZN(n30) );
  INV_X1 U54 ( .A(n30), .ZN(n66) );
  AOI22_X1 U55 ( .A1(ffAOut[2]), .A2(n42), .B1(a[2]), .B2(n4), .ZN(n31) );
  INV_X1 U56 ( .A(n31), .ZN(n67) );
  AOI22_X1 U57 ( .A1(n6), .A2(n42), .B1(a[1]), .B2(n4), .ZN(n32) );
  INV_X1 U58 ( .A(n32), .ZN(n68) );
  AOI22_X1 U59 ( .A1(ffAOut[0]), .A2(n42), .B1(a[0]), .B2(n4), .ZN(n33) );
  INV_X1 U60 ( .A(n33), .ZN(n69) );
  AOI22_X1 U61 ( .A1(ffBOut[7]), .A2(n42), .B1(b[7]), .B2(n4), .ZN(n35) );
  INV_X1 U62 ( .A(n35), .ZN(n70) );
  AOI22_X1 U63 ( .A1(ffBOut[6]), .A2(n42), .B1(b[6]), .B2(n4), .ZN(n36) );
  INV_X1 U64 ( .A(n36), .ZN(n71) );
  AOI22_X1 U65 ( .A1(ffBOut[5]), .A2(n42), .B1(b[5]), .B2(n4), .ZN(n37) );
  INV_X1 U66 ( .A(n37), .ZN(n72) );
  AOI22_X1 U67 ( .A1(ffBOut[4]), .A2(n42), .B1(b[4]), .B2(n4), .ZN(n38) );
  INV_X1 U68 ( .A(n38), .ZN(n73) );
  AOI22_X1 U69 ( .A1(ffBOut[3]), .A2(n42), .B1(b[3]), .B2(n4), .ZN(n39) );
  INV_X1 U70 ( .A(n39), .ZN(n74) );
  AOI22_X1 U71 ( .A1(ffBOut[2]), .A2(n42), .B1(b[2]), .B2(n4), .ZN(n40) );
  INV_X1 U72 ( .A(n40), .ZN(n75) );
  AOI22_X1 U73 ( .A1(ffBOut[1]), .A2(n42), .B1(b[1]), .B2(n4), .ZN(n41) );
  INV_X1 U74 ( .A(n41), .ZN(n76) );
  AOI22_X1 U75 ( .A1(ffBOut[0]), .A2(n42), .B1(b[0]), .B2(n4), .ZN(n43) );
  INV_X1 U76 ( .A(n43), .ZN(n77) );
  AOI22_X1 U77 ( .A1(f[0]), .A2(n44), .B1(adderOut[0]), .B2(n3), .ZN(n45) );
  INV_X1 U78 ( .A(n45), .ZN(n61) );
endmodule


module mvm3_part2_DW01_add_1 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16, n17,
         n18, n19, n20, n22, n24, n25, n26, n27, n28, n30, n32, n33, n34, n35,
         n36, n38, n40, n41, n42, n43, n44, n46, n48, n49, n50, n51, n53, n55,
         n56, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n75, n76, n78, n80, n82, n86, n87, n88, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n160, n161, n162, n163, n164, n165, n166, n167, n168;

  FA_X1 U3 ( .A(A[14]), .B(B[14]), .CI(n17), .CO(n16), .S(SUM[14]) );
  OR2_X1 U108 ( .A1(A[0]), .A2(B[0]), .ZN(n144) );
  CLKBUF_X1 U109 ( .A(n69), .Z(n145) );
  AND2_X1 U110 ( .A1(A[4]), .A2(B[4]), .ZN(n165) );
  CLKBUF_X1 U111 ( .A(n66), .Z(n146) );
  CLKBUF_X1 U112 ( .A(n64), .Z(n147) );
  INV_X1 U113 ( .A(n70), .ZN(n148) );
  CLKBUF_X1 U114 ( .A(n25), .Z(n149) );
  AOI21_X1 U115 ( .B1(n63), .B2(n148), .A(n147), .ZN(n150) );
  OAI21_X1 U116 ( .B1(n168), .B2(n34), .A(n35), .ZN(n151) );
  CLKBUF_X1 U117 ( .A(n20), .Z(n152) );
  OAI21_X1 U118 ( .B1(n150), .B2(n50), .A(n51), .ZN(n153) );
  AOI21_X1 U119 ( .B1(n49), .B2(n157), .A(n46), .ZN(n154) );
  AOI21_X1 U120 ( .B1(n33), .B2(n162), .A(n30), .ZN(n155) );
  XNOR2_X1 U121 ( .A(B[15]), .B(A[15]), .ZN(n156) );
  OR2_X1 U122 ( .A1(A[6]), .A2(B[6]), .ZN(n157) );
  OR2_X1 U123 ( .A1(A[5]), .A2(B[5]), .ZN(n161) );
  OR2_X1 U124 ( .A1(A[4]), .A2(B[4]), .ZN(n160) );
  NOR2_X1 U125 ( .A1(A[3]), .A2(B[3]), .ZN(n158) );
  INV_X1 U126 ( .A(n71), .ZN(n70) );
  INV_X1 U127 ( .A(n24), .ZN(n22) );
  INV_X1 U128 ( .A(n32), .ZN(n30) );
  INV_X1 U129 ( .A(n48), .ZN(n46) );
  NAND2_X1 U130 ( .A1(n160), .A2(n161), .ZN(n50) );
  INV_X1 U131 ( .A(n55), .ZN(n53) );
  NAND2_X1 U132 ( .A1(n80), .A2(n35), .ZN(n6) );
  NAND2_X1 U133 ( .A1(n157), .A2(n48), .ZN(n9) );
  NAND2_X1 U134 ( .A1(n78), .A2(n27), .ZN(n4) );
  INV_X1 U135 ( .A(n26), .ZN(n78) );
  NAND2_X1 U136 ( .A1(n76), .A2(n19), .ZN(n2) );
  INV_X1 U137 ( .A(n18), .ZN(n76) );
  NAND2_X1 U138 ( .A1(n82), .A2(n43), .ZN(n8) );
  INV_X1 U139 ( .A(n42), .ZN(n82) );
  NAND2_X1 U140 ( .A1(n164), .A2(n24), .ZN(n3) );
  NAND2_X1 U141 ( .A1(n162), .A2(n32), .ZN(n5) );
  NAND2_X1 U142 ( .A1(n163), .A2(n40), .ZN(n7) );
  XOR2_X1 U143 ( .A(n56), .B(n10), .Z(SUM[5]) );
  NAND2_X1 U144 ( .A1(n161), .A2(n55), .ZN(n10) );
  AOI21_X1 U145 ( .B1(n61), .B2(n160), .A(n165), .ZN(n56) );
  XOR2_X1 U146 ( .A(n70), .B(n13), .Z(SUM[2]) );
  INV_X1 U147 ( .A(n68), .ZN(n87) );
  XNOR2_X1 U148 ( .A(n61), .B(n11), .ZN(SUM[4]) );
  NAND2_X1 U149 ( .A1(n160), .A2(n60), .ZN(n11) );
  INV_X1 U150 ( .A(n165), .ZN(n60) );
  XNOR2_X1 U151 ( .A(n67), .B(n12), .ZN(SUM[3]) );
  NAND2_X1 U152 ( .A1(n86), .A2(n146), .ZN(n12) );
  INV_X1 U153 ( .A(n34), .ZN(n80) );
  INV_X1 U154 ( .A(n40), .ZN(n38) );
  NAND2_X1 U155 ( .A1(n88), .A2(n73), .ZN(n14) );
  INV_X1 U156 ( .A(n72), .ZN(n88) );
  AND2_X1 U157 ( .A1(n144), .A2(n166), .ZN(SUM[0]) );
  NOR2_X1 U158 ( .A1(A[2]), .A2(B[2]), .ZN(n68) );
  NAND2_X1 U159 ( .A1(A[12]), .A2(B[12]), .ZN(n24) );
  NAND2_X1 U160 ( .A1(A[10]), .A2(B[10]), .ZN(n32) );
  NAND2_X1 U161 ( .A1(A[6]), .A2(B[6]), .ZN(n48) );
  NAND2_X1 U162 ( .A1(A[8]), .A2(B[8]), .ZN(n40) );
  NAND2_X1 U163 ( .A1(A[11]), .A2(B[11]), .ZN(n27) );
  NAND2_X1 U164 ( .A1(A[9]), .A2(B[9]), .ZN(n35) );
  NAND2_X1 U165 ( .A1(A[13]), .A2(B[13]), .ZN(n19) );
  NAND2_X1 U166 ( .A1(A[7]), .A2(B[7]), .ZN(n43) );
  NOR2_X1 U167 ( .A1(A[3]), .A2(B[3]), .ZN(n65) );
  NAND2_X1 U168 ( .A1(B[2]), .A2(A[2]), .ZN(n69) );
  NOR2_X1 U169 ( .A1(A[11]), .A2(B[11]), .ZN(n26) );
  NOR2_X1 U170 ( .A1(A[9]), .A2(B[9]), .ZN(n34) );
  NOR2_X1 U171 ( .A1(A[13]), .A2(B[13]), .ZN(n18) );
  NOR2_X1 U172 ( .A1(A[7]), .A2(B[7]), .ZN(n42) );
  OR2_X1 U173 ( .A1(A[10]), .A2(B[10]), .ZN(n162) );
  OR2_X1 U174 ( .A1(A[8]), .A2(B[8]), .ZN(n163) );
  OR2_X1 U175 ( .A1(A[12]), .A2(B[12]), .ZN(n164) );
  AOI21_X1 U176 ( .B1(n63), .B2(n71), .A(n64), .ZN(n62) );
  AOI21_X1 U177 ( .B1(n161), .B2(n165), .A(n53), .ZN(n51) );
  AOI21_X1 U178 ( .B1(n153), .B2(n157), .A(n46), .ZN(n44) );
  OAI21_X1 U179 ( .B1(n62), .B2(n50), .A(n51), .ZN(n49) );
  AOI21_X1 U180 ( .B1(n151), .B2(n162), .A(n30), .ZN(n28) );
  CLKBUF_X1 U181 ( .A(n75), .Z(n166) );
  XNOR2_X1 U182 ( .A(n16), .B(n156), .ZN(SUM[15]) );
  CLKBUF_X1 U183 ( .A(n41), .Z(n167) );
  AOI21_X1 U184 ( .B1(n167), .B2(n163), .A(n38), .ZN(n168) );
  OAI21_X1 U185 ( .B1(n154), .B2(n42), .A(n43), .ZN(n41) );
  AOI21_X1 U186 ( .B1(n41), .B2(n163), .A(n38), .ZN(n36) );
  OAI21_X1 U187 ( .B1(n70), .B2(n68), .A(n145), .ZN(n67) );
  NAND2_X1 U188 ( .A1(n87), .A2(n145), .ZN(n13) );
  OAI21_X1 U189 ( .B1(n36), .B2(n34), .A(n35), .ZN(n33) );
  XNOR2_X1 U190 ( .A(n167), .B(n7), .ZN(SUM[8]) );
  NAND2_X1 U191 ( .A1(A[3]), .A2(B[3]), .ZN(n66) );
  XOR2_X1 U192 ( .A(n44), .B(n8), .Z(SUM[7]) );
  XNOR2_X1 U193 ( .A(n153), .B(n9), .ZN(SUM[6]) );
  XNOR2_X1 U194 ( .A(n149), .B(n3), .ZN(SUM[12]) );
  NAND2_X1 U195 ( .A1(A[5]), .A2(B[5]), .ZN(n55) );
  INV_X1 U196 ( .A(n150), .ZN(n61) );
  OAI21_X1 U197 ( .B1(n155), .B2(n26), .A(n27), .ZN(n25) );
  XNOR2_X1 U198 ( .A(n151), .B(n5), .ZN(SUM[10]) );
  XOR2_X1 U199 ( .A(n28), .B(n4), .Z(SUM[11]) );
  XOR2_X1 U200 ( .A(n168), .B(n6), .Z(SUM[9]) );
  NAND2_X1 U201 ( .A1(A[1]), .A2(B[1]), .ZN(n73) );
  NOR2_X1 U202 ( .A1(A[1]), .A2(B[1]), .ZN(n72) );
  XOR2_X1 U203 ( .A(n152), .B(n2), .Z(SUM[13]) );
  OAI21_X1 U204 ( .B1(n20), .B2(n18), .A(n19), .ZN(n17) );
  AOI21_X1 U205 ( .B1(n25), .B2(n164), .A(n22), .ZN(n20) );
  XOR2_X1 U206 ( .A(n14), .B(n166), .Z(SUM[1]) );
  OAI21_X1 U207 ( .B1(n72), .B2(n75), .A(n73), .ZN(n71) );
  NAND2_X1 U208 ( .A1(A[0]), .A2(B[0]), .ZN(n75) );
  INV_X1 U209 ( .A(n158), .ZN(n86) );
  NOR2_X1 U210 ( .A1(n68), .A2(n158), .ZN(n63) );
  OAI21_X1 U211 ( .B1(n65), .B2(n69), .A(n66), .ZN(n64) );
endmodule


module mvm3_part2 ( clk, reset, s_valid, m_ready, data_in, m_valid, s_ready, 
        data_out );
  input [7:0] data_in;
  output [15:0] data_out;
  input clk, reset, s_valid, m_ready;
  output m_valid, s_ready;
  wire   wr_en_m, wr_en_x, wr_en_b, \next_state[2] , N75, N76, N77, N78, N79,
         N80, store_complete, N83, N84, N85, \m_ptr[0] , valid_in, clear_mac,
         N167, N168, N169, N176, N177, N178, N179, N205, N229, N0, N1,
         valid_out, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265,
         N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, N276,
         N277, N278, N279, N280, N281, N282, N283, N284, N285, N286, N287, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n118, n119,
         n120, n121, n123, n124, n125, n128, n129, n131, n132, n137, n138,
         n139, n141, n142, n143, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n201, n202, n203, n204, n205, n229, n230, n231, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n299, n300, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         \rem_270/u_div/PartRem[3][2] , \rem_270/u_div/PartRem[3][1] ,
         \rem_270/u_div/PartRem[2][2] , \rem_270/u_div/PartRem[2][1] ,
         \rem_270/u_div/PartRem[1][2] , \rem_270/u_div/PartRem[1][1] ,
         \rem_270/u_div/SumTmp[3][1] , \rem_270/u_div/SumTmp[2][1] ,
         \rem_270/u_div/SumTmp[1][1] , \rem_270/u_div/SumTmp[0][1] ,
         \rem_270/quotient[3] , n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520;
  wire   [7:0] in_m;
  wire   [3:0] addr_m;
  wire   [7:0] in_x;
  wire   [1:0] addr_x;
  wire   [7:0] in_b;
  wire   [1:0] addr_b;
  wire   [2:0] state;
  wire   [3:0] in_ptr;
  wire   [2:0] load_ptr;
  wire   [3:0] out_ctr;
  wire   [1:0] out_ptr;
  wire   [15:0] f;
  wire   [4:2] \r484/carry ;
  wire   [4:2] \r482/carry ;

  DFF_X1 \out_ctr_reg[3]  ( .D(n488), .CK(clk), .Q(out_ctr[3]), .QN(n143) );
  DFF_X1 \out_ctr_reg[0]  ( .D(n489), .CK(clk), .Q(out_ctr[0]), .QN(n146) );
  DFF_X1 \out_ctr_reg[1]  ( .D(n490), .CK(clk), .Q(out_ctr[1]), .QN(n398) );
  DFF_X1 \out_ctr_reg[2]  ( .D(n491), .CK(clk), .Q(out_ctr[2]), .QN(n399) );
  DFF_X1 out_valid_reg ( .D(n373), .CK(clk), .QN(n128) );
  DFF_X1 \state_reg[2]  ( .D(n372), .CK(clk), .Q(state[2]), .QN(n118) );
  DFF_X1 \in_ptr_reg[3]  ( .D(n364), .CK(clk), .Q(in_ptr[3]), .QN(n132) );
  DFF_X1 \in_ptr_reg[0]  ( .D(n363), .CK(clk), .Q(in_ptr[0]), .QN(n139) );
  DFF_X1 \in_ptr_reg[1]  ( .D(n362), .CK(clk), .Q(in_ptr[1]), .QN(n138) );
  DFF_X1 \in_ptr_reg[2]  ( .D(n361), .CK(clk), .Q(in_ptr[2]), .QN(n137) );
  DFF_X1 s_ready_reg ( .D(n360), .CK(clk), .Q(s_ready), .QN(n125) );
  DFF_X1 \load_ptr_reg[0]  ( .D(n368), .CK(clk), .Q(load_ptr[0]), .QN(n124) );
  DFF_X1 \load_ptr_reg[1]  ( .D(n367), .CK(clk), .Q(load_ptr[1]), .QN(n123) );
  DFF_X1 \load_ptr_reg[2]  ( .D(n369), .CK(clk), .Q(load_ptr[2]), .QN(n121) );
  DFF_X1 \addr_b_reg[0]  ( .D(n358), .CK(clk), .Q(addr_b[0]), .QN(n149) );
  DFF_X1 \addr_b_reg[1]  ( .D(n359), .CK(clk), .Q(addr_b[1]), .QN(n148) );
  DFF_X1 \m_ptr_reg[1]  ( .D(n366), .CK(clk), .QN(n141) );
  DFF_X1 \m_ptr_reg[0]  ( .D(n365), .CK(clk), .Q(\m_ptr[0] ), .QN(n142) );
  DFF_X1 \addr_x_reg[1]  ( .D(n356), .CK(clk), .Q(addr_x[1]), .QN(n147) );
  DFF_X1 \acc_buff_reg[0][0]  ( .D(n353), .CK(clk), .QN(n197) );
  DFF_X1 \acc_buff_reg[2][0]  ( .D(n321), .CK(clk), .QN(n165) );
  DFF_X1 \acc_buff_reg[1][0]  ( .D(n337), .CK(clk), .QN(n181) );
  DFF_X1 \acc_buff_reg[2][1]  ( .D(n320), .CK(clk), .QN(n164) );
  DFF_X1 \acc_buff_reg[1][1]  ( .D(n336), .CK(clk), .QN(n180) );
  DFF_X1 \acc_buff_reg[0][1]  ( .D(n352), .CK(clk), .QN(n196) );
  DFF_X1 \acc_buff_reg[2][2]  ( .D(n319), .CK(clk), .QN(n163) );
  DFF_X1 \acc_buff_reg[1][2]  ( .D(n335), .CK(clk), .QN(n179) );
  DFF_X1 \acc_buff_reg[0][2]  ( .D(n351), .CK(clk), .QN(n195) );
  DFF_X1 \acc_buff_reg[2][3]  ( .D(n318), .CK(clk), .QN(n162) );
  DFF_X1 \acc_buff_reg[1][3]  ( .D(n334), .CK(clk), .QN(n178) );
  DFF_X1 \acc_buff_reg[0][3]  ( .D(n350), .CK(clk), .QN(n194) );
  DFF_X1 \acc_buff_reg[2][4]  ( .D(n317), .CK(clk), .QN(n161) );
  DFF_X1 \acc_buff_reg[1][4]  ( .D(n333), .CK(clk), .QN(n177) );
  DFF_X1 \acc_buff_reg[0][4]  ( .D(n349), .CK(clk), .QN(n193) );
  DFF_X1 \acc_buff_reg[2][5]  ( .D(n316), .CK(clk), .QN(n160) );
  DFF_X1 \acc_buff_reg[1][5]  ( .D(n332), .CK(clk), .QN(n176) );
  DFF_X1 \acc_buff_reg[0][5]  ( .D(n348), .CK(clk), .QN(n192) );
  DFF_X1 \acc_buff_reg[2][6]  ( .D(n315), .CK(clk), .QN(n159) );
  DFF_X1 \acc_buff_reg[1][6]  ( .D(n331), .CK(clk), .QN(n175) );
  DFF_X1 \acc_buff_reg[0][6]  ( .D(n347), .CK(clk), .QN(n191) );
  DFF_X1 \acc_buff_reg[2][7]  ( .D(n314), .CK(clk), .QN(n158) );
  DFF_X1 \acc_buff_reg[1][7]  ( .D(n330), .CK(clk), .QN(n174) );
  DFF_X1 \acc_buff_reg[0][7]  ( .D(n346), .CK(clk), .QN(n190) );
  DFF_X1 \acc_buff_reg[2][8]  ( .D(n313), .CK(clk), .QN(n157) );
  DFF_X1 \acc_buff_reg[1][8]  ( .D(n329), .CK(clk), .QN(n173) );
  DFF_X1 \acc_buff_reg[0][8]  ( .D(n345), .CK(clk), .QN(n189) );
  DFF_X1 \acc_buff_reg[2][9]  ( .D(n312), .CK(clk), .QN(n156) );
  DFF_X1 \acc_buff_reg[1][9]  ( .D(n328), .CK(clk), .QN(n172) );
  DFF_X1 \acc_buff_reg[0][9]  ( .D(n344), .CK(clk), .QN(n188) );
  DFF_X1 \acc_buff_reg[2][10]  ( .D(n311), .CK(clk), .QN(n155) );
  DFF_X1 \acc_buff_reg[1][10]  ( .D(n327), .CK(clk), .QN(n171) );
  DFF_X1 \acc_buff_reg[0][10]  ( .D(n343), .CK(clk), .QN(n187) );
  DFF_X1 \acc_buff_reg[2][11]  ( .D(n310), .CK(clk), .QN(n154) );
  DFF_X1 \acc_buff_reg[1][11]  ( .D(n326), .CK(clk), .QN(n170) );
  DFF_X1 \acc_buff_reg[0][11]  ( .D(n342), .CK(clk), .QN(n186) );
  DFF_X1 \acc_buff_reg[2][12]  ( .D(n309), .CK(clk), .QN(n153) );
  DFF_X1 \acc_buff_reg[1][12]  ( .D(n325), .CK(clk), .QN(n169) );
  DFF_X1 \acc_buff_reg[0][12]  ( .D(n341), .CK(clk), .QN(n185) );
  DFF_X1 \acc_buff_reg[2][13]  ( .D(n308), .CK(clk), .QN(n152) );
  DFF_X1 \acc_buff_reg[1][13]  ( .D(n324), .CK(clk), .QN(n168) );
  DFF_X1 \acc_buff_reg[0][13]  ( .D(n340), .CK(clk), .QN(n184) );
  DFF_X1 \acc_buff_reg[2][14]  ( .D(n307), .CK(clk), .QN(n151) );
  DFF_X1 \acc_buff_reg[1][14]  ( .D(n323), .CK(clk), .QN(n167) );
  DFF_X1 \acc_buff_reg[0][14]  ( .D(n339), .CK(clk), .QN(n183) );
  DFF_X1 \acc_buff_reg[2][15]  ( .D(n306), .CK(clk), .QN(n150) );
  DFF_X1 \acc_buff_reg[1][15]  ( .D(n322), .CK(clk), .QN(n166) );
  DFF_X1 \acc_buff_reg[0][15]  ( .D(n338), .CK(clk), .QN(n182) );
  DFF_X1 store_complete_reg ( .D(n305), .CK(clk), .Q(store_complete), .QN(n198) );
  XOR2_X1 U8 ( .A(state[0]), .B(state[1]), .Z(n56) );
  MUX2_X1 U12 ( .A(n57), .B(n54), .S(state[2]), .Z(n58) );
  MUX2_X1 U13 ( .A(N76), .B(N79), .S(state[1]), .Z(n59) );
  MUX2_X1 U15 ( .A(n60), .B(n55), .S(state[2]), .Z(n61) );
  NAND3_X1 U299 ( .A1(n240), .A2(n238), .A3(n241), .ZN(n239) );
  NAND3_X1 U300 ( .A1(n264), .A2(n149), .A3(n266), .ZN(n265) );
  NAND3_X1 U301 ( .A1(n266), .A2(n264), .A3(n268), .ZN(n267) );
  NAND3_X1 U302 ( .A1(n202), .A2(n203), .A3(n275), .ZN(n270) );
  NAND3_X1 U303 ( .A1(N168), .A2(N167), .A3(N169), .ZN(n278) );
  NAND3_X1 U304 ( .A1(n279), .A2(n496), .A3(n229), .ZN(n280) );
  NAND3_X1 U305 ( .A1(n288), .A2(n124), .A3(n287), .ZN(n289) );
  NAND3_X1 U306 ( .A1(n287), .A2(n288), .A3(n291), .ZN(n290) );
  NAND3_X1 U307 ( .A1(n507), .A2(n505), .A3(n292), .ZN(n288) );
  NAND3_X1 U308 ( .A1(n513), .A2(n475), .A3(n253), .ZN(n204) );
  NAND3_X1 U309 ( .A1(state[1]), .A2(n118), .A3(state[0]), .ZN(n281) );
  memory_WIDTH8_SIZE9_LOGSIZE4 memM ( .clk(clk), .data_in(data_in), .data_out(
        in_m), .addr(addr_m), .wr_en(wr_en_m) );
  memory_WIDTH8_SIZE3_LOGSIZE2_0 memx ( .clk(clk), .data_in(data_in), 
        .data_out(in_x), .addr(addr_x), .wr_en(wr_en_x) );
  memory_WIDTH8_SIZE3_LOGSIZE2_1 memb ( .clk(clk), .data_in(data_in), 
        .data_out(in_b), .addr(addr_b), .wr_en(wr_en_b) );
  part2_mac mac ( .clk(clk), .reset(clear_mac), .a(in_m), .b(in_x), .valid_in(
        valid_in), .f(f), .valid_out(valid_out) );
  MUX2_X1 \rem_270/u_div/u_mx_PartRem_0_0_0  ( .A(N176), .B(addr_m[0]), .S(
        n485), .Z(N0) );
  MUX2_X1 \rem_270/u_div/u_mx_PartRem_0_0_1  ( .A(
        \rem_270/u_div/PartRem[1][1] ), .B(\rem_270/u_div/SumTmp[0][1] ), .S(
        n485), .Z(N1) );
  MUX2_X1 \rem_270/u_div/u_mx_PartRem_0_1_0  ( .A(N177), .B(n480), .S(n484), 
        .Z(\rem_270/u_div/PartRem[1][1] ) );
  MUX2_X1 \rem_270/u_div/u_mx_PartRem_0_1_1  ( .A(
        \rem_270/u_div/PartRem[2][1] ), .B(\rem_270/u_div/SumTmp[1][1] ), .S(
        n484), .Z(\rem_270/u_div/PartRem[1][2] ) );
  MUX2_X1 \rem_270/u_div/u_mx_PartRem_0_2_0  ( .A(N178), .B(n481), .S(n483), 
        .Z(\rem_270/u_div/PartRem[2][1] ) );
  MUX2_X1 \rem_270/u_div/u_mx_PartRem_0_2_1  ( .A(
        \rem_270/u_div/PartRem[3][1] ), .B(\rem_270/u_div/SumTmp[2][1] ), .S(
        n483), .Z(\rem_270/u_div/PartRem[2][2] ) );
  MUX2_X1 \rem_270/u_div/u_mx_PartRem_0_3_0  ( .A(N179), .B(n482), .S(
        \rem_270/quotient[3] ), .Z(\rem_270/u_div/PartRem[3][1] ) );
  MUX2_X1 \rem_270/u_div/u_mx_PartRem_0_3_1  ( .A(N229), .B(
        \rem_270/u_div/SumTmp[3][1] ), .S(\rem_270/quotient[3] ), .Z(
        \rem_270/u_div/PartRem[3][2] ) );
  HA_X1 \r484/U1_1_1  ( .A(addr_m[1]), .B(addr_m[0]), .CO(\r484/carry [2]), 
        .S(N177) );
  HA_X1 \r484/U1_1_2  ( .A(addr_m[2]), .B(\r484/carry [2]), .CO(
        \r484/carry [3]), .S(N178) );
  HA_X1 \r484/U1_1_3  ( .A(addr_m[3]), .B(\r484/carry [3]), .CO(N229), .S(N179) );
  HA_X1 \r482/U1_1_1  ( .A(in_ptr[1]), .B(in_ptr[0]), .CO(\r482/carry [2]), 
        .S(N167) );
  HA_X1 \r482/U1_1_2  ( .A(in_ptr[2]), .B(\r482/carry [2]), .CO(
        \r482/carry [3]), .S(N168) );
  HA_X1 \r482/U1_1_3  ( .A(in_ptr[3]), .B(\r482/carry [3]), .CO(N205), .S(N169) );
  mvm3_part2_DW01_add_1 add_279 ( .A({N256, N257, N258, N259, N260, N261, N262, 
        N263, N264, N265, N266, N267, N268, N269, N270, N271}), .B(f), .CI(
        1'b0), .SUM({N287, N286, N285, N284, N283, N282, N281, N280, N279, 
        N278, N277, N276, N275, N274, N273, N272}) );
  DFF_X1 \out_ptr_reg[0]  ( .D(n354), .CK(clk), .Q(out_ptr[0]), .QN(n131) );
  DFF_X1 \state_reg[0]  ( .D(n370), .CK(clk), .Q(state[0]), .QN(n120) );
  DFF_X1 \state_reg[1]  ( .D(n371), .CK(clk), .Q(state[1]), .QN(n119) );
  DFF_X1 m_valid_reg ( .D(n503), .CK(clk), .Q(m_valid) );
  DFF_X1 valid_in_reg ( .D(n357), .CK(clk), .Q(valid_in) );
  DFF_X1 clear_mac_reg ( .D(n494), .CK(clk), .Q(clear_mac) );
  DFF_X1 \addr_m_reg[0]  ( .D(n500), .CK(clk), .Q(addr_m[0]), .QN(N176) );
  DFF_X1 \addr_m_reg[3]  ( .D(n497), .CK(clk), .Q(addr_m[3]) );
  DFF_X1 \addr_m_reg[2]  ( .D(n498), .CK(clk), .Q(addr_m[2]) );
  DFF_X1 \addr_m_reg[1]  ( .D(n499), .CK(clk), .Q(addr_m[1]) );
  DFF_X1 \addr_x_reg[0]  ( .D(n486), .CK(clk), .Q(addr_x[0]) );
  DFF_X1 \out_ptr_reg[1]  ( .D(n355), .CK(clk), .Q(out_ptr[1]), .QN(n129) );
  BUF_X2 U319 ( .A(n465), .Z(n397) );
  INV_X1 U320 ( .A(valid_out), .ZN(n492) );
  NOR3_X1 U321 ( .A1(n299), .A2(reset), .A3(n272), .ZN(n253) );
  AND2_X1 U322 ( .A1(n496), .A2(n476), .ZN(n383) );
  BUF_X1 U323 ( .A(n421), .Z(n391) );
  XNOR2_X1 U324 ( .A(n421), .B(out_ctr[1]), .ZN(n425) );
  AND2_X1 U325 ( .A1(out_ctr[2]), .A2(out_ctr[3]), .ZN(n384) );
  OR2_X1 U326 ( .A1(n399), .A2(n143), .ZN(n385) );
  OR2_X1 U327 ( .A1(n399), .A2(n143), .ZN(n419) );
  CLKBUF_X3 U328 ( .A(n466), .Z(n390) );
  OAI21_X1 U329 ( .B1(n425), .B2(n146), .A(n424), .ZN(n386) );
  INV_X1 U330 ( .A(n410), .ZN(n387) );
  NAND2_X2 U331 ( .A1(n458), .A2(n473), .ZN(n460) );
  OAI211_X2 U332 ( .C1(n433), .C2(n397), .A(n383), .B(n427), .ZN(n458) );
  NAND2_X2 U333 ( .A1(n461), .A2(n473), .ZN(n463) );
  OAI211_X2 U334 ( .C1(n464), .C2(n433), .A(n383), .B(n432), .ZN(n461) );
  OAI221_X4 U335 ( .B1(n390), .B2(n433), .C1(load_ptr[0]), .C2(n429), .A(n383), 
        .ZN(n467) );
  XNOR2_X1 U336 ( .A(n423), .B(n388), .ZN(n424) );
  NAND2_X1 U337 ( .A1(n387), .A2(n385), .ZN(n388) );
  BUF_X2 U338 ( .A(n466), .Z(n396) );
  OR2_X2 U339 ( .A1(n386), .A2(n391), .ZN(n465) );
  NAND2_X1 U340 ( .A1(n419), .A2(out_ctr[2]), .ZN(n389) );
  INV_X1 U341 ( .A(n275), .ZN(n509) );
  NOR2_X1 U342 ( .A1(n476), .A2(n255), .ZN(n275) );
  INV_X1 U343 ( .A(n252), .ZN(n502) );
  INV_X1 U344 ( .A(n204), .ZN(n504) );
  INV_X1 U345 ( .A(n293), .ZN(n513) );
  INV_X1 U346 ( .A(n241), .ZN(n520) );
  AOI21_X1 U347 ( .B1(n248), .B2(n505), .A(n501), .ZN(n257) );
  NAND4_X1 U348 ( .A1(n253), .A2(n281), .A3(n475), .A4(n509), .ZN(n279) );
  AOI22_X1 U349 ( .A1(n293), .A2(n496), .B1(n474), .B2(n273), .ZN(n292) );
  AOI22_X1 U350 ( .A1(n229), .A2(N205), .B1(n519), .B2(n231), .ZN(n254) );
  INV_X1 U351 ( .A(n262), .ZN(n519) );
  INV_X1 U352 ( .A(n478), .ZN(n484) );
  NOR2_X1 U353 ( .A1(n201), .A2(n202), .ZN(wr_en_m) );
  NAND4_X1 U354 ( .A1(n475), .A2(n514), .A3(n270), .A4(n271), .ZN(n264) );
  AOI221_X1 U355 ( .B1(n272), .B2(n273), .C1(N205), .C2(n229), .A(n274), .ZN(
        n271) );
  OAI211_X1 U356 ( .C1(n476), .C2(n510), .A(n253), .B(n254), .ZN(n252) );
  INV_X1 U357 ( .A(wr_en_x), .ZN(n510) );
  OAI211_X1 U358 ( .C1(n262), .C2(n475), .A(n513), .B(n253), .ZN(n283) );
  INV_X1 U359 ( .A(n261), .ZN(n501) );
  OAI211_X1 U360 ( .C1(n202), .C2(n509), .A(n253), .B(n254), .ZN(n261) );
  NOR2_X1 U361 ( .A1(n255), .A2(n203), .ZN(wr_en_x) );
  NAND2_X1 U362 ( .A1(n496), .A2(n281), .ZN(n274) );
  NAND2_X1 U363 ( .A1(n272), .A2(n496), .ZN(n269) );
  INV_X1 U364 ( .A(N177), .ZN(n480) );
  INV_X1 U365 ( .A(N178), .ZN(n481) );
  INV_X1 U366 ( .A(N179), .ZN(n482) );
  NAND2_X1 U367 ( .A1(n476), .A2(n281), .ZN(n293) );
  OR2_X1 U368 ( .A1(n201), .A2(n282), .ZN(n255) );
  AND3_X1 U369 ( .A1(n508), .A2(n203), .A3(n202), .ZN(wr_en_b) );
  INV_X1 U370 ( .A(n201), .ZN(n508) );
  INV_X1 U371 ( .A(n291), .ZN(n518) );
  NAND2_X1 U372 ( .A1(n294), .A2(n230), .ZN(n273) );
  INV_X1 U373 ( .A(n299), .ZN(n514) );
  XOR2_X1 U374 ( .A(n416), .B(n415), .Z(n392) );
  INV_X1 U375 ( .A(n477), .ZN(n483) );
  INV_X1 U376 ( .A(n240), .ZN(n507) );
  INV_X1 U377 ( .A(n244), .ZN(n506) );
  INV_X1 U378 ( .A(n479), .ZN(n485) );
  NOR3_X1 U379 ( .A1(state[0]), .A2(state[1]), .A3(n118), .ZN(n231) );
  NOR3_X1 U380 ( .A1(state[1]), .A2(state[2]), .A3(n120), .ZN(n229) );
  NOR3_X1 U381 ( .A1(state[0]), .A2(state[2]), .A3(n119), .ZN(n272) );
  NOR3_X1 U382 ( .A1(n139), .A2(n203), .A3(n138), .ZN(n282) );
  NOR3_X1 U383 ( .A1(state[1]), .A2(state[2]), .A3(state[0]), .ZN(n299) );
  NOR3_X1 U384 ( .A1(n124), .A2(load_ptr[2]), .A3(n123), .ZN(n291) );
  NOR3_X1 U385 ( .A1(n502), .A2(addr_x[0]), .A3(n248), .ZN(n249) );
  NOR3_X1 U386 ( .A1(state[1]), .A2(state[0]), .A3(N85), .ZN(n51) );
  OAI222_X1 U387 ( .A1(n181), .A2(n131), .B1(n197), .B2(n520), .C1(n165), .C2(
        n129), .ZN(data_out[0]) );
  OAI222_X1 U388 ( .A1(n180), .A2(n131), .B1(n196), .B2(n520), .C1(n164), .C2(
        n129), .ZN(data_out[1]) );
  OAI222_X1 U389 ( .A1(n179), .A2(n131), .B1(n195), .B2(n520), .C1(n163), .C2(
        n129), .ZN(data_out[2]) );
  OAI222_X1 U390 ( .A1(n178), .A2(n131), .B1(n194), .B2(n520), .C1(n162), .C2(
        n129), .ZN(data_out[3]) );
  OAI222_X1 U391 ( .A1(n177), .A2(n131), .B1(n193), .B2(n520), .C1(n161), .C2(
        n129), .ZN(data_out[4]) );
  OAI222_X1 U392 ( .A1(n176), .A2(n131), .B1(n192), .B2(n520), .C1(n160), .C2(
        n129), .ZN(data_out[5]) );
  OAI222_X1 U393 ( .A1(n175), .A2(n131), .B1(n191), .B2(n520), .C1(n159), .C2(
        n129), .ZN(data_out[6]) );
  OAI222_X1 U394 ( .A1(n174), .A2(n131), .B1(n190), .B2(n520), .C1(n158), .C2(
        n129), .ZN(data_out[7]) );
  OAI222_X1 U395 ( .A1(n173), .A2(n131), .B1(n189), .B2(n520), .C1(n157), .C2(
        n129), .ZN(data_out[8]) );
  OAI222_X1 U396 ( .A1(n172), .A2(n131), .B1(n188), .B2(n520), .C1(n156), .C2(
        n129), .ZN(data_out[9]) );
  NOR2_X1 U397 ( .A1(n514), .A2(reset), .ZN(n240) );
  AND2_X1 U398 ( .A1(n272), .A2(n121), .ZN(n287) );
  NOR2_X1 U399 ( .A1(n128), .A2(n507), .ZN(n244) );
  NOR2_X1 U400 ( .A1(n141), .A2(n142), .ZN(n262) );
  AOI21_X1 U401 ( .B1(n124), .B2(n287), .A(n493), .ZN(n285) );
  INV_X1 U402 ( .A(n288), .ZN(n493) );
  OAI22_X1 U403 ( .A1(n142), .A2(n283), .B1(\m_ptr[0] ), .B2(n505), .ZN(n365)
         );
  NAND2_X1 U404 ( .A1(in_b[7]), .A2(n428), .ZN(n443) );
  NAND2_X1 U405 ( .A1(in_b[7]), .A2(n430), .ZN(n444) );
  NAND2_X1 U406 ( .A1(in_b[7]), .A2(n434), .ZN(n445) );
  OAI22_X1 U407 ( .A1(n137), .A2(n279), .B1(n516), .B2(n280), .ZN(n361) );
  INV_X1 U408 ( .A(N168), .ZN(n516) );
  OAI22_X1 U409 ( .A1(n138), .A2(n279), .B1(n517), .B2(n280), .ZN(n362) );
  INV_X1 U410 ( .A(N167), .ZN(n517) );
  OAI22_X1 U411 ( .A1(n139), .A2(n279), .B1(in_ptr[0]), .B2(n280), .ZN(n363)
         );
  OAI22_X1 U412 ( .A1(n132), .A2(n279), .B1(n515), .B2(n280), .ZN(n364) );
  INV_X1 U413 ( .A(N169), .ZN(n515) );
  OAI22_X1 U414 ( .A1(n128), .A2(n495), .B1(n296), .B2(n297), .ZN(n373) );
  INV_X1 U415 ( .A(n296), .ZN(n495) );
  NOR2_X1 U416 ( .A1(n238), .A2(n229), .ZN(n296) );
  OAI22_X1 U417 ( .A1(n245), .A2(n147), .B1(n502), .B2(n246), .ZN(n356) );
  NOR2_X1 U418 ( .A1(n249), .A2(n502), .ZN(n245) );
  AOI22_X1 U419 ( .A1(n247), .A2(addr_x[0]), .B1(N1), .B2(n473), .ZN(n246) );
  NOR2_X1 U420 ( .A1(addr_x[1]), .A2(n248), .ZN(n247) );
  OAI22_X1 U421 ( .A1(n125), .A2(n204), .B1(n277), .B2(n248), .ZN(n360) );
  NOR4_X1 U422 ( .A1(n278), .A2(in_ptr[0]), .A3(N205), .A4(n255), .ZN(n277) );
  NAND2_X1 U423 ( .A1(in_ptr[3]), .A2(in_ptr[2]), .ZN(n203) );
  NOR2_X1 U424 ( .A1(out_ptr[0]), .A2(out_ptr[1]), .ZN(n241) );
  OAI21_X1 U425 ( .B1(load_ptr[2]), .B2(n269), .A(n248), .ZN(n266) );
  OAI21_X1 U426 ( .B1(N77), .B2(state[1]), .A(state[0]), .ZN(n52) );
  NOR2_X1 U427 ( .A1(n282), .A2(n118), .ZN(N77) );
  OAI21_X1 U428 ( .B1(n238), .B2(n129), .A(n242), .ZN(n355) );
  NAND4_X1 U429 ( .A1(out_ptr[0]), .A2(n240), .A3(n238), .A4(n129), .ZN(n242)
         );
  NAND2_X1 U430 ( .A1(n203), .A2(n276), .ZN(n202) );
  OAI21_X1 U431 ( .B1(in_ptr[0]), .B2(in_ptr[1]), .A(in_ptr[3]), .ZN(n276) );
  OAI21_X1 U432 ( .B1(n204), .B2(n198), .A(n205), .ZN(n305) );
  OAI21_X1 U433 ( .B1(n262), .B2(n505), .A(n263), .ZN(n357) );
  NAND2_X1 U434 ( .A1(valid_in), .A2(n504), .ZN(n263) );
  OAI21_X1 U435 ( .B1(n238), .B2(n131), .A(n239), .ZN(n354) );
  OAI21_X1 U436 ( .B1(n264), .B2(n148), .A(n267), .ZN(n359) );
  XNOR2_X1 U437 ( .A(n148), .B(addr_b[0]), .ZN(n268) );
  OAI21_X1 U438 ( .B1(n264), .B2(n149), .A(n265), .ZN(n358) );
  NOR2_X1 U439 ( .A1(n291), .A2(n118), .ZN(N80) );
  AOI21_X1 U440 ( .B1(N83), .B2(n119), .A(state[0]), .ZN(n54) );
  NAND2_X1 U441 ( .A1(s_valid), .A2(s_ready), .ZN(n201) );
  NAND2_X1 U442 ( .A1(n123), .A2(n124), .ZN(n294) );
  OR3_X1 U443 ( .A1(N205), .A2(reset), .A3(n476), .ZN(n248) );
  OAI21_X1 U444 ( .B1(n285), .B2(n123), .A(n286), .ZN(n367) );
  NAND4_X1 U445 ( .A1(n287), .A2(load_ptr[0]), .A3(n288), .A4(n123), .ZN(n286)
         );
  OR3_X1 U446 ( .A1(n300), .A2(n231), .A3(n274), .ZN(n238) );
  AND3_X1 U447 ( .A1(m_ready), .A2(n299), .A3(m_valid), .ZN(n300) );
  OAI21_X1 U448 ( .B1(n285), .B2(n121), .A(n290), .ZN(n369) );
  NAND2_X1 U449 ( .A1(n294), .A2(n121), .ZN(n230) );
  AND2_X1 U450 ( .A1(n394), .A2(n418), .ZN(n393) );
  NOR2_X1 U451 ( .A1(n492), .A2(n402), .ZN(n394) );
  NOR2_X1 U452 ( .A1(n244), .A2(n295), .ZN(n370) );
  NOR2_X1 U453 ( .A1(n511), .A2(reset), .ZN(n295) );
  INV_X1 U454 ( .A(n58), .ZN(n511) );
  OAI22_X1 U455 ( .A1(n284), .A2(n141), .B1(n505), .B2(n142), .ZN(n366) );
  AND2_X1 U456 ( .A1(n505), .A2(n283), .ZN(n284) );
  INV_X1 U457 ( .A(in_b[6]), .ZN(n487) );
  INV_X1 U458 ( .A(n258), .ZN(n498) );
  AOI22_X1 U459 ( .A1(N178), .A2(n257), .B1(addr_m[2]), .B2(n501), .ZN(n258)
         );
  OAI22_X1 U460 ( .A1(N78), .A2(n119), .B1(n50), .B2(n120), .ZN(n57) );
  NAND2_X1 U461 ( .A1(n120), .A2(n518), .ZN(N78) );
  AND2_X1 U462 ( .A1(N75), .A2(n119), .ZN(n50) );
  NOR2_X1 U463 ( .A1(n282), .A2(n120), .ZN(N75) );
  NAND2_X1 U464 ( .A1(n59), .A2(n56), .ZN(n60) );
  NAND2_X1 U465 ( .A1(n119), .A2(n518), .ZN(N79) );
  INV_X1 U466 ( .A(n260), .ZN(n500) );
  AOI22_X1 U467 ( .A1(N176), .A2(n257), .B1(addr_m[0]), .B2(n501), .ZN(n260)
         );
  OAI222_X1 U468 ( .A1(n166), .A2(n390), .B1(n182), .B2(n397), .C1(n150), .C2(
        n464), .ZN(N256) );
  INV_X1 U469 ( .A(n259), .ZN(n499) );
  AOI22_X1 U470 ( .A1(N177), .A2(n257), .B1(addr_m[1]), .B2(n501), .ZN(n259)
         );
  INV_X1 U471 ( .A(n250), .ZN(n486) );
  AOI211_X1 U472 ( .C1(addr_x[0]), .C2(n502), .A(n251), .B(n249), .ZN(n250) );
  AND3_X1 U473 ( .A1(n473), .A2(n252), .A3(N0), .ZN(n251) );
  INV_X1 U474 ( .A(n256), .ZN(n497) );
  AOI22_X1 U475 ( .A1(N179), .A2(n257), .B1(addr_m[3]), .B2(n501), .ZN(n256)
         );
  AND3_X1 U476 ( .A1(n506), .A2(n496), .A3(\next_state[2] ), .ZN(n372) );
  OAI211_X1 U477 ( .C1(n118), .C2(n51), .A(n52), .B(n53), .ZN(\next_state[2] )
         );
  NAND2_X1 U478 ( .A1(N80), .A2(state[1]), .ZN(n53) );
  AND3_X1 U479 ( .A1(n506), .A2(n496), .A3(n512), .ZN(n371) );
  INV_X1 U480 ( .A(n61), .ZN(n512) );
  AOI21_X1 U481 ( .B1(N84), .B2(n120), .A(state[1]), .ZN(n55) );
  OR2_X1 U482 ( .A1(state[1]), .A2(n282), .ZN(N76) );
  INV_X1 U483 ( .A(n304), .ZN(n494) );
  AOI21_X1 U484 ( .B1(clear_mac), .B2(n504), .A(n274), .ZN(n304) );
  INV_X1 U485 ( .A(n243), .ZN(n503) );
  AOI21_X1 U486 ( .B1(n504), .B2(m_valid), .A(n244), .ZN(n243) );
  INV_X1 U487 ( .A(reset), .ZN(n496) );
  INV_X1 U488 ( .A(n391), .ZN(n464) );
  OAI22_X1 U489 ( .A1(n384), .A2(n420), .B1(n422), .B2(n398), .ZN(n421) );
  OAI22_X1 U490 ( .A1(n384), .A2(n420), .B1(n389), .B2(n398), .ZN(n395) );
  INV_X1 U491 ( .A(n386), .ZN(n466) );
  INV_X1 U492 ( .A(n231), .ZN(n475) );
  NAND2_X1 U493 ( .A1(n231), .A2(n496), .ZN(n505) );
  OAI21_X1 U494 ( .B1(n124), .B2(n288), .A(n289), .ZN(n368) );
  INV_X1 U495 ( .A(out_ctr[2]), .ZN(n410) );
  NAND2_X1 U496 ( .A1(n410), .A2(n398), .ZN(n400) );
  OR3_X1 U497 ( .A1(n420), .A2(n146), .A3(n400), .ZN(n404) );
  INV_X1 U498 ( .A(n505), .ZN(n473) );
  INV_X1 U499 ( .A(n229), .ZN(n476) );
  INV_X1 U500 ( .A(n404), .ZN(n472) );
  INV_X1 U501 ( .A(n400), .ZN(n401) );
  INV_X1 U502 ( .A(out_ctr[3]), .ZN(n420) );
  AOI21_X1 U503 ( .B1(n401), .B2(n146), .A(n420), .ZN(n402) );
  OAI21_X1 U504 ( .B1(n472), .B2(n394), .A(n231), .ZN(n403) );
  NAND3_X1 U505 ( .A1(n253), .A2(n476), .A3(n403), .ZN(n411) );
  NAND3_X1 U506 ( .A1(n404), .A2(n473), .A3(n411), .ZN(n412) );
  NAND2_X1 U507 ( .A1(out_ctr[1]), .A2(out_ctr[0]), .ZN(n409) );
  INV_X1 U508 ( .A(n409), .ZN(n405) );
  NAND2_X1 U509 ( .A1(n387), .A2(n405), .ZN(n406) );
  XOR2_X1 U510 ( .A(n406), .B(out_ctr[3]), .Z(n413) );
  OAI22_X1 U511 ( .A1(n412), .A2(n413), .B1(n420), .B2(n411), .ZN(n488) );
  INV_X1 U512 ( .A(n412), .ZN(n408) );
  INV_X1 U513 ( .A(n411), .ZN(n407) );
  MUX2_X1 U514 ( .A(n408), .B(n407), .S(out_ctr[0]), .Z(n489) );
  XOR2_X1 U515 ( .A(n409), .B(n387), .Z(n414) );
  OAI22_X1 U516 ( .A1(n414), .A2(n412), .B1(n410), .B2(n411), .ZN(n491) );
  XOR2_X1 U517 ( .A(n146), .B(out_ctr[1]), .Z(n415) );
  OAI22_X1 U518 ( .A1(n415), .A2(n412), .B1(n398), .B2(n411), .ZN(n490) );
  OAI21_X1 U519 ( .B1(n415), .B2(n414), .A(n413), .ZN(n416) );
  NAND3_X1 U520 ( .A1(n392), .A2(n416), .A3(out_ctr[0]), .ZN(n417) );
  OAI21_X1 U521 ( .B1(out_ctr[0]), .B2(n392), .A(n417), .ZN(n418) );
  NAND2_X1 U522 ( .A1(n393), .A2(n231), .ZN(n433) );
  NAND2_X1 U523 ( .A1(n385), .A2(out_ctr[2]), .ZN(n422) );
  NAND2_X1 U524 ( .A1(n395), .A2(out_ctr[1]), .ZN(n423) );
  INV_X1 U525 ( .A(n230), .ZN(n426) );
  NAND2_X1 U526 ( .A1(n272), .A2(n426), .ZN(n429) );
  INV_X1 U527 ( .A(n429), .ZN(n431) );
  NAND3_X1 U528 ( .A1(load_ptr[0]), .A2(n431), .A3(n123), .ZN(n427) );
  INV_X1 U529 ( .A(N287), .ZN(n435) );
  INV_X1 U530 ( .A(n269), .ZN(n474) );
  NAND2_X1 U531 ( .A1(n458), .A2(n474), .ZN(n459) );
  INV_X1 U532 ( .A(n459), .ZN(n428) );
  OAI221_X1 U533 ( .B1(n460), .B2(n435), .C1(n182), .C2(n458), .A(n443), .ZN(
        n338) );
  NAND2_X1 U534 ( .A1(n467), .A2(n473), .ZN(n471) );
  NAND2_X1 U535 ( .A1(n467), .A2(n474), .ZN(n469) );
  INV_X1 U536 ( .A(n469), .ZN(n430) );
  OAI221_X1 U537 ( .B1(n435), .B2(n471), .C1(n166), .C2(n467), .A(n444), .ZN(
        n322) );
  NAND3_X1 U538 ( .A1(load_ptr[1]), .A2(load_ptr[0]), .A3(n431), .ZN(n432) );
  NAND2_X1 U539 ( .A1(n461), .A2(n474), .ZN(n462) );
  INV_X1 U540 ( .A(n462), .ZN(n434) );
  OAI221_X1 U541 ( .B1(n463), .B2(n435), .C1(n150), .C2(n461), .A(n445), .ZN(
        n306) );
  INV_X1 U542 ( .A(N286), .ZN(n436) );
  OAI221_X1 U543 ( .B1(n460), .B2(n436), .C1(n183), .C2(n458), .A(n443), .ZN(
        n339) );
  OAI221_X1 U544 ( .B1(n471), .B2(n436), .C1(n167), .C2(n467), .A(n444), .ZN(
        n323) );
  OAI221_X1 U545 ( .B1(n463), .B2(n436), .C1(n151), .C2(n461), .A(n445), .ZN(
        n307) );
  OAI222_X1 U546 ( .A1(n167), .A2(n390), .B1(n183), .B2(n397), .C1(n151), .C2(
        n464), .ZN(N257) );
  INV_X1 U547 ( .A(N285), .ZN(n437) );
  OAI221_X1 U548 ( .B1(n460), .B2(n437), .C1(n184), .C2(n458), .A(n443), .ZN(
        n340) );
  OAI221_X1 U549 ( .B1(n471), .B2(n437), .C1(n168), .C2(n467), .A(n444), .ZN(
        n324) );
  OAI221_X1 U550 ( .B1(n463), .B2(n437), .C1(n152), .C2(n461), .A(n445), .ZN(
        n308) );
  OAI222_X1 U551 ( .A1(n168), .A2(n390), .B1(n184), .B2(n397), .C1(n152), .C2(
        n464), .ZN(N258) );
  INV_X1 U552 ( .A(N284), .ZN(n438) );
  OAI221_X1 U553 ( .B1(n460), .B2(n438), .C1(n185), .C2(n458), .A(n443), .ZN(
        n341) );
  OAI221_X1 U554 ( .B1(n471), .B2(n438), .C1(n169), .C2(n467), .A(n444), .ZN(
        n325) );
  OAI221_X1 U555 ( .B1(n463), .B2(n438), .C1(n153), .C2(n461), .A(n445), .ZN(
        n309) );
  OAI222_X1 U556 ( .A1(n169), .A2(n390), .B1(n185), .B2(n397), .C1(n153), .C2(
        n464), .ZN(N259) );
  INV_X1 U557 ( .A(N283), .ZN(n439) );
  OAI221_X1 U558 ( .B1(n460), .B2(n439), .C1(n186), .C2(n458), .A(n443), .ZN(
        n342) );
  OAI221_X1 U559 ( .B1(n471), .B2(n439), .C1(n170), .C2(n467), .A(n444), .ZN(
        n326) );
  OAI221_X1 U560 ( .B1(n463), .B2(n439), .C1(n154), .C2(n461), .A(n445), .ZN(
        n310) );
  OAI222_X1 U561 ( .A1(n170), .A2(n390), .B1(n186), .B2(n397), .C1(n154), .C2(
        n464), .ZN(N260) );
  INV_X1 U562 ( .A(N282), .ZN(n440) );
  OAI221_X1 U563 ( .B1(n460), .B2(n440), .C1(n187), .C2(n458), .A(n443), .ZN(
        n343) );
  OAI221_X1 U564 ( .B1(n471), .B2(n440), .C1(n171), .C2(n467), .A(n444), .ZN(
        n327) );
  OAI221_X1 U565 ( .B1(n463), .B2(n440), .C1(n155), .C2(n461), .A(n445), .ZN(
        n311) );
  OAI222_X1 U566 ( .A1(n171), .A2(n390), .B1(n187), .B2(n397), .C1(n155), .C2(
        n464), .ZN(N261) );
  INV_X1 U567 ( .A(N281), .ZN(n441) );
  OAI221_X1 U568 ( .B1(n460), .B2(n441), .C1(n188), .C2(n458), .A(n443), .ZN(
        n344) );
  OAI221_X1 U569 ( .B1(n471), .B2(n441), .C1(n172), .C2(n467), .A(n444), .ZN(
        n328) );
  OAI221_X1 U570 ( .B1(n463), .B2(n441), .C1(n156), .C2(n461), .A(n445), .ZN(
        n312) );
  OAI222_X1 U571 ( .A1(n172), .A2(n390), .B1(n188), .B2(n397), .C1(n156), .C2(
        n464), .ZN(N262) );
  INV_X1 U572 ( .A(N280), .ZN(n442) );
  OAI221_X1 U573 ( .B1(n460), .B2(n442), .C1(n189), .C2(n458), .A(n443), .ZN(
        n345) );
  OAI221_X1 U574 ( .B1(n471), .B2(n442), .C1(n173), .C2(n467), .A(n444), .ZN(
        n329) );
  OAI221_X1 U575 ( .B1(n463), .B2(n442), .C1(n157), .C2(n461), .A(n445), .ZN(
        n313) );
  OAI222_X1 U576 ( .A1(n173), .A2(n390), .B1(n189), .B2(n397), .C1(n157), .C2(
        n464), .ZN(N263) );
  INV_X1 U577 ( .A(N279), .ZN(n446) );
  OAI221_X1 U578 ( .B1(n460), .B2(n446), .C1(n190), .C2(n458), .A(n443), .ZN(
        n346) );
  OAI221_X1 U579 ( .B1(n471), .B2(n446), .C1(n174), .C2(n467), .A(n444), .ZN(
        n330) );
  OAI221_X1 U580 ( .B1(n463), .B2(n446), .C1(n158), .C2(n461), .A(n445), .ZN(
        n314) );
  OAI222_X1 U581 ( .A1(n174), .A2(n390), .B1(n190), .B2(n397), .C1(n158), .C2(
        n464), .ZN(N264) );
  INV_X1 U582 ( .A(N278), .ZN(n447) );
  OAI222_X1 U583 ( .A1(n460), .A2(n447), .B1(n487), .B2(n459), .C1(n191), .C2(
        n458), .ZN(n347) );
  OAI222_X1 U584 ( .A1(n471), .A2(n447), .B1(n487), .B2(n469), .C1(n175), .C2(
        n467), .ZN(n331) );
  OAI222_X1 U585 ( .A1(n463), .A2(n447), .B1(n487), .B2(n462), .C1(n159), .C2(
        n461), .ZN(n315) );
  OAI222_X1 U586 ( .A1(n175), .A2(n390), .B1(n191), .B2(n397), .C1(n159), .C2(
        n464), .ZN(N265) );
  INV_X1 U587 ( .A(N277), .ZN(n449) );
  INV_X1 U588 ( .A(in_b[5]), .ZN(n448) );
  OAI222_X1 U589 ( .A1(n460), .A2(n449), .B1(n459), .B2(n448), .C1(n192), .C2(
        n458), .ZN(n348) );
  OAI222_X1 U590 ( .A1(n471), .A2(n449), .B1(n469), .B2(n448), .C1(n176), .C2(
        n467), .ZN(n332) );
  OAI222_X1 U591 ( .A1(n463), .A2(n449), .B1(n462), .B2(n448), .C1(n160), .C2(
        n461), .ZN(n316) );
  OAI222_X1 U592 ( .A1(n176), .A2(n396), .B1(n192), .B2(n465), .C1(n160), .C2(
        n464), .ZN(N266) );
  INV_X1 U593 ( .A(N276), .ZN(n451) );
  INV_X1 U594 ( .A(in_b[4]), .ZN(n450) );
  OAI222_X1 U595 ( .A1(n460), .A2(n451), .B1(n459), .B2(n450), .C1(n193), .C2(
        n458), .ZN(n349) );
  OAI222_X1 U596 ( .A1(n471), .A2(n451), .B1(n469), .B2(n450), .C1(n177), .C2(
        n467), .ZN(n333) );
  OAI222_X1 U597 ( .A1(n463), .A2(n451), .B1(n462), .B2(n450), .C1(n161), .C2(
        n461), .ZN(n317) );
  OAI222_X1 U598 ( .A1(n177), .A2(n390), .B1(n193), .B2(n465), .C1(n161), .C2(
        n464), .ZN(N267) );
  INV_X1 U599 ( .A(N275), .ZN(n453) );
  INV_X1 U600 ( .A(in_b[3]), .ZN(n452) );
  OAI222_X1 U601 ( .A1(n460), .A2(n453), .B1(n459), .B2(n452), .C1(n194), .C2(
        n458), .ZN(n350) );
  OAI222_X1 U602 ( .A1(n471), .A2(n453), .B1(n469), .B2(n452), .C1(n178), .C2(
        n467), .ZN(n334) );
  OAI222_X1 U603 ( .A1(n463), .A2(n453), .B1(n462), .B2(n452), .C1(n162), .C2(
        n461), .ZN(n318) );
  OAI222_X1 U604 ( .A1(n178), .A2(n396), .B1(n194), .B2(n465), .C1(n162), .C2(
        n464), .ZN(N268) );
  INV_X1 U605 ( .A(N274), .ZN(n455) );
  INV_X1 U606 ( .A(in_b[2]), .ZN(n454) );
  OAI222_X1 U607 ( .A1(n460), .A2(n455), .B1(n459), .B2(n454), .C1(n195), .C2(
        n458), .ZN(n351) );
  OAI222_X1 U608 ( .A1(n471), .A2(n455), .B1(n469), .B2(n454), .C1(n179), .C2(
        n467), .ZN(n335) );
  OAI222_X1 U609 ( .A1(n463), .A2(n455), .B1(n462), .B2(n454), .C1(n163), .C2(
        n461), .ZN(n319) );
  OAI222_X1 U610 ( .A1(n179), .A2(n396), .B1(n195), .B2(n465), .C1(n163), .C2(
        n464), .ZN(N269) );
  INV_X1 U611 ( .A(N273), .ZN(n457) );
  INV_X1 U612 ( .A(in_b[1]), .ZN(n456) );
  OAI222_X1 U613 ( .A1(n460), .A2(n457), .B1(n459), .B2(n456), .C1(n196), .C2(
        n458), .ZN(n352) );
  OAI222_X1 U614 ( .A1(n471), .A2(n457), .B1(n469), .B2(n456), .C1(n180), .C2(
        n467), .ZN(n336) );
  OAI222_X1 U615 ( .A1(n463), .A2(n457), .B1(n462), .B2(n456), .C1(n164), .C2(
        n461), .ZN(n320) );
  OAI222_X1 U616 ( .A1(n180), .A2(n396), .B1(n196), .B2(n465), .C1(n164), .C2(
        n464), .ZN(N270) );
  INV_X1 U617 ( .A(N272), .ZN(n470) );
  INV_X1 U618 ( .A(in_b[0]), .ZN(n468) );
  OAI222_X1 U619 ( .A1(n470), .A2(n460), .B1(n468), .B2(n459), .C1(n197), .C2(
        n458), .ZN(n353) );
  OAI222_X1 U620 ( .A1(n470), .A2(n463), .B1(n468), .B2(n462), .C1(n165), .C2(
        n461), .ZN(n321) );
  OAI222_X1 U621 ( .A1(n181), .A2(n396), .B1(n197), .B2(n465), .C1(n165), .C2(
        n464), .ZN(N271) );
  OAI222_X1 U622 ( .A1(n471), .A2(n470), .B1(n469), .B2(n468), .C1(n181), .C2(
        n467), .ZN(n337) );
  AOI22_X1 U623 ( .A1(n472), .A2(n473), .B1(n240), .B2(n129), .ZN(n297) );
  NAND2_X1 U624 ( .A1(n473), .A2(n393), .ZN(n205) );
  NOR3_X1 U625 ( .A1(n118), .A2(store_complete), .A3(n472), .ZN(N85) );
  AOI21_X1 U626 ( .B1(n119), .B2(n198), .A(n472), .ZN(N84) );
  AOI21_X1 U627 ( .B1(n120), .B2(n198), .A(n472), .ZN(N83) );
  OAI222_X1 U628 ( .A1(n131), .A2(n171), .B1(n520), .B2(n187), .C1(n129), .C2(
        n155), .ZN(data_out[10]) );
  OAI222_X1 U629 ( .A1(n131), .A2(n170), .B1(n520), .B2(n186), .C1(n129), .C2(
        n154), .ZN(data_out[11]) );
  OAI222_X1 U630 ( .A1(n131), .A2(n169), .B1(n520), .B2(n185), .C1(n129), .C2(
        n153), .ZN(data_out[12]) );
  OAI222_X1 U631 ( .A1(n131), .A2(n168), .B1(n520), .B2(n184), .C1(n129), .C2(
        n152), .ZN(data_out[13]) );
  OAI222_X1 U632 ( .A1(n131), .A2(n167), .B1(n520), .B2(n183), .C1(n129), .C2(
        n151), .ZN(data_out[14]) );
  OAI222_X1 U633 ( .A1(n131), .A2(n166), .B1(n520), .B2(n182), .C1(n129), .C2(
        n150), .ZN(data_out[15]) );
  XOR2_X1 U634 ( .A(N179), .B(N229), .Z(\rem_270/u_div/SumTmp[3][1] ) );
  AND2_X1 U635 ( .A1(N179), .A2(N229), .ZN(\rem_270/quotient[3] ) );
  XOR2_X1 U636 ( .A(N178), .B(\rem_270/u_div/PartRem[3][1] ), .Z(
        \rem_270/u_div/SumTmp[2][1] ) );
  AOI21_X1 U637 ( .B1(N178), .B2(\rem_270/u_div/PartRem[3][1] ), .A(
        \rem_270/u_div/PartRem[3][2] ), .ZN(n477) );
  XOR2_X1 U638 ( .A(N177), .B(\rem_270/u_div/PartRem[2][1] ), .Z(
        \rem_270/u_div/SumTmp[1][1] ) );
  AOI21_X1 U639 ( .B1(N177), .B2(\rem_270/u_div/PartRem[2][1] ), .A(
        \rem_270/u_div/PartRem[2][2] ), .ZN(n478) );
  XOR2_X1 U640 ( .A(N176), .B(\rem_270/u_div/PartRem[1][1] ), .Z(
        \rem_270/u_div/SumTmp[0][1] ) );
  AOI21_X1 U641 ( .B1(N176), .B2(\rem_270/u_div/PartRem[1][1] ), .A(
        \rem_270/u_div/PartRem[1][2] ), .ZN(n479) );
endmodule

