
module part2_mac_DW01_add_1 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16, n17,
         n18, n19, n20, n22, n24, n25, n26, n27, n28, n30, n32, n33, n34, n35,
         n36, n38, n40, n41, n42, n43, n44, n46, n48, n49, n50, n51, n52, n54,
         n56, n57, n58, n59, n60, n62, n64, n65, n66, n67, n69, n70, n72, n74,
         n76, n78, n80, n82, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n154, n155, n156;

  FA_X1 U3 ( .A(A[14]), .B(B[14]), .CI(n17), .CO(n16), .S(SUM[14]) );
  AOI21_X1 U102 ( .B1(n49), .B2(n148), .A(n46), .ZN(n138) );
  CLKBUF_X1 U103 ( .A(n25), .Z(n139) );
  CLKBUF_X1 U104 ( .A(n33), .Z(n140) );
  CLKBUF_X1 U105 ( .A(n57), .Z(n141) );
  AOI21_X1 U106 ( .B1(n57), .B2(n149), .A(n54), .ZN(n142) );
  AOI21_X1 U107 ( .B1(n33), .B2(n151), .A(n30), .ZN(n143) );
  CLKBUF_X1 U108 ( .A(n41), .Z(n144) );
  AOI21_X1 U109 ( .B1(n41), .B2(n147), .A(n38), .ZN(n145) );
  CLKBUF_X1 U110 ( .A(n65), .Z(n146) );
  INV_X1 U111 ( .A(n40), .ZN(n38) );
  INV_X1 U112 ( .A(n32), .ZN(n30) );
  INV_X1 U113 ( .A(n48), .ZN(n46) );
  INV_X1 U114 ( .A(n56), .ZN(n54) );
  INV_X1 U115 ( .A(n24), .ZN(n22) );
  INV_X1 U116 ( .A(n18), .ZN(n70) );
  INV_X1 U117 ( .A(n26), .ZN(n72) );
  INV_X1 U118 ( .A(n34), .ZN(n74) );
  INV_X1 U119 ( .A(n42), .ZN(n76) );
  INV_X1 U120 ( .A(n50), .ZN(n78) );
  NAND2_X1 U121 ( .A1(n80), .A2(n59), .ZN(n12) );
  INV_X1 U122 ( .A(n58), .ZN(n80) );
  INV_X1 U123 ( .A(n64), .ZN(n62) );
  XOR2_X1 U124 ( .A(B[15]), .B(A[15]), .Z(n1) );
  NAND2_X1 U125 ( .A1(n78), .A2(n51), .ZN(n10) );
  NAND2_X1 U126 ( .A1(n74), .A2(n35), .ZN(n6) );
  NAND2_X1 U127 ( .A1(n76), .A2(n43), .ZN(n8) );
  NAND2_X1 U128 ( .A1(n149), .A2(n56), .ZN(n11) );
  NOR2_X1 U129 ( .A1(A[7]), .A2(B[7]), .ZN(n42) );
  NOR2_X1 U130 ( .A1(A[5]), .A2(B[5]), .ZN(n50) );
  NOR2_X1 U131 ( .A1(A[3]), .A2(B[3]), .ZN(n58) );
  NOR2_X1 U132 ( .A1(A[11]), .A2(B[11]), .ZN(n26) );
  NOR2_X1 U133 ( .A1(A[13]), .A2(B[13]), .ZN(n18) );
  NOR2_X1 U134 ( .A1(A[9]), .A2(B[9]), .ZN(n34) );
  NAND2_X1 U135 ( .A1(A[8]), .A2(B[8]), .ZN(n40) );
  NAND2_X1 U136 ( .A1(A[6]), .A2(B[6]), .ZN(n48) );
  NAND2_X1 U137 ( .A1(A[4]), .A2(B[4]), .ZN(n56) );
  NAND2_X1 U138 ( .A1(A[12]), .A2(B[12]), .ZN(n24) );
  NAND2_X1 U139 ( .A1(A[7]), .A2(B[7]), .ZN(n43) );
  NAND2_X1 U140 ( .A1(A[5]), .A2(B[5]), .ZN(n51) );
  NAND2_X1 U141 ( .A1(A[3]), .A2(B[3]), .ZN(n59) );
  NAND2_X1 U142 ( .A1(A[13]), .A2(B[13]), .ZN(n19) );
  NAND2_X1 U143 ( .A1(A[11]), .A2(B[11]), .ZN(n27) );
  NAND2_X1 U144 ( .A1(A[9]), .A2(B[9]), .ZN(n35) );
  OR2_X1 U145 ( .A1(A[8]), .A2(B[8]), .ZN(n147) );
  OR2_X1 U146 ( .A1(A[6]), .A2(B[6]), .ZN(n148) );
  OR2_X1 U147 ( .A1(A[4]), .A2(B[4]), .ZN(n149) );
  OR2_X1 U148 ( .A1(A[12]), .A2(B[12]), .ZN(n150) );
  OR2_X1 U149 ( .A1(A[10]), .A2(B[10]), .ZN(n151) );
  OR2_X1 U150 ( .A1(A[2]), .A2(B[2]), .ZN(n152) );
  NAND2_X1 U151 ( .A1(n150), .A2(n24), .ZN(n3) );
  NAND2_X1 U152 ( .A1(n72), .A2(n27), .ZN(n4) );
  NAND2_X1 U153 ( .A1(n70), .A2(n19), .ZN(n2) );
  NAND2_X1 U154 ( .A1(n147), .A2(n40), .ZN(n7) );
  NAND2_X1 U155 ( .A1(n148), .A2(n48), .ZN(n9) );
  NAND2_X1 U156 ( .A1(n151), .A2(n32), .ZN(n5) );
  XOR2_X1 U157 ( .A(n16), .B(n1), .Z(SUM[15]) );
  AND2_X1 U158 ( .A1(n154), .A2(n69), .ZN(SUM[0]) );
  OR2_X1 U159 ( .A1(A[0]), .A2(B[0]), .ZN(n154) );
  NAND2_X1 U160 ( .A1(A[10]), .A2(B[10]), .ZN(n32) );
  NAND2_X1 U161 ( .A1(n82), .A2(n67), .ZN(n14) );
  XOR2_X1 U162 ( .A(n14), .B(n69), .Z(SUM[1]) );
  NAND2_X1 U163 ( .A1(A[0]), .A2(B[0]), .ZN(n69) );
  AOI21_X1 U164 ( .B1(n146), .B2(n152), .A(n62), .ZN(n155) );
  AOI21_X1 U165 ( .B1(n65), .B2(n152), .A(n62), .ZN(n60) );
  INV_X1 U166 ( .A(n66), .ZN(n82) );
  XNOR2_X1 U167 ( .A(n144), .B(n7), .ZN(SUM[8]) );
  OAI21_X1 U168 ( .B1(n138), .B2(n42), .A(n43), .ZN(n41) );
  AOI21_X1 U169 ( .B1(n49), .B2(n148), .A(n46), .ZN(n44) );
  XNOR2_X1 U170 ( .A(n146), .B(n13), .ZN(SUM[2]) );
  AOI21_X1 U171 ( .B1(n144), .B2(n147), .A(n38), .ZN(n36) );
  XOR2_X1 U172 ( .A(n44), .B(n8), .Z(SUM[7]) );
  XNOR2_X1 U173 ( .A(n49), .B(n9), .ZN(SUM[6]) );
  OAI21_X1 U174 ( .B1(n142), .B2(n50), .A(n51), .ZN(n49) );
  AOI21_X1 U175 ( .B1(n141), .B2(n149), .A(n54), .ZN(n52) );
  XNOR2_X1 U176 ( .A(n141), .B(n11), .ZN(SUM[4]) );
  XOR2_X1 U177 ( .A(n52), .B(n10), .Z(SUM[5]) );
  NAND2_X1 U178 ( .A1(n152), .A2(n64), .ZN(n13) );
  NAND2_X1 U179 ( .A1(A[2]), .A2(B[2]), .ZN(n64) );
  NOR2_X1 U180 ( .A1(A[1]), .A2(B[1]), .ZN(n66) );
  OAI21_X1 U181 ( .B1(n66), .B2(n69), .A(n67), .ZN(n65) );
  OAI21_X1 U182 ( .B1(n60), .B2(n58), .A(n59), .ZN(n57) );
  CLKBUF_X1 U183 ( .A(n20), .Z(n156) );
  XNOR2_X1 U184 ( .A(n139), .B(n3), .ZN(SUM[12]) );
  XOR2_X1 U185 ( .A(n28), .B(n4), .Z(SUM[11]) );
  AOI21_X1 U186 ( .B1(n25), .B2(n150), .A(n22), .ZN(n20) );
  OAI21_X1 U187 ( .B1(n143), .B2(n26), .A(n27), .ZN(n25) );
  AOI21_X1 U188 ( .B1(n140), .B2(n151), .A(n30), .ZN(n28) );
  XNOR2_X1 U189 ( .A(n140), .B(n5), .ZN(SUM[10]) );
  XOR2_X1 U190 ( .A(n155), .B(n12), .Z(SUM[3]) );
  OAI21_X1 U191 ( .B1(n145), .B2(n34), .A(n35), .ZN(n33) );
  NAND2_X1 U192 ( .A1(A[1]), .A2(B[1]), .ZN(n67) );
  OAI21_X1 U193 ( .B1(n20), .B2(n18), .A(n19), .ZN(n17) );
  XOR2_X1 U194 ( .A(n36), .B(n6), .Z(SUM[9]) );
  XOR2_X1 U195 ( .A(n156), .B(n2), .Z(SUM[13]) );
endmodule


module part2_mac_DW_mult_tc_1 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n3, n7, n8, n9, n10, n11, n12, n15, n16, n17, n18, n19, n20, n21, n22,
         n24, n25, n26, n30, n31, n35, n36, n38, n39, n40, n41, n42, n43, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n65, n66, n67, n68, n69, n70, n71, n72, n73, n75, n77, n78,
         n80, n81, n84, n85, n86, n87, n90, n91, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n139, n140, n143, n145, n146, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n227, n228, n230, n231, n232, n233,
         n234, n235, n236, n238, n240, n241, n242, n243, n244, n245, n246,
         n247, n255, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392;
  assign n146 = a[0];
  assign n227 = b[0];
  assign n244 = a[7];
  assign n245 = a[5];
  assign n246 = a[3];
  assign n247 = a[1];

  FA_X1 U109 ( .A(n153), .B(n100), .CI(n160), .CO(n96), .S(n97) );
  FA_X1 U112 ( .A(n108), .B(n155), .CI(n105), .CO(n102), .S(n103) );
  FA_X1 U113 ( .A(n110), .B(n161), .CI(n168), .CO(n104), .S(n105) );
  FA_X1 U114 ( .A(n114), .B(n116), .CI(n109), .CO(n106), .S(n107) );
  FA_X1 U115 ( .A(n162), .B(n156), .CI(n111), .CO(n108), .S(n109) );
  FA_X1 U121 ( .A(n126), .B(n123), .CI(n121), .CO(n118), .S(n119) );
  FA_X1 U122 ( .A(n177), .B(n164), .CI(n170), .CO(n120), .S(n121) );
  HA_X1 U123 ( .A(n148), .B(n158), .CO(n122), .S(n123) );
  FA_X1 U124 ( .A(n130), .B(n165), .CI(n127), .CO(n124), .S(n125) );
  FA_X1 U125 ( .A(n178), .B(n159), .CI(n171), .CO(n126), .S(n127) );
  FA_X1 U126 ( .A(n172), .B(n179), .CI(n131), .CO(n128), .S(n129) );
  HA_X1 U127 ( .A(n149), .B(n166), .CO(n130), .S(n131) );
  FA_X1 U128 ( .A(n180), .B(n167), .CI(n173), .CO(n132), .S(n133) );
  HA_X1 U129 ( .A(n174), .B(n181), .CO(n134), .S(n135) );
  BUF_X2 U249 ( .A(n245), .Z(n380) );
  OR2_X1 U250 ( .A1(n99), .A2(n102), .ZN(n362) );
  XOR2_X1 U251 ( .A(n174), .B(n181), .Z(n285) );
  BUF_X2 U252 ( .A(n386), .Z(n366) );
  NOR2_X1 U253 ( .A1(n103), .A2(n106), .ZN(n286) );
  OR2_X1 U254 ( .A1(n247), .A2(a[2]), .ZN(n389) );
  XNOR2_X1 U255 ( .A(n115), .B(n364), .ZN(n287) );
  BUF_X2 U256 ( .A(n245), .Z(n381) );
  OR2_X1 U257 ( .A1(a[2]), .A2(n247), .ZN(n288) );
  NAND2_X1 U258 ( .A1(n288), .A2(n388), .ZN(n383) );
  NAND2_X1 U259 ( .A1(n320), .A2(n321), .ZN(n289) );
  OAI22_X1 U260 ( .A1(n363), .A2(n187), .B1(n186), .B2(n391), .ZN(n154) );
  AOI21_X1 U261 ( .B1(n323), .B2(n383), .A(n202), .ZN(n290) );
  INV_X1 U262 ( .A(n290), .ZN(n168) );
  NOR2_X1 U263 ( .A1(n55), .A2(n327), .ZN(n50) );
  OR2_X2 U264 ( .A1(n367), .A2(n369), .ZN(n233) );
  BUF_X2 U265 ( .A(n341), .Z(n391) );
  NOR2_X1 U266 ( .A1(n133), .A2(n134), .ZN(n67) );
  INV_X1 U267 ( .A(n65), .ZN(n291) );
  CLKBUF_X1 U268 ( .A(n359), .Z(n292) );
  AND2_X1 U269 ( .A1(n102), .A2(n99), .ZN(n359) );
  AOI21_X1 U270 ( .B1(n352), .B2(n66), .A(n291), .ZN(n293) );
  OR2_X2 U271 ( .A1(n129), .A2(n132), .ZN(n352) );
  CLKBUF_X1 U272 ( .A(n247), .Z(n294) );
  CLKBUF_X1 U273 ( .A(n247), .Z(n295) );
  NOR3_X1 U274 ( .A1(n297), .A2(n298), .A3(n299), .ZN(product[15]) );
  AND2_X1 U275 ( .A1(n15), .A2(n94), .ZN(n297) );
  AND2_X1 U276 ( .A1(n15), .A2(n152), .ZN(n298) );
  AND2_X1 U277 ( .A1(n152), .A2(n94), .ZN(n299) );
  INV_X1 U278 ( .A(n310), .ZN(n300) );
  NOR2_X1 U279 ( .A1(n327), .A2(n55), .ZN(n301) );
  XOR2_X1 U280 ( .A(n242), .B(b[4]), .Z(n205) );
  CLKBUF_X1 U281 ( .A(n247), .Z(n302) );
  AOI21_X1 U282 ( .B1(n352), .B2(n66), .A(n360), .ZN(n303) );
  BUF_X1 U283 ( .A(n243), .Z(n304) );
  CLKBUF_X1 U284 ( .A(n368), .Z(n305) );
  OAI21_X2 U285 ( .B1(n69), .B2(n67), .A(n68), .ZN(n66) );
  NAND2_X1 U286 ( .A1(n317), .A2(n255), .ZN(n306) );
  NAND2_X1 U287 ( .A1(n231), .A2(n255), .ZN(n307) );
  XOR2_X1 U288 ( .A(n243), .B(b[6]), .Z(n212) );
  CLKBUF_X1 U289 ( .A(n55), .Z(n353) );
  XOR2_X1 U290 ( .A(n152), .B(n94), .Z(n308) );
  XOR2_X1 U291 ( .A(n15), .B(n308), .Z(product[14]) );
  OR2_X1 U292 ( .A1(n46), .A2(n286), .ZN(n309) );
  INV_X1 U293 ( .A(n318), .ZN(n310) );
  XOR2_X1 U294 ( .A(n101), .B(n154), .Z(n311) );
  XOR2_X1 U295 ( .A(n104), .B(n311), .Z(n99) );
  NAND2_X1 U296 ( .A1(n104), .A2(n101), .ZN(n312) );
  NAND2_X1 U297 ( .A1(n104), .A2(n154), .ZN(n313) );
  NAND2_X1 U298 ( .A1(n101), .A2(n154), .ZN(n314) );
  NAND3_X1 U299 ( .A1(n312), .A2(n313), .A3(n314), .ZN(n98) );
  NAND2_X1 U300 ( .A1(n317), .A2(n255), .ZN(n315) );
  NAND2_X1 U301 ( .A1(n231), .A2(n255), .ZN(n316) );
  NAND2_X1 U302 ( .A1(n379), .A2(n378), .ZN(n317) );
  NAND2_X1 U303 ( .A1(n317), .A2(n255), .ZN(n235) );
  NAND2_X1 U304 ( .A1(n246), .A2(n319), .ZN(n320) );
  NAND2_X1 U305 ( .A1(n318), .A2(a[2]), .ZN(n321) );
  NAND2_X1 U306 ( .A1(n320), .A2(n321), .ZN(n230) );
  INV_X1 U307 ( .A(n246), .ZN(n318) );
  INV_X1 U308 ( .A(a[2]), .ZN(n319) );
  CLKBUF_X1 U309 ( .A(n47), .Z(n322) );
  NAND2_X1 U310 ( .A1(n238), .A2(n230), .ZN(n323) );
  NOR2_X1 U311 ( .A1(n106), .A2(n103), .ZN(n324) );
  OAI21_X1 U312 ( .B1(n56), .B2(n52), .A(n53), .ZN(n325) );
  NOR2_X1 U313 ( .A1(n25), .A2(n20), .ZN(n326) );
  NOR2_X1 U314 ( .A1(n287), .A2(n118), .ZN(n327) );
  XOR2_X1 U315 ( .A(n10), .B(n69), .Z(product[4]) );
  XOR2_X1 U316 ( .A(n11), .B(n73), .Z(product[3]) );
  AOI21_X1 U317 ( .B1(n292), .B2(n344), .A(n357), .ZN(n328) );
  OR2_X2 U318 ( .A1(n98), .A2(n97), .ZN(n344) );
  OAI21_X1 U319 ( .B1(n61), .B2(n59), .A(n60), .ZN(n329) );
  NOR2_X1 U320 ( .A1(n112), .A2(n107), .ZN(n46) );
  INV_X1 U321 ( .A(n20), .ZN(n81) );
  INV_X1 U322 ( .A(n357), .ZN(n30) );
  INV_X1 U323 ( .A(n292), .ZN(n35) );
  OAI21_X1 U324 ( .B1(n303), .B2(n59), .A(n60), .ZN(n58) );
  NOR2_X1 U325 ( .A1(n113), .A2(n118), .ZN(n52) );
  INV_X1 U326 ( .A(n94), .ZN(n95) );
  NOR2_X1 U327 ( .A1(n96), .A2(n95), .ZN(n20) );
  NAND2_X1 U328 ( .A1(n96), .A2(n95), .ZN(n21) );
  NAND2_X1 U329 ( .A1(n90), .A2(n68), .ZN(n10) );
  INV_X1 U330 ( .A(n136), .ZN(n152) );
  NAND2_X1 U331 ( .A1(n330), .A2(n331), .ZN(n158) );
  OR2_X1 U332 ( .A1(n232), .A2(n191), .ZN(n330) );
  OR2_X1 U333 ( .A1(n190), .A2(n342), .ZN(n331) );
  OR2_X1 U334 ( .A1(n183), .A2(n151), .ZN(n332) );
  OR2_X1 U335 ( .A1(n182), .A2(n175), .ZN(n333) );
  OR2_X1 U336 ( .A1(n227), .A2(n240), .ZN(n192) );
  OR2_X1 U337 ( .A1(n227), .A2(n300), .ZN(n210) );
  OR2_X1 U338 ( .A1(n227), .A2(n304), .ZN(n219) );
  XOR2_X1 U339 ( .A(n48), .B(n334), .Z(product[9]) );
  AND2_X1 U340 ( .A1(n85), .A2(n322), .ZN(n334) );
  XOR2_X1 U341 ( .A(n57), .B(n7), .Z(product[7]) );
  AND2_X1 U342 ( .A1(n227), .A2(n137), .ZN(n159) );
  AND2_X1 U343 ( .A1(n227), .A2(n143), .ZN(n175) );
  AND2_X1 U344 ( .A1(n332), .A2(n80), .ZN(product[1]) );
  XOR2_X1 U345 ( .A(n242), .B(b[5]), .Z(n204) );
  XNOR2_X1 U346 ( .A(n22), .B(n336), .ZN(product[13]) );
  AND2_X1 U347 ( .A1(n81), .A2(n21), .ZN(n336) );
  XNOR2_X1 U348 ( .A(n31), .B(n337), .ZN(product[12]) );
  AND2_X1 U349 ( .A1(n344), .A2(n30), .ZN(n337) );
  NAND2_X1 U350 ( .A1(n347), .A2(n35), .ZN(n3) );
  XOR2_X1 U351 ( .A(n54), .B(n338), .Z(product[8]) );
  AND2_X1 U352 ( .A1(n86), .A2(n53), .ZN(n338) );
  AND2_X1 U353 ( .A1(n227), .A2(n146), .ZN(product[0]) );
  XNOR2_X1 U354 ( .A(n12), .B(n78), .ZN(product[2]) );
  XNOR2_X1 U355 ( .A(n43), .B(n339), .ZN(product[10]) );
  AND2_X1 U356 ( .A1(n84), .A2(n42), .ZN(n339) );
  NAND2_X1 U357 ( .A1(n103), .A2(n106), .ZN(n42) );
  XOR2_X1 U358 ( .A(n244), .B(a[6]), .Z(n340) );
  XNOR2_X1 U359 ( .A(n380), .B(a[6]), .ZN(n341) );
  XNOR2_X1 U360 ( .A(n380), .B(a[6]), .ZN(n342) );
  XNOR2_X1 U361 ( .A(n381), .B(a[6]), .ZN(n236) );
  AOI21_X1 U362 ( .B1(n301), .B2(n329), .A(n51), .ZN(n343) );
  NAND2_X1 U363 ( .A1(n348), .A2(n230), .ZN(n345) );
  CLKBUF_X1 U364 ( .A(n352), .Z(n346) );
  INV_X1 U365 ( .A(n100), .ZN(n101) );
  AND2_X1 U366 ( .A1(n227), .A2(n140), .ZN(n167) );
  CLKBUF_X1 U367 ( .A(n362), .Z(n347) );
  NAND2_X1 U368 ( .A1(n388), .A2(n389), .ZN(n348) );
  INV_X1 U369 ( .A(n242), .ZN(n349) );
  OAI22_X1 U370 ( .A1(n316), .A2(n215), .B1(n214), .B2(n255), .ZN(n180) );
  OAI22_X1 U371 ( .A1(n316), .A2(n214), .B1(n213), .B2(n255), .ZN(n179) );
  CLKBUF_X1 U372 ( .A(n125), .Z(n350) );
  AND2_X1 U373 ( .A1(n362), .A2(n344), .ZN(n351) );
  INV_X1 U374 ( .A(n327), .ZN(n86) );
  INV_X1 U375 ( .A(n67), .ZN(n90) );
  INV_X1 U376 ( .A(n360), .ZN(n65) );
  AND2_X1 U377 ( .A1(n148), .A2(n158), .ZN(n354) );
  NOR2_X1 U378 ( .A1(n119), .A2(n124), .ZN(n55) );
  INV_X1 U379 ( .A(n353), .ZN(n87) );
  OR2_X1 U380 ( .A1(n350), .A2(n128), .ZN(n355) );
  NAND2_X1 U381 ( .A1(n355), .A2(n60), .ZN(n8) );
  CLKBUF_X1 U382 ( .A(n56), .Z(n356) );
  AND2_X1 U383 ( .A1(n98), .A2(n97), .ZN(n357) );
  NAND2_X1 U384 ( .A1(n346), .A2(n65), .ZN(n9) );
  OR2_X1 U385 ( .A1(n227), .A2(n241), .ZN(n201) );
  INV_X1 U386 ( .A(n46), .ZN(n85) );
  CLKBUF_X1 U387 ( .A(n246), .Z(n358) );
  INV_X1 U388 ( .A(n77), .ZN(n75) );
  NAND2_X1 U389 ( .A1(n333), .A2(n77), .ZN(n12) );
  INV_X1 U390 ( .A(n71), .ZN(n91) );
  OAI22_X1 U391 ( .A1(n307), .A2(n213), .B1(n212), .B2(n255), .ZN(n178) );
  INV_X1 U392 ( .A(n322), .ZN(n45) );
  OAI22_X1 U393 ( .A1(n235), .A2(n212), .B1(n211), .B2(n255), .ZN(n177) );
  AND2_X1 U394 ( .A1(n129), .A2(n132), .ZN(n360) );
  XNOR2_X1 U395 ( .A(n361), .B(n354), .ZN(n115) );
  XNOR2_X1 U396 ( .A(n176), .B(n163), .ZN(n361) );
  NAND2_X1 U397 ( .A1(n340), .A2(n341), .ZN(n363) );
  XNOR2_X1 U398 ( .A(n115), .B(n364), .ZN(n113) );
  XNOR2_X1 U399 ( .A(n120), .B(n117), .ZN(n364) );
  AOI21_X1 U400 ( .B1(n333), .B2(n78), .A(n75), .ZN(n73) );
  INV_X1 U401 ( .A(n324), .ZN(n84) );
  NOR2_X1 U402 ( .A1(n46), .A2(n324), .ZN(n39) );
  NOR2_X1 U403 ( .A1(n103), .A2(n106), .ZN(n41) );
  BUF_X1 U404 ( .A(n386), .Z(n365) );
  NAND2_X1 U405 ( .A1(n133), .A2(n134), .ZN(n68) );
  NAND2_X1 U406 ( .A1(n87), .A2(n356), .ZN(n7) );
  OAI21_X1 U407 ( .B1(n57), .B2(n353), .A(n356), .ZN(n54) );
  NOR2_X1 U408 ( .A1(n285), .A2(n150), .ZN(n71) );
  XNOR2_X1 U409 ( .A(n380), .B(a[4]), .ZN(n367) );
  INV_X1 U410 ( .A(n328), .ZN(n24) );
  NAND2_X1 U411 ( .A1(n125), .A2(n128), .ZN(n60) );
  NOR2_X1 U412 ( .A1(n125), .A2(n128), .ZN(n59) );
  NAND2_X1 U413 ( .A1(n287), .A2(n118), .ZN(n53) );
  NAND2_X1 U414 ( .A1(n119), .A2(n124), .ZN(n56) );
  OR2_X2 U415 ( .A1(n367), .A2(n369), .ZN(n368) );
  XNOR2_X1 U416 ( .A(n244), .B(b[7]), .ZN(n184) );
  XNOR2_X1 U417 ( .A(n244), .B(b[6]), .ZN(n185) );
  XNOR2_X1 U418 ( .A(n244), .B(b[5]), .ZN(n186) );
  XNOR2_X1 U419 ( .A(n244), .B(b[4]), .ZN(n187) );
  INV_X1 U420 ( .A(n80), .ZN(n78) );
  OAI22_X1 U421 ( .A1(n315), .A2(n304), .B1(n219), .B2(n255), .ZN(n151) );
  OR2_X1 U422 ( .A1(n169), .A2(n157), .ZN(n116) );
  XNOR2_X1 U423 ( .A(n169), .B(n157), .ZN(n117) );
  NAND2_X1 U424 ( .A1(n362), .A2(n344), .ZN(n25) );
  XOR2_X1 U425 ( .A(n246), .B(a[4]), .Z(n369) );
  NAND2_X1 U426 ( .A1(n176), .A2(n163), .ZN(n370) );
  NAND2_X1 U427 ( .A1(n122), .A2(n176), .ZN(n371) );
  NAND2_X1 U428 ( .A1(n163), .A2(n354), .ZN(n372) );
  NAND3_X1 U429 ( .A1(n372), .A2(n371), .A3(n370), .ZN(n114) );
  NAND2_X1 U430 ( .A1(n120), .A2(n117), .ZN(n373) );
  NAND2_X1 U431 ( .A1(n120), .A2(n115), .ZN(n374) );
  NAND2_X1 U432 ( .A1(n117), .A2(n115), .ZN(n375) );
  NAND3_X1 U433 ( .A1(n373), .A2(n374), .A3(n375), .ZN(n112) );
  NAND2_X1 U434 ( .A1(n247), .A2(n377), .ZN(n378) );
  NAND2_X1 U435 ( .A1(n376), .A2(n146), .ZN(n379) );
  NAND2_X1 U436 ( .A1(n379), .A2(n378), .ZN(n231) );
  INV_X1 U437 ( .A(n247), .ZN(n376) );
  INV_X1 U438 ( .A(n146), .ZN(n377) );
  INV_X1 U439 ( .A(n329), .ZN(n57) );
  XOR2_X1 U440 ( .A(n8), .B(n293), .Z(product[6]) );
  INV_X1 U441 ( .A(n244), .ZN(n240) );
  XNOR2_X1 U442 ( .A(n244), .B(b[3]), .ZN(n188) );
  XNOR2_X1 U443 ( .A(n244), .B(b[2]), .ZN(n189) );
  NAND2_X1 U444 ( .A1(n289), .A2(n348), .ZN(n382) );
  NAND2_X1 U445 ( .A1(n388), .A2(n389), .ZN(n384) );
  OAI22_X1 U446 ( .A1(n234), .A2(n203), .B1(n383), .B2(n202), .ZN(n385) );
  NAND2_X1 U447 ( .A1(n238), .A2(n289), .ZN(n234) );
  NAND2_X1 U448 ( .A1(n388), .A2(n389), .ZN(n238) );
  AOI21_X1 U449 ( .B1(n352), .B2(n66), .A(n360), .ZN(n61) );
  OAI22_X1 U450 ( .A1(n316), .A2(n218), .B1(n217), .B2(n255), .ZN(n183) );
  INV_X1 U451 ( .A(n385), .ZN(n111) );
  INV_X1 U452 ( .A(n145), .ZN(n176) );
  XNOR2_X1 U453 ( .A(n246), .B(a[4]), .ZN(n386) );
  XNOR2_X1 U454 ( .A(n9), .B(n66), .ZN(product[5]) );
  NAND2_X1 U455 ( .A1(n182), .A2(n175), .ZN(n77) );
  OAI22_X1 U456 ( .A1(n315), .A2(n217), .B1(n216), .B2(n255), .ZN(n182) );
  OAI22_X1 U457 ( .A1(n211), .A2(n315), .B1(n211), .B2(n255), .ZN(n145) );
  OAI22_X1 U458 ( .A1(n306), .A2(n216), .B1(n215), .B2(n255), .ZN(n181) );
  INV_X1 U459 ( .A(n139), .ZN(n160) );
  CLKBUF_X1 U460 ( .A(n247), .Z(n387) );
  NAND2_X1 U461 ( .A1(n247), .A2(a[2]), .ZN(n388) );
  NAND2_X1 U462 ( .A1(n228), .A2(n342), .ZN(n390) );
  XOR2_X1 U463 ( .A(n244), .B(a[6]), .Z(n228) );
  NAND2_X1 U464 ( .A1(n228), .A2(n236), .ZN(n232) );
  NAND2_X1 U465 ( .A1(n183), .A2(n151), .ZN(n80) );
  OAI21_X1 U466 ( .B1(n49), .B2(n309), .A(n38), .ZN(n392) );
  OAI21_X1 U467 ( .B1(n343), .B2(n309), .A(n38), .ZN(n36) );
  XNOR2_X1 U468 ( .A(n244), .B(n227), .ZN(n191) );
  XNOR2_X1 U469 ( .A(n244), .B(b[1]), .ZN(n190) );
  INV_X1 U470 ( .A(n70), .ZN(n69) );
  OAI21_X1 U471 ( .B1(n26), .B2(n20), .A(n21), .ZN(n19) );
  NOR2_X1 U472 ( .A1(n25), .A2(n20), .ZN(n18) );
  AOI21_X1 U473 ( .B1(n359), .B2(n344), .A(n357), .ZN(n26) );
  NAND2_X1 U474 ( .A1(n91), .A2(n72), .ZN(n11) );
  OAI21_X1 U475 ( .B1(n73), .B2(n71), .A(n72), .ZN(n70) );
  OAI22_X1 U476 ( .A1(n305), .A2(n199), .B1(n198), .B2(n365), .ZN(n165) );
  OAI22_X1 U477 ( .A1(n368), .A2(n197), .B1(n196), .B2(n365), .ZN(n163) );
  OAI22_X1 U478 ( .A1(n233), .A2(n198), .B1(n197), .B2(n366), .ZN(n164) );
  OAI22_X1 U479 ( .A1(n368), .A2(n194), .B1(n193), .B2(n365), .ZN(n100) );
  OAI22_X1 U480 ( .A1(n196), .A2(n368), .B1(n195), .B2(n365), .ZN(n162) );
  INV_X1 U481 ( .A(n366), .ZN(n140) );
  OAI22_X1 U482 ( .A1(n193), .A2(n305), .B1(n193), .B2(n366), .ZN(n139) );
  OAI22_X1 U483 ( .A1(n368), .A2(n195), .B1(n194), .B2(n366), .ZN(n161) );
  XNOR2_X1 U484 ( .A(n349), .B(b[3]), .ZN(n206) );
  OAI22_X1 U485 ( .A1(n233), .A2(n241), .B1(n201), .B2(n365), .ZN(n149) );
  OAI22_X1 U486 ( .A1(n233), .A2(n200), .B1(n199), .B2(n366), .ZN(n166) );
  XNOR2_X1 U487 ( .A(n310), .B(b[2]), .ZN(n207) );
  INV_X1 U488 ( .A(n246), .ZN(n242) );
  XNOR2_X1 U489 ( .A(n358), .B(b[6]), .ZN(n203) );
  XNOR2_X1 U490 ( .A(n310), .B(n227), .ZN(n209) );
  XNOR2_X1 U491 ( .A(n358), .B(b[7]), .ZN(n202) );
  XNOR2_X1 U492 ( .A(n310), .B(b[1]), .ZN(n208) );
  OAI22_X1 U493 ( .A1(n184), .A2(n390), .B1(n184), .B2(n391), .ZN(n136) );
  OAI22_X1 U494 ( .A1(n363), .A2(n185), .B1(n184), .B2(n391), .ZN(n94) );
  OAI22_X1 U495 ( .A1(n390), .A2(n188), .B1(n187), .B2(n391), .ZN(n155) );
  OAI22_X1 U496 ( .A1(n363), .A2(n190), .B1(n189), .B2(n391), .ZN(n157) );
  OAI22_X1 U497 ( .A1(n390), .A2(n186), .B1(n185), .B2(n391), .ZN(n153) );
  OAI22_X1 U498 ( .A1(n363), .A2(n189), .B1(n188), .B2(n342), .ZN(n156) );
  INV_X1 U499 ( .A(n342), .ZN(n137) );
  OAI22_X1 U500 ( .A1(n390), .A2(n240), .B1(n192), .B2(n342), .ZN(n148) );
  XNOR2_X1 U501 ( .A(n381), .B(b[2]), .ZN(n198) );
  XNOR2_X1 U502 ( .A(n381), .B(b[3]), .ZN(n197) );
  XNOR2_X1 U503 ( .A(n381), .B(b[4]), .ZN(n196) );
  XNOR2_X1 U504 ( .A(n381), .B(b[5]), .ZN(n195) );
  XNOR2_X1 U505 ( .A(n381), .B(b[7]), .ZN(n193) );
  XNOR2_X1 U506 ( .A(n381), .B(n227), .ZN(n200) );
  XNOR2_X1 U507 ( .A(n381), .B(b[6]), .ZN(n194) );
  XNOR2_X1 U508 ( .A(n381), .B(b[1]), .ZN(n199) );
  INV_X1 U509 ( .A(n381), .ZN(n241) );
  AOI21_X1 U510 ( .B1(n48), .B2(n85), .A(n45), .ZN(n43) );
  NAND2_X1 U511 ( .A1(n135), .A2(n150), .ZN(n72) );
  INV_X1 U512 ( .A(n40), .ZN(n38) );
  AOI21_X1 U513 ( .B1(n40), .B2(n18), .A(n19), .ZN(n17) );
  OAI21_X1 U514 ( .B1(n47), .B2(n41), .A(n42), .ZN(n40) );
  NAND2_X1 U515 ( .A1(n107), .A2(n112), .ZN(n47) );
  AOI21_X1 U516 ( .B1(n50), .B2(n58), .A(n325), .ZN(n49) );
  OAI21_X1 U517 ( .B1(n52), .B2(n56), .A(n53), .ZN(n51) );
  NAND2_X1 U518 ( .A1(n39), .A2(n326), .ZN(n16) );
  XNOR2_X1 U519 ( .A(n392), .B(n3), .ZN(product[11]) );
  AOI21_X1 U520 ( .B1(n392), .B2(n347), .A(n292), .ZN(n31) );
  AOI21_X1 U521 ( .B1(n36), .B2(n351), .A(n24), .ZN(n22) );
  OAI21_X1 U522 ( .B1(n49), .B2(n16), .A(n17), .ZN(n15) );
  INV_X1 U523 ( .A(n343), .ZN(n48) );
  OAI22_X1 U524 ( .A1(n382), .A2(n204), .B1(n203), .B2(n383), .ZN(n169) );
  OAI22_X1 U525 ( .A1(n382), .A2(n207), .B1(n206), .B2(n384), .ZN(n172) );
  OAI22_X1 U526 ( .A1(n345), .A2(n206), .B1(n383), .B2(n205), .ZN(n171) );
  OAI22_X1 U527 ( .A1(n345), .A2(n205), .B1(n204), .B2(n384), .ZN(n170) );
  OAI22_X1 U528 ( .A1(n382), .A2(n208), .B1(n207), .B2(n384), .ZN(n173) );
  OAI22_X1 U529 ( .A1(n382), .A2(n300), .B1(n210), .B2(n383), .ZN(n150) );
  OAI22_X1 U530 ( .A1(n234), .A2(n203), .B1(n202), .B2(n383), .ZN(n110) );
  XNOR2_X1 U531 ( .A(n387), .B(b[5]), .ZN(n213) );
  XNOR2_X1 U532 ( .A(n387), .B(b[4]), .ZN(n214) );
  XNOR2_X1 U533 ( .A(n294), .B(b[7]), .ZN(n211) );
  INV_X1 U534 ( .A(n384), .ZN(n143) );
  OAI22_X1 U535 ( .A1(n323), .A2(n209), .B1(n208), .B2(n384), .ZN(n174) );
  XNOR2_X1 U536 ( .A(n295), .B(b[3]), .ZN(n215) );
  XNOR2_X1 U537 ( .A(n302), .B(b[2]), .ZN(n216) );
  XNOR2_X1 U538 ( .A(n302), .B(n227), .ZN(n218) );
  XNOR2_X1 U539 ( .A(n302), .B(b[1]), .ZN(n217) );
  INV_X1 U540 ( .A(n247), .ZN(n243) );
  INV_X2 U541 ( .A(n146), .ZN(n255) );
endmodule


module part2_mac ( clk, reset, a, b, valid_in, f, valid_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] f;
  input clk, reset, valid_in;
  output valid_out;
  wire   N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41,
         N42, N43, n109, n110, n111, n112, n113, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227;
  wire   [7:0] a_reg;
  wire   [7:0] b_reg;
  wire   [15:0] mul_w;
  wire   [15:0] multa;

  DFF_X1 \a_reg_reg[4]  ( .D(n207), .CK(clk), .Q(a_reg[4]), .QN(n118) );
  DFF_X1 \multa_reg[14]  ( .D(n213), .CK(clk), .Q(multa[14]) );
  DFF_X1 \multa_reg[13]  ( .D(n214), .CK(clk), .Q(multa[13]) );
  DFF_X1 \multa_reg[12]  ( .D(n215), .CK(clk), .Q(multa[12]) );
  DFF_X1 \multa_reg[9]  ( .D(n218), .CK(clk), .Q(multa[9]) );
  DFF_X1 \f_reg_reg[0]  ( .D(n196), .CK(clk), .Q(f[0]) );
  part2_mac_DW01_add_1 add_69 ( .A(f), .B(multa), .CI(1'b0), .SUM({N43, N42, 
        N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28})
         );
  part2_mac_DW_mult_tc_1 mult_57 ( .a({n121, a_reg[6:2], n123, a_reg[0]}), .b(
        b_reg), .product(mul_w) );
  DFF_X1 \a_reg_reg[3]  ( .D(n208), .CK(clk), .Q(a_reg[3]), .QN(n124) );
  DFF_X1 \a_reg_reg[1]  ( .D(n210), .CK(clk), .QN(n122) );
  DFF_X1 \a_reg_reg[7]  ( .D(n205), .CK(clk), .Q(a_reg[7]), .QN(n120) );
  DFF_X1 \multa_reg[10]  ( .D(n217), .CK(clk), .Q(multa[10]) );
  DFF_X1 valid_out_reg ( .D(n112), .CK(clk), .Q(valid_out) );
  DFF_X1 enable_f_reg ( .D(n110), .CK(clk), .QN(n111) );
  DFF_X1 \f_reg_reg[2]  ( .D(n194), .CK(clk), .Q(f[2]) );
  DFF_X1 \multa_reg[0]  ( .D(n227), .CK(clk), .Q(multa[0]) );
  DFF_X1 \f_reg_reg[1]  ( .D(n195), .CK(clk), .Q(f[1]) );
  DFF_X1 enable_multa_reg ( .D(n180), .CK(clk), .QN(n109) );
  DFF_X1 \f_reg_reg[3]  ( .D(n193), .CK(clk), .Q(f[3]) );
  DFF_X1 \f_reg_reg[4]  ( .D(n192), .CK(clk), .Q(f[4]) );
  DFF_X1 \b_reg_reg[7]  ( .D(n197), .CK(clk), .Q(b_reg[7]) );
  DFF_X1 \b_reg_reg[6]  ( .D(n198), .CK(clk), .Q(b_reg[6]) );
  DFF_X1 \b_reg_reg[5]  ( .D(n199), .CK(clk), .Q(b_reg[5]) );
  DFF_X1 \b_reg_reg[4]  ( .D(n200), .CK(clk), .Q(b_reg[4]) );
  DFF_X1 \b_reg_reg[3]  ( .D(n201), .CK(clk), .Q(b_reg[3]) );
  DFF_X1 \b_reg_reg[2]  ( .D(n202), .CK(clk), .Q(b_reg[2]) );
  DFF_X1 \b_reg_reg[1]  ( .D(n203), .CK(clk), .Q(b_reg[1]) );
  DFF_X1 \a_reg_reg[6]  ( .D(n206), .CK(clk), .Q(a_reg[6]) );
  DFF_X1 \a_reg_reg[2]  ( .D(n209), .CK(clk), .Q(a_reg[2]) );
  DFF_X1 \a_reg_reg[0]  ( .D(n211), .CK(clk), .Q(a_reg[0]) );
  DFF_X1 \b_reg_reg[0]  ( .D(n204), .CK(clk), .Q(b_reg[0]) );
  DFF_X1 \f_reg_reg[6]  ( .D(n190), .CK(clk), .Q(f[6]) );
  DFF_X1 \multa_reg[1]  ( .D(n226), .CK(clk), .Q(multa[1]) );
  DFF_X1 \f_reg_reg[5]  ( .D(n191), .CK(clk), .Q(f[5]) );
  DFF_X1 \multa_reg[2]  ( .D(n225), .CK(clk), .Q(multa[2]) );
  DFF_X1 \f_reg_reg[7]  ( .D(n189), .CK(clk), .Q(f[7]) );
  DFF_X1 \f_reg_reg[8]  ( .D(n188), .CK(clk), .Q(f[8]) );
  DFF_X1 \multa_reg[3]  ( .D(n224), .CK(clk), .Q(multa[3]) );
  DFF_X1 \f_reg_reg[9]  ( .D(n187), .CK(clk), .Q(f[9]) );
  DFF_X1 \f_reg_reg[10]  ( .D(n186), .CK(clk), .Q(f[10]) );
  DFF_X1 \multa_reg[4]  ( .D(n223), .CK(clk), .Q(multa[4]) );
  DFF_X1 \f_reg_reg[11]  ( .D(n185), .CK(clk), .Q(f[11]) );
  DFF_X1 \f_reg_reg[12]  ( .D(n184), .CK(clk), .Q(f[12]) );
  DFF_X1 \multa_reg[5]  ( .D(n222), .CK(clk), .Q(multa[5]) );
  DFF_X1 \f_reg_reg[13]  ( .D(n183), .CK(clk), .Q(f[13]) );
  DFF_X1 \multa_reg[6]  ( .D(n221), .CK(clk), .Q(multa[6]) );
  DFF_X1 \multa_reg[7]  ( .D(n220), .CK(clk), .Q(multa[7]) );
  DFF_X1 \multa_reg[8]  ( .D(n219), .CK(clk), .Q(multa[8]) );
  DFF_X1 \f_reg_reg[14]  ( .D(n182), .CK(clk), .Q(f[14]) );
  DFF_X1 \multa_reg[11]  ( .D(n216), .CK(clk), .Q(multa[11]) );
  DFF_X1 \f_reg_reg[15]  ( .D(n181), .CK(clk), .Q(f[15]) );
  SDFF_X1 \a_reg_reg[5]  ( .D(1'b1), .SI(1'b0), .SE(n145), .CK(clk), .Q(
        a_reg[5]) );
  DFF_X2 \multa_reg[15]  ( .D(n212), .CK(clk), .Q(multa[15]) );
  INV_X1 U109 ( .A(n160), .ZN(n176) );
  NOR2_X1 U112 ( .A1(reset), .A2(n109), .ZN(n110) );
  NOR2_X1 U113 ( .A1(reset), .A2(n111), .ZN(n112) );
  AOI22_X1 U114 ( .A1(mul_w[15]), .A2(n116), .B1(n176), .B2(multa[15]), .ZN(
        n161) );
  AOI22_X1 U115 ( .A1(mul_w[10]), .A2(n116), .B1(n176), .B2(multa[10]), .ZN(
        n166) );
  AOI22_X1 U116 ( .A1(mul_w[9]), .A2(n116), .B1(n176), .B2(multa[9]), .ZN(n167) );
  AOI22_X1 U117 ( .A1(mul_w[13]), .A2(n116), .B1(n176), .B2(multa[13]), .ZN(
        n163) );
  AOI22_X1 U118 ( .A1(mul_w[12]), .A2(n116), .B1(n176), .B2(multa[12]), .ZN(
        n164) );
  CLKBUF_X1 U119 ( .A(n123), .Z(n113) );
  INV_X1 U120 ( .A(n142), .ZN(n180) );
  INV_X1 U121 ( .A(n126), .ZN(n178) );
  AND2_X1 U122 ( .A1(n126), .A2(n159), .ZN(n115) );
  AND2_X1 U123 ( .A1(n160), .A2(n159), .ZN(n116) );
  AND2_X1 U124 ( .A1(n142), .A2(n159), .ZN(n117) );
  INV_X1 U125 ( .A(n118), .ZN(n119) );
  INV_X2 U126 ( .A(n120), .ZN(n121) );
  INV_X1 U127 ( .A(n124), .ZN(n125) );
  INV_X2 U128 ( .A(n122), .ZN(n123) );
  INV_X1 U129 ( .A(reset), .ZN(n159) );
  NAND2_X1 U130 ( .A1(valid_in), .A2(n159), .ZN(n142) );
  NAND2_X1 U131 ( .A1(n159), .A2(n111), .ZN(n126) );
  AOI22_X1 U132 ( .A1(f[15]), .A2(n178), .B1(N43), .B2(n115), .ZN(n127) );
  INV_X1 U133 ( .A(n127), .ZN(n181) );
  AOI22_X1 U134 ( .A1(f[14]), .A2(n178), .B1(N42), .B2(n115), .ZN(n128) );
  INV_X1 U135 ( .A(n128), .ZN(n182) );
  AOI22_X1 U136 ( .A1(f[13]), .A2(n178), .B1(N41), .B2(n115), .ZN(n129) );
  INV_X1 U137 ( .A(n129), .ZN(n183) );
  AOI22_X1 U138 ( .A1(f[12]), .A2(n178), .B1(N40), .B2(n115), .ZN(n130) );
  INV_X1 U139 ( .A(n130), .ZN(n184) );
  AOI22_X1 U140 ( .A1(f[11]), .A2(n178), .B1(N39), .B2(n115), .ZN(n131) );
  INV_X1 U141 ( .A(n131), .ZN(n185) );
  AOI22_X1 U142 ( .A1(f[10]), .A2(n178), .B1(N38), .B2(n115), .ZN(n132) );
  INV_X1 U143 ( .A(n132), .ZN(n186) );
  AOI22_X1 U144 ( .A1(f[9]), .A2(n178), .B1(N37), .B2(n115), .ZN(n133) );
  INV_X1 U145 ( .A(n133), .ZN(n187) );
  AOI22_X1 U146 ( .A1(f[8]), .A2(n178), .B1(N36), .B2(n115), .ZN(n134) );
  INV_X1 U147 ( .A(n134), .ZN(n188) );
  AOI22_X1 U148 ( .A1(f[7]), .A2(n178), .B1(N35), .B2(n115), .ZN(n135) );
  INV_X1 U149 ( .A(n135), .ZN(n189) );
  AOI22_X1 U150 ( .A1(f[6]), .A2(n178), .B1(N34), .B2(n115), .ZN(n136) );
  INV_X1 U151 ( .A(n136), .ZN(n190) );
  AOI22_X1 U152 ( .A1(f[5]), .A2(n178), .B1(N33), .B2(n115), .ZN(n137) );
  INV_X1 U153 ( .A(n137), .ZN(n191) );
  AOI22_X1 U154 ( .A1(f[4]), .A2(n178), .B1(N32), .B2(n115), .ZN(n138) );
  INV_X1 U155 ( .A(n138), .ZN(n192) );
  AOI22_X1 U156 ( .A1(f[3]), .A2(n178), .B1(N31), .B2(n115), .ZN(n139) );
  INV_X1 U157 ( .A(n139), .ZN(n193) );
  AOI22_X1 U158 ( .A1(f[2]), .A2(n178), .B1(N30), .B2(n115), .ZN(n140) );
  INV_X1 U159 ( .A(n140), .ZN(n194) );
  AOI22_X1 U160 ( .A1(f[1]), .A2(n178), .B1(N29), .B2(n115), .ZN(n141) );
  INV_X1 U161 ( .A(n141), .ZN(n195) );
  AOI22_X1 U162 ( .A1(a[7]), .A2(n180), .B1(a_reg[7]), .B2(n117), .ZN(n143) );
  INV_X1 U163 ( .A(n143), .ZN(n205) );
  AOI22_X1 U164 ( .A1(a[6]), .A2(n180), .B1(a_reg[6]), .B2(n117), .ZN(n144) );
  INV_X1 U165 ( .A(n144), .ZN(n206) );
  AOI22_X1 U166 ( .A1(a[5]), .A2(n180), .B1(a_reg[5]), .B2(n117), .ZN(n145) );
  AOI22_X1 U167 ( .A1(a[4]), .A2(n180), .B1(n119), .B2(n117), .ZN(n146) );
  INV_X1 U168 ( .A(n146), .ZN(n207) );
  AOI22_X1 U169 ( .A1(a[3]), .A2(n180), .B1(n125), .B2(n117), .ZN(n147) );
  INV_X1 U170 ( .A(n147), .ZN(n208) );
  AOI22_X1 U171 ( .A1(a[2]), .A2(n180), .B1(a_reg[2]), .B2(n117), .ZN(n148) );
  INV_X1 U172 ( .A(n148), .ZN(n209) );
  AOI22_X1 U173 ( .A1(a[1]), .A2(n180), .B1(n113), .B2(n117), .ZN(n149) );
  INV_X1 U174 ( .A(n149), .ZN(n210) );
  AOI22_X1 U175 ( .A1(a[0]), .A2(n180), .B1(a_reg[0]), .B2(n117), .ZN(n150) );
  INV_X1 U176 ( .A(n150), .ZN(n211) );
  AOI22_X1 U177 ( .A1(b[7]), .A2(n180), .B1(b_reg[7]), .B2(n117), .ZN(n151) );
  INV_X1 U178 ( .A(n151), .ZN(n197) );
  AOI22_X1 U179 ( .A1(b[6]), .A2(n180), .B1(b_reg[6]), .B2(n117), .ZN(n152) );
  INV_X1 U180 ( .A(n152), .ZN(n198) );
  AOI22_X1 U181 ( .A1(b[5]), .A2(n180), .B1(b_reg[5]), .B2(n117), .ZN(n153) );
  INV_X1 U182 ( .A(n153), .ZN(n199) );
  AOI22_X1 U183 ( .A1(b[4]), .A2(n180), .B1(b_reg[4]), .B2(n117), .ZN(n154) );
  INV_X1 U184 ( .A(n154), .ZN(n200) );
  AOI22_X1 U185 ( .A1(b[3]), .A2(n180), .B1(b_reg[3]), .B2(n117), .ZN(n155) );
  INV_X1 U186 ( .A(n155), .ZN(n201) );
  AOI22_X1 U187 ( .A1(b[2]), .A2(n180), .B1(b_reg[2]), .B2(n117), .ZN(n156) );
  INV_X1 U188 ( .A(n156), .ZN(n202) );
  AOI22_X1 U189 ( .A1(b[1]), .A2(n180), .B1(b_reg[1]), .B2(n117), .ZN(n157) );
  INV_X1 U190 ( .A(n157), .ZN(n203) );
  AOI22_X1 U191 ( .A1(b[0]), .A2(n180), .B1(b_reg[0]), .B2(n117), .ZN(n158) );
  INV_X1 U192 ( .A(n158), .ZN(n204) );
  NAND2_X1 U193 ( .A1(n159), .A2(n109), .ZN(n160) );
  INV_X1 U194 ( .A(n161), .ZN(n212) );
  AOI22_X1 U195 ( .A1(multa[14]), .A2(n176), .B1(mul_w[14]), .B2(n116), .ZN(
        n162) );
  INV_X1 U196 ( .A(n162), .ZN(n213) );
  INV_X1 U197 ( .A(n163), .ZN(n214) );
  INV_X1 U198 ( .A(n164), .ZN(n215) );
  AOI22_X1 U199 ( .A1(multa[11]), .A2(n176), .B1(mul_w[11]), .B2(n116), .ZN(
        n165) );
  INV_X1 U200 ( .A(n165), .ZN(n216) );
  INV_X1 U201 ( .A(n166), .ZN(n217) );
  INV_X1 U202 ( .A(n167), .ZN(n218) );
  AOI22_X1 U203 ( .A1(multa[8]), .A2(n176), .B1(mul_w[8]), .B2(n116), .ZN(n168) );
  INV_X1 U204 ( .A(n168), .ZN(n219) );
  AOI22_X1 U205 ( .A1(multa[7]), .A2(n176), .B1(mul_w[7]), .B2(n116), .ZN(n169) );
  INV_X1 U206 ( .A(n169), .ZN(n220) );
  AOI22_X1 U207 ( .A1(multa[6]), .A2(n176), .B1(mul_w[6]), .B2(n116), .ZN(n170) );
  INV_X1 U208 ( .A(n170), .ZN(n221) );
  AOI22_X1 U209 ( .A1(multa[5]), .A2(n176), .B1(mul_w[5]), .B2(n116), .ZN(n171) );
  INV_X1 U210 ( .A(n171), .ZN(n222) );
  AOI22_X1 U211 ( .A1(multa[4]), .A2(n176), .B1(mul_w[4]), .B2(n116), .ZN(n172) );
  INV_X1 U212 ( .A(n172), .ZN(n223) );
  AOI22_X1 U213 ( .A1(multa[3]), .A2(n176), .B1(mul_w[3]), .B2(n116), .ZN(n173) );
  INV_X1 U214 ( .A(n173), .ZN(n224) );
  AOI22_X1 U215 ( .A1(multa[2]), .A2(n176), .B1(mul_w[2]), .B2(n116), .ZN(n174) );
  INV_X1 U216 ( .A(n174), .ZN(n225) );
  AOI22_X1 U217 ( .A1(multa[1]), .A2(n176), .B1(mul_w[1]), .B2(n116), .ZN(n175) );
  INV_X1 U218 ( .A(n175), .ZN(n226) );
  AOI22_X1 U219 ( .A1(multa[0]), .A2(n176), .B1(mul_w[0]), .B2(n116), .ZN(n177) );
  INV_X1 U220 ( .A(n177), .ZN(n227) );
  AOI22_X1 U221 ( .A1(f[0]), .A2(n178), .B1(N28), .B2(n115), .ZN(n179) );
  INV_X1 U222 ( .A(n179), .ZN(n196) );
endmodule

