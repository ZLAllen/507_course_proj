
module memory_WIDTH16_SIZE4_LOGSIZE3 ( clk, data_in, data_out, addr, wr_en );
  input [15:0] data_in;
  output [15:0] data_out;
  input [2:0] addr;
  input clk, wr_en;
  wire   N6, N7, \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] ,
         \mem[3][11] , \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] ,
         \mem[3][6] , \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] ,
         \mem[3][1] , \mem[3][0] , \mem[2][15] , \mem[2][14] , \mem[2][13] ,
         \mem[2][12] , \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] ,
         \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] ,
         \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][15] , \mem[1][14] ,
         \mem[1][13] , \mem[1][12] , \mem[1][11] , \mem[1][10] , \mem[1][9] ,
         \mem[1][8] , \mem[1][7] , \mem[1][6] , \mem[1][5] , \mem[1][4] ,
         \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] , \mem[0][15] ,
         \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] , \mem[0][10] ,
         \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] , \mem[0][5] ,
         \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N8,
         N9, N10, N11, N12, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n1, n4, n5, n6, n7, n8, n9, n12,
         n13, n14, n15, n16, n17, n18, n19, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211;
  assign N6 = addr[0];
  assign N7 = addr[1];

  DFF_X1 \data_out_reg[15]  ( .D(N8), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \data_out_reg[13]  ( .D(N10), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \data_out_reg[11]  ( .D(N12), .CK(clk), .QN(n9) );
  DFF_X1 \data_out_reg[5]  ( .D(N18), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[3]  ( .D(N20), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[1]  ( .D(N22), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N23), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[3][15]  ( .D(n152), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n151), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n150), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n149), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n148), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n147), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n146), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n145), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n144), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n143), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n142), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n141), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n140), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n139), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n138), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n137), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n136), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n135), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n134), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n133), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n132), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n131), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n130), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n129), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n128), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n127), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n126), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n125), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n124), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n123), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n122), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n121), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n120), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n119), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n118), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n117), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n116), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n115), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n114), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n113), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n112), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n111), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n110), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n109), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n108), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n107), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n106), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n105), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n104), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n103), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n102), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n101), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n100), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n99), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n98), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n97), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n96), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n95), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n94), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n93), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n92), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n91), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n90), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n89), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U151 ( .A1(n4), .A2(n195), .A3(n194), .ZN(n20) );
  NAND3_X1 U152 ( .A1(n4), .A2(n195), .A3(n193), .ZN(n38) );
  NAND3_X1 U153 ( .A1(n37), .A2(n194), .A3(N7), .ZN(n55) );
  NAND3_X1 U154 ( .A1(n37), .A2(n193), .A3(N7), .ZN(n72) );
  DFF_X1 \data_out_reg[4]  ( .D(N19), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N21), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[6]  ( .D(N17), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[8]  ( .D(N15), .CK(clk), .Q(data_out[8]) );
  SDFF_X2 \data_out_reg[10]  ( .D(n168), .SI(n167), .SE(N7), .CK(clk), .Q(
        data_out[10]) );
  DFF_X1 \data_out_reg[12]  ( .D(N11), .CK(clk), .Q(data_out[12]) );
  DFF_X2 \data_out_reg[14]  ( .D(N9), .CK(clk), .Q(data_out[14]) );
  DFF_X2 \data_out_reg[9]  ( .D(N14), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \data_out_reg[7]  ( .D(N16), .CK(clk), .QN(n1) );
  INV_X2 U3 ( .A(n1), .ZN(data_out[7]) );
  INV_X1 U4 ( .A(addr[2]), .ZN(n12) );
  BUF_X1 U5 ( .A(n20), .Z(n191) );
  AND2_X1 U6 ( .A1(wr_en), .A2(n12), .ZN(n4) );
  AND2_X1 U7 ( .A1(wr_en), .A2(n12), .ZN(n37) );
  BUF_X1 U8 ( .A(n55), .Z(n5) );
  BUF_X1 U9 ( .A(n55), .Z(n187) );
  BUF_X1 U10 ( .A(n38), .Z(n190) );
  BUF_X1 U11 ( .A(n72), .Z(n184) );
  BUF_X2 U12 ( .A(n20), .Z(n6) );
  BUF_X2 U13 ( .A(n72), .Z(n183) );
  BUF_X2 U14 ( .A(n72), .Z(n182) );
  BUF_X1 U15 ( .A(n38), .Z(n7) );
  BUF_X1 U16 ( .A(n38), .Z(n8) );
  INV_X2 U17 ( .A(n9), .ZN(data_out[11]) );
  BUF_X2 U18 ( .A(n55), .Z(n186) );
  BUF_X2 U19 ( .A(n55), .Z(n185) );
  BUF_X2 U20 ( .A(n20), .Z(n192) );
  BUF_X1 U21 ( .A(n72), .Z(n13) );
  BUF_X1 U22 ( .A(n38), .Z(n189) );
  BUF_X1 U23 ( .A(n38), .Z(n188) );
  BUF_X1 U24 ( .A(n193), .Z(n180) );
  BUF_X1 U25 ( .A(n193), .Z(n181) );
  BUF_X1 U26 ( .A(n193), .Z(n179) );
  INV_X1 U27 ( .A(N7), .ZN(n195) );
  INV_X1 U28 ( .A(data_in[0]), .ZN(n211) );
  INV_X1 U29 ( .A(data_in[1]), .ZN(n210) );
  INV_X1 U30 ( .A(data_in[2]), .ZN(n209) );
  INV_X1 U31 ( .A(data_in[3]), .ZN(n208) );
  INV_X1 U32 ( .A(data_in[4]), .ZN(n207) );
  INV_X1 U33 ( .A(data_in[5]), .ZN(n206) );
  INV_X1 U34 ( .A(data_in[6]), .ZN(n205) );
  INV_X1 U35 ( .A(data_in[7]), .ZN(n204) );
  INV_X1 U36 ( .A(data_in[8]), .ZN(n203) );
  INV_X1 U37 ( .A(data_in[9]), .ZN(n202) );
  INV_X1 U38 ( .A(data_in[10]), .ZN(n201) );
  INV_X1 U39 ( .A(data_in[11]), .ZN(n200) );
  INV_X1 U40 ( .A(data_in[12]), .ZN(n199) );
  INV_X1 U41 ( .A(data_in[13]), .ZN(n198) );
  INV_X1 U42 ( .A(data_in[14]), .ZN(n197) );
  INV_X1 U43 ( .A(data_in[15]), .ZN(n196) );
  OAI21_X1 U44 ( .B1(n204), .B2(n182), .A(n80), .ZN(n144) );
  NAND2_X1 U45 ( .A1(\mem[3][7] ), .A2(n183), .ZN(n80) );
  OAI21_X1 U46 ( .B1(n204), .B2(n186), .A(n63), .ZN(n128) );
  NAND2_X1 U47 ( .A1(\mem[2][7] ), .A2(n185), .ZN(n63) );
  OAI21_X1 U48 ( .B1(n204), .B2(n189), .A(n46), .ZN(n112) );
  NAND2_X1 U49 ( .A1(\mem[1][7] ), .A2(n7), .ZN(n46) );
  OAI21_X1 U50 ( .B1(n191), .B2(n203), .A(n29), .ZN(n97) );
  NAND2_X1 U51 ( .A1(\mem[0][8] ), .A2(n192), .ZN(n29) );
  OAI21_X1 U52 ( .B1(n6), .B2(n202), .A(n30), .ZN(n98) );
  NAND2_X1 U53 ( .A1(\mem[0][9] ), .A2(n192), .ZN(n30) );
  OAI21_X1 U54 ( .B1(n191), .B2(n201), .A(n31), .ZN(n99) );
  NAND2_X1 U55 ( .A1(\mem[0][10] ), .A2(n192), .ZN(n31) );
  OAI21_X1 U56 ( .B1(n6), .B2(n200), .A(n32), .ZN(n100) );
  NAND2_X1 U57 ( .A1(\mem[0][11] ), .A2(n192), .ZN(n32) );
  OAI21_X1 U58 ( .B1(n191), .B2(n199), .A(n33), .ZN(n101) );
  NAND2_X1 U59 ( .A1(\mem[0][12] ), .A2(n192), .ZN(n33) );
  OAI21_X1 U60 ( .B1(n6), .B2(n198), .A(n34), .ZN(n102) );
  NAND2_X1 U61 ( .A1(\mem[0][13] ), .A2(n6), .ZN(n34) );
  OAI21_X1 U62 ( .B1(n6), .B2(n197), .A(n35), .ZN(n103) );
  NAND2_X1 U63 ( .A1(\mem[0][14] ), .A2(n6), .ZN(n35) );
  OAI21_X1 U64 ( .B1(n191), .B2(n207), .A(n25), .ZN(n93) );
  NAND2_X1 U65 ( .A1(\mem[0][4] ), .A2(n6), .ZN(n25) );
  OAI21_X1 U66 ( .B1(n6), .B2(n206), .A(n26), .ZN(n94) );
  NAND2_X1 U67 ( .A1(\mem[0][5] ), .A2(n191), .ZN(n26) );
  OAI21_X1 U68 ( .B1(n192), .B2(n205), .A(n27), .ZN(n95) );
  NAND2_X1 U69 ( .A1(\mem[0][6] ), .A2(n6), .ZN(n27) );
  OAI21_X1 U70 ( .B1(n191), .B2(n204), .A(n28), .ZN(n96) );
  NAND2_X1 U71 ( .A1(\mem[0][7] ), .A2(n192), .ZN(n28) );
  OAI21_X1 U72 ( .B1(n6), .B2(n211), .A(n21), .ZN(n89) );
  NAND2_X1 U73 ( .A1(\mem[0][0] ), .A2(n192), .ZN(n21) );
  OAI21_X1 U74 ( .B1(n191), .B2(n210), .A(n22), .ZN(n90) );
  NAND2_X1 U75 ( .A1(\mem[0][1] ), .A2(n192), .ZN(n22) );
  OAI21_X1 U76 ( .B1(n6), .B2(n209), .A(n23), .ZN(n91) );
  NAND2_X1 U77 ( .A1(\mem[0][2] ), .A2(n192), .ZN(n23) );
  OAI21_X1 U78 ( .B1(n6), .B2(n208), .A(n24), .ZN(n92) );
  NAND2_X1 U79 ( .A1(\mem[0][3] ), .A2(n192), .ZN(n24) );
  OAI21_X1 U80 ( .B1(n6), .B2(n196), .A(n36), .ZN(n104) );
  NAND2_X1 U81 ( .A1(\mem[0][15] ), .A2(n192), .ZN(n36) );
  OAI21_X1 U82 ( .B1(n207), .B2(n182), .A(n77), .ZN(n141) );
  NAND2_X1 U83 ( .A1(\mem[3][4] ), .A2(n13), .ZN(n77) );
  OAI21_X1 U84 ( .B1(n206), .B2(n182), .A(n78), .ZN(n142) );
  NAND2_X1 U85 ( .A1(\mem[3][5] ), .A2(n182), .ZN(n78) );
  OAI21_X1 U86 ( .B1(n205), .B2(n183), .A(n79), .ZN(n143) );
  NAND2_X1 U87 ( .A1(\mem[3][6] ), .A2(n183), .ZN(n79) );
  OAI21_X1 U88 ( .B1(n207), .B2(n186), .A(n60), .ZN(n125) );
  NAND2_X1 U89 ( .A1(\mem[2][4] ), .A2(n185), .ZN(n60) );
  OAI21_X1 U90 ( .B1(n206), .B2(n5), .A(n61), .ZN(n126) );
  NAND2_X1 U91 ( .A1(\mem[2][5] ), .A2(n185), .ZN(n61) );
  OAI21_X1 U92 ( .B1(n205), .B2(n187), .A(n62), .ZN(n127) );
  NAND2_X1 U93 ( .A1(\mem[2][6] ), .A2(n185), .ZN(n62) );
  OAI21_X1 U94 ( .B1(n207), .B2(n7), .A(n43), .ZN(n109) );
  NAND2_X1 U95 ( .A1(\mem[1][4] ), .A2(n7), .ZN(n43) );
  OAI21_X1 U96 ( .B1(n206), .B2(n7), .A(n44), .ZN(n110) );
  NAND2_X1 U97 ( .A1(\mem[1][5] ), .A2(n189), .ZN(n44) );
  OAI21_X1 U98 ( .B1(n205), .B2(n189), .A(n45), .ZN(n111) );
  NAND2_X1 U99 ( .A1(\mem[1][6] ), .A2(n190), .ZN(n45) );
  OAI21_X1 U100 ( .B1(n211), .B2(n184), .A(n73), .ZN(n137) );
  NAND2_X1 U101 ( .A1(\mem[3][0] ), .A2(n183), .ZN(n73) );
  OAI21_X1 U102 ( .B1(n210), .B2(n183), .A(n74), .ZN(n138) );
  NAND2_X1 U103 ( .A1(\mem[3][1] ), .A2(n182), .ZN(n74) );
  OAI21_X1 U104 ( .B1(n209), .B2(n184), .A(n75), .ZN(n139) );
  NAND2_X1 U105 ( .A1(\mem[3][2] ), .A2(n13), .ZN(n75) );
  OAI21_X1 U106 ( .B1(n208), .B2(n182), .A(n76), .ZN(n140) );
  NAND2_X1 U107 ( .A1(\mem[3][3] ), .A2(n183), .ZN(n76) );
  OAI21_X1 U108 ( .B1(n196), .B2(n182), .A(n88), .ZN(n152) );
  NAND2_X1 U109 ( .A1(\mem[3][15] ), .A2(n13), .ZN(n88) );
  OAI21_X1 U110 ( .B1(n203), .B2(n183), .A(n81), .ZN(n145) );
  NAND2_X1 U111 ( .A1(\mem[3][8] ), .A2(n184), .ZN(n81) );
  OAI21_X1 U112 ( .B1(n202), .B2(n183), .A(n82), .ZN(n146) );
  NAND2_X1 U113 ( .A1(\mem[3][9] ), .A2(n182), .ZN(n82) );
  OAI21_X1 U114 ( .B1(n201), .B2(n183), .A(n83), .ZN(n147) );
  NAND2_X1 U115 ( .A1(\mem[3][10] ), .A2(n182), .ZN(n83) );
  OAI21_X1 U116 ( .B1(n200), .B2(n184), .A(n84), .ZN(n148) );
  NAND2_X1 U117 ( .A1(\mem[3][11] ), .A2(n182), .ZN(n84) );
  OAI21_X1 U118 ( .B1(n199), .B2(n184), .A(n85), .ZN(n149) );
  NAND2_X1 U119 ( .A1(\mem[3][12] ), .A2(n13), .ZN(n85) );
  OAI21_X1 U120 ( .B1(n198), .B2(n182), .A(n86), .ZN(n150) );
  NAND2_X1 U121 ( .A1(\mem[3][13] ), .A2(n13), .ZN(n86) );
  OAI21_X1 U122 ( .B1(n197), .B2(n184), .A(n87), .ZN(n151) );
  NAND2_X1 U123 ( .A1(\mem[3][14] ), .A2(n13), .ZN(n87) );
  OAI21_X1 U124 ( .B1(n211), .B2(n186), .A(n56), .ZN(n121) );
  NAND2_X1 U125 ( .A1(\mem[2][0] ), .A2(n5), .ZN(n56) );
  OAI21_X1 U126 ( .B1(n210), .B2(n186), .A(n57), .ZN(n122) );
  NAND2_X1 U127 ( .A1(\mem[2][1] ), .A2(n187), .ZN(n57) );
  OAI21_X1 U128 ( .B1(n209), .B2(n5), .A(n58), .ZN(n123) );
  NAND2_X1 U129 ( .A1(\mem[2][2] ), .A2(n186), .ZN(n58) );
  OAI21_X1 U130 ( .B1(n208), .B2(n187), .A(n59), .ZN(n124) );
  NAND2_X1 U131 ( .A1(\mem[2][3] ), .A2(n186), .ZN(n59) );
  OAI21_X1 U132 ( .B1(n196), .B2(n186), .A(n71), .ZN(n136) );
  NAND2_X1 U133 ( .A1(\mem[2][15] ), .A2(n186), .ZN(n71) );
  OAI21_X1 U134 ( .B1(n203), .B2(n5), .A(n64), .ZN(n129) );
  NAND2_X1 U135 ( .A1(\mem[2][8] ), .A2(n185), .ZN(n64) );
  OAI21_X1 U136 ( .B1(n202), .B2(n187), .A(n65), .ZN(n130) );
  NAND2_X1 U137 ( .A1(\mem[2][9] ), .A2(n185), .ZN(n65) );
  OAI21_X1 U138 ( .B1(n201), .B2(n186), .A(n66), .ZN(n131) );
  NAND2_X1 U139 ( .A1(\mem[2][10] ), .A2(n185), .ZN(n66) );
  OAI21_X1 U140 ( .B1(n200), .B2(n186), .A(n67), .ZN(n132) );
  NAND2_X1 U141 ( .A1(\mem[2][11] ), .A2(n185), .ZN(n67) );
  OAI21_X1 U142 ( .B1(n199), .B2(n186), .A(n68), .ZN(n133) );
  NAND2_X1 U143 ( .A1(\mem[2][12] ), .A2(n185), .ZN(n68) );
  OAI21_X1 U144 ( .B1(n198), .B2(n5), .A(n69), .ZN(n134) );
  NAND2_X1 U145 ( .A1(\mem[2][13] ), .A2(n185), .ZN(n69) );
  OAI21_X1 U146 ( .B1(n197), .B2(n187), .A(n70), .ZN(n135) );
  NAND2_X1 U147 ( .A1(\mem[2][14] ), .A2(n185), .ZN(n70) );
  OAI21_X1 U148 ( .B1(n211), .B2(n188), .A(n39), .ZN(n105) );
  NAND2_X1 U149 ( .A1(\mem[1][0] ), .A2(n188), .ZN(n39) );
  OAI21_X1 U150 ( .B1(n210), .B2(n189), .A(n40), .ZN(n106) );
  NAND2_X1 U155 ( .A1(\mem[1][1] ), .A2(n8), .ZN(n40) );
  OAI21_X1 U156 ( .B1(n209), .B2(n188), .A(n41), .ZN(n107) );
  NAND2_X1 U157 ( .A1(\mem[1][2] ), .A2(n188), .ZN(n41) );
  OAI21_X1 U158 ( .B1(n208), .B2(n190), .A(n42), .ZN(n108) );
  NAND2_X1 U159 ( .A1(\mem[1][3] ), .A2(n189), .ZN(n42) );
  OAI21_X1 U160 ( .B1(n196), .B2(n190), .A(n54), .ZN(n120) );
  NAND2_X1 U161 ( .A1(\mem[1][15] ), .A2(n190), .ZN(n54) );
  OAI21_X1 U162 ( .B1(n203), .B2(n190), .A(n47), .ZN(n113) );
  NAND2_X1 U163 ( .A1(\mem[1][8] ), .A2(n8), .ZN(n47) );
  OAI21_X1 U164 ( .B1(n202), .B2(n189), .A(n48), .ZN(n114) );
  NAND2_X1 U165 ( .A1(\mem[1][9] ), .A2(n8), .ZN(n48) );
  OAI21_X1 U166 ( .B1(n201), .B2(n188), .A(n49), .ZN(n115) );
  NAND2_X1 U167 ( .A1(\mem[1][10] ), .A2(n7), .ZN(n49) );
  OAI21_X1 U168 ( .B1(n200), .B2(n190), .A(n50), .ZN(n116) );
  NAND2_X1 U169 ( .A1(\mem[1][11] ), .A2(n8), .ZN(n50) );
  OAI21_X1 U170 ( .B1(n199), .B2(n7), .A(n51), .ZN(n117) );
  NAND2_X1 U171 ( .A1(\mem[1][12] ), .A2(n8), .ZN(n51) );
  OAI21_X1 U172 ( .B1(n198), .B2(n7), .A(n52), .ZN(n118) );
  NAND2_X1 U173 ( .A1(\mem[1][13] ), .A2(n189), .ZN(n52) );
  OAI21_X1 U174 ( .B1(n197), .B2(n188), .A(n53), .ZN(n119) );
  NAND2_X1 U175 ( .A1(\mem[1][14] ), .A2(n8), .ZN(n53) );
  MUX2_X1 U176 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n179), .Z(n14) );
  MUX2_X1 U177 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n179), .Z(n15) );
  MUX2_X1 U178 ( .A(n15), .B(n14), .S(N7), .Z(N23) );
  MUX2_X1 U179 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n179), .Z(n16) );
  MUX2_X1 U180 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n179), .Z(n17) );
  MUX2_X1 U181 ( .A(n17), .B(n16), .S(N7), .Z(N22) );
  MUX2_X1 U182 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n179), .Z(n18) );
  MUX2_X1 U183 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n179), .Z(n19) );
  MUX2_X1 U184 ( .A(n19), .B(n18), .S(N7), .Z(N21) );
  MUX2_X1 U185 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n179), .Z(n153) );
  MUX2_X1 U186 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n179), .Z(n154) );
  MUX2_X1 U187 ( .A(n154), .B(n153), .S(N7), .Z(N20) );
  MUX2_X1 U188 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n180), .Z(n155) );
  MUX2_X1 U189 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n180), .Z(n156) );
  MUX2_X1 U190 ( .A(n156), .B(n155), .S(N7), .Z(N19) );
  MUX2_X1 U191 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n180), .Z(n157) );
  MUX2_X1 U192 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n180), .Z(n158) );
  MUX2_X1 U193 ( .A(n158), .B(n157), .S(N7), .Z(N18) );
  MUX2_X1 U194 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n180), .Z(n159) );
  MUX2_X1 U195 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n180), .Z(n160) );
  MUX2_X1 U196 ( .A(n160), .B(n159), .S(N7), .Z(N17) );
  MUX2_X1 U197 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n180), .Z(n161) );
  MUX2_X1 U198 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n180), .Z(n162) );
  MUX2_X1 U199 ( .A(n162), .B(n161), .S(N7), .Z(N16) );
  MUX2_X1 U200 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n180), .Z(n163) );
  MUX2_X1 U201 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n180), .Z(n164) );
  MUX2_X1 U202 ( .A(n164), .B(n163), .S(N7), .Z(N15) );
  MUX2_X1 U203 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n180), .Z(n165) );
  MUX2_X1 U204 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n180), .Z(n166) );
  MUX2_X1 U205 ( .A(n166), .B(n165), .S(N7), .Z(N14) );
  MUX2_X1 U206 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n181), .Z(n167) );
  MUX2_X1 U207 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n181), .Z(n168) );
  MUX2_X1 U208 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n181), .Z(n169) );
  MUX2_X1 U209 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n181), .Z(n170) );
  MUX2_X1 U210 ( .A(n170), .B(n169), .S(N7), .Z(N12) );
  MUX2_X1 U211 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n181), .Z(n171) );
  MUX2_X1 U212 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n181), .Z(n172) );
  MUX2_X1 U213 ( .A(n172), .B(n171), .S(N7), .Z(N11) );
  MUX2_X1 U214 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n181), .Z(n173) );
  MUX2_X1 U215 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n181), .Z(n174) );
  MUX2_X1 U216 ( .A(n174), .B(n173), .S(N7), .Z(N10) );
  MUX2_X1 U217 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n181), .Z(n175) );
  MUX2_X1 U218 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n181), .Z(n176) );
  MUX2_X1 U219 ( .A(n176), .B(n175), .S(N7), .Z(N9) );
  MUX2_X1 U220 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(n181), .Z(n177) );
  MUX2_X1 U221 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(n181), .Z(n178) );
  MUX2_X1 U222 ( .A(n178), .B(n177), .S(N7), .Z(N8) );
  INV_X1 U223 ( .A(n194), .ZN(n193) );
  INV_X1 U224 ( .A(N6), .ZN(n194) );
endmodule


module layer1_8_4_8_16_W_rom_0 ( clk, addr, z );
  input [2:0] addr;
  output [15:0] z;
  input clk;
  wire   N14, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n1, n2, n4, n35, n36;
  assign z[1] = 1'b0;
  assign N14 = addr[0];

  DFF_X1 \z_reg[15]  ( .D(n34), .CK(clk), .Q(z[15]), .QN(n5) );
  DFF_X1 \z_reg[14]  ( .D(n33), .CK(clk), .Q(z[14]), .QN(n6) );
  DFF_X1 \z_reg[13]  ( .D(n32), .CK(clk), .Q(z[13]), .QN(n7) );
  DFF_X1 \z_reg[12]  ( .D(n31), .CK(clk), .Q(z[12]), .QN(n8) );
  DFF_X1 \z_reg[11]  ( .D(n30), .CK(clk), .Q(z[11]), .QN(n9) );
  DFF_X1 \z_reg[10]  ( .D(n29), .CK(clk), .Q(z[10]), .QN(n10) );
  DFF_X1 \z_reg[9]  ( .D(n28), .CK(clk), .Q(z[9]), .QN(n11) );
  DFF_X1 \z_reg[8]  ( .D(n27), .CK(clk), .Q(z[8]), .QN(n12) );
  DFF_X1 \z_reg[7]  ( .D(n26), .CK(clk), .Q(z[7]), .QN(n13) );
  DFF_X1 \z_reg[6]  ( .D(n25), .CK(clk), .Q(z[6]), .QN(n14) );
  DFF_X1 \z_reg[5]  ( .D(n24), .CK(clk), .Q(z[5]), .QN(n15) );
  DFF_X1 \z_reg[4]  ( .D(n23), .CK(clk), .Q(z[4]), .QN(n16) );
  DFF_X1 \z_reg[3]  ( .D(n22), .CK(clk), .Q(z[3]), .QN(n17) );
  DFF_X1 \z_reg[2]  ( .D(n21), .CK(clk), .Q(z[2]), .QN(n18) );
  DFF_X1 \z_reg[0]  ( .D(n20), .CK(clk), .Q(z[0]), .QN(n19) );
  INV_X1 U3 ( .A(addr[2]), .ZN(n36) );
  OAI21_X1 U4 ( .B1(n36), .B2(n8), .A(n3), .ZN(n31) );
  OAI21_X1 U5 ( .B1(n36), .B2(n7), .A(n3), .ZN(n32) );
  OAI21_X1 U6 ( .B1(n36), .B2(n6), .A(n3), .ZN(n33) );
  OAI21_X1 U7 ( .B1(n36), .B2(n5), .A(n3), .ZN(n34) );
  NAND2_X1 U8 ( .A1(N14), .A2(n36), .ZN(n3) );
  INV_X1 U9 ( .A(addr[1]), .ZN(n35) );
  NAND2_X1 U10 ( .A1(n36), .A2(n35), .ZN(n4) );
  MUX2_X1 U11 ( .A(N14), .B(n19), .S(addr[2]), .Z(n1) );
  NAND2_X1 U12 ( .A1(n4), .A2(n1), .ZN(n20) );
  OAI21_X1 U13 ( .B1(n18), .B2(n36), .A(n3), .ZN(n21) );
  OAI211_X1 U14 ( .C1(n17), .C2(n36), .A(n4), .B(n3), .ZN(n22) );
  MUX2_X1 U15 ( .A(n35), .B(n16), .S(addr[2]), .Z(n2) );
  NAND2_X1 U16 ( .A1(n3), .A2(n2), .ZN(n23) );
  OAI222_X1 U17 ( .A1(n3), .A2(n35), .B1(N14), .B2(n4), .C1(n15), .C2(n36), 
        .ZN(n24) );
  OAI21_X1 U18 ( .B1(n14), .B2(n36), .A(n3), .ZN(n25) );
  OAI21_X1 U19 ( .B1(n13), .B2(n36), .A(n3), .ZN(n26) );
  OAI21_X1 U20 ( .B1(n12), .B2(n36), .A(n3), .ZN(n27) );
  OAI21_X1 U21 ( .B1(n11), .B2(n36), .A(n3), .ZN(n28) );
  OAI21_X1 U23 ( .B1(n10), .B2(n36), .A(n3), .ZN(n29) );
  OAI21_X1 U24 ( .B1(n9), .B2(n36), .A(n3), .ZN(n30) );
endmodule


module layer1_8_4_8_16_B_rom_0 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b0;
  assign z[14] = 1'b0;
  assign z[13] = 1'b0;
  assign z[12] = 1'b0;
  assign z[11] = 1'b0;
  assign z[10] = 1'b0;
  assign z[9] = 1'b0;
  assign z[8] = 1'b0;
  assign z[7] = 1'b0;
  assign z[6] = 1'b0;
  assign z[5] = 1'b1;
  assign z[4] = 1'b1;
  assign z[3] = 1'b1;
  assign z[2] = 1'b1;
  assign z[1] = 1'b0;
  assign z[0] = 1'b1;

endmodule


module layer1_8_4_8_16_W_rom_1 ( clk, addr, z );
  input [2:0] addr;
  output [15:0] z;
  input clk;
  wire   n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n1, n2, n3, n4, n5, n6, n7, n22, n23, n24;
  assign z[15] = 1'b1;
  assign z[14] = 1'b1;
  assign z[13] = 1'b1;
  assign z[12] = 1'b1;
  assign z[11] = 1'b1;
  assign z[10] = 1'b1;
  assign z[9] = 1'b1;
  assign z[8] = 1'b1;
  assign z[7] = 1'b1;

  DFF_X1 \z_reg[6]  ( .D(n21), .CK(clk), .Q(z[6]), .QN(n8) );
  DFF_X1 \z_reg[5]  ( .D(n20), .CK(clk), .Q(z[5]), .QN(n9) );
  DFF_X1 \z_reg[4]  ( .D(n19), .CK(clk), .Q(z[4]), .QN(n10) );
  DFF_X1 \z_reg[3]  ( .D(n18), .CK(clk), .Q(z[3]), .QN(n11) );
  DFF_X1 \z_reg[2]  ( .D(n17), .CK(clk), .Q(z[2]), .QN(n12) );
  DFF_X1 \z_reg[1]  ( .D(n16), .CK(clk), .Q(z[1]), .QN(n13) );
  DFF_X1 \z_reg[0]  ( .D(n15), .CK(clk), .Q(z[0]), .QN(n14) );
  INV_X1 U3 ( .A(addr[0]), .ZN(n1) );
  INV_X1 U4 ( .A(addr[2]), .ZN(n24) );
  NAND2_X1 U5 ( .A1(n1), .A2(n24), .ZN(n23) );
  INV_X1 U6 ( .A(n23), .ZN(n2) );
  INV_X1 U7 ( .A(addr[1]), .ZN(n7) );
  NAND2_X1 U8 ( .A1(n2), .A2(n7), .ZN(n5) );
  NAND2_X1 U9 ( .A1(addr[1]), .A2(addr[0]), .ZN(n3) );
  MUX2_X1 U10 ( .A(n3), .B(n14), .S(addr[2]), .Z(n4) );
  NAND2_X1 U11 ( .A1(n5), .A2(n4), .ZN(n15) );
  NAND3_X1 U12 ( .A1(addr[0]), .A2(n24), .A3(n7), .ZN(n22) );
  OAI21_X1 U13 ( .B1(n13), .B2(n24), .A(n22), .ZN(n16) );
  OAI21_X1 U14 ( .B1(n12), .B2(n24), .A(n5), .ZN(n17) );
  MUX2_X1 U15 ( .A(addr[1]), .B(n11), .S(addr[2]), .Z(n6) );
  NAND2_X1 U16 ( .A1(n23), .A2(n6), .ZN(n18) );
  OAI221_X1 U26 ( .B1(n23), .B2(n7), .C1(n10), .C2(n24), .A(n22), .ZN(n19) );
  OAI21_X1 U27 ( .B1(n9), .B2(n24), .A(n22), .ZN(n20) );
  OAI21_X1 U28 ( .B1(n8), .B2(n24), .A(n23), .ZN(n21) );
endmodule


module layer1_8_4_8_16_B_rom_1 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b0;
  assign z[14] = 1'b0;
  assign z[13] = 1'b0;
  assign z[12] = 1'b0;
  assign z[11] = 1'b0;
  assign z[10] = 1'b0;
  assign z[9] = 1'b0;
  assign z[8] = 1'b0;
  assign z[7] = 1'b0;
  assign z[6] = 1'b1;
  assign z[5] = 1'b1;
  assign z[4] = 1'b1;
  assign z[3] = 1'b1;
  assign z[2] = 1'b1;
  assign z[1] = 1'b1;
  assign z[0] = 1'b0;

endmodule


module layer1_8_4_8_16_W_rom_2 ( clk, addr, z );
  input [2:0] addr;
  output [15:0] z;
  input clk;
  wire   n2, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n1, n3, n4, n5, n6, n39, n40, n41, n42;

  DFF_X1 \z_reg[15]  ( .D(n38), .CK(clk), .Q(z[15]), .QN(n7) );
  DFF_X1 \z_reg[14]  ( .D(n37), .CK(clk), .Q(z[14]), .QN(n8) );
  DFF_X1 \z_reg[13]  ( .D(n36), .CK(clk), .Q(z[13]), .QN(n9) );
  DFF_X1 \z_reg[12]  ( .D(n35), .CK(clk), .Q(z[12]), .QN(n10) );
  DFF_X1 \z_reg[11]  ( .D(n34), .CK(clk), .Q(z[11]), .QN(n11) );
  DFF_X1 \z_reg[10]  ( .D(n33), .CK(clk), .Q(z[10]), .QN(n12) );
  DFF_X1 \z_reg[9]  ( .D(n32), .CK(clk), .Q(z[9]), .QN(n13) );
  DFF_X1 \z_reg[8]  ( .D(n31), .CK(clk), .Q(z[8]), .QN(n14) );
  DFF_X1 \z_reg[7]  ( .D(n30), .CK(clk), .Q(z[7]), .QN(n15) );
  DFF_X1 \z_reg[6]  ( .D(n29), .CK(clk), .Q(z[6]), .QN(n16) );
  DFF_X1 \z_reg[5]  ( .D(n28), .CK(clk), .Q(z[5]), .QN(n17) );
  DFF_X1 \z_reg[4]  ( .D(n27), .CK(clk), .Q(z[4]), .QN(n18) );
  DFF_X1 \z_reg[3]  ( .D(n26), .CK(clk), .Q(z[3]), .QN(n19) );
  DFF_X1 \z_reg[2]  ( .D(n25), .CK(clk), .Q(z[2]), .QN(n20) );
  DFF_X1 \z_reg[1]  ( .D(n24), .CK(clk), .Q(z[1]), .QN(n21) );
  DFF_X1 \z_reg[0]  ( .D(n23), .CK(clk), .Q(z[0]), .QN(n22) );
  INV_X1 U3 ( .A(addr[2]), .ZN(n42) );
  OAI21_X1 U4 ( .B1(n42), .B2(n10), .A(n2), .ZN(n35) );
  OAI21_X1 U5 ( .B1(n42), .B2(n9), .A(n2), .ZN(n36) );
  OAI21_X1 U6 ( .B1(n42), .B2(n8), .A(n2), .ZN(n37) );
  OAI21_X1 U7 ( .B1(n42), .B2(n7), .A(n2), .ZN(n38) );
  NAND3_X1 U8 ( .A1(addr[0]), .A2(addr[1]), .A3(n42), .ZN(n2) );
  OAI21_X1 U9 ( .B1(n22), .B2(n42), .A(n2), .ZN(n23) );
  INV_X1 U10 ( .A(addr[0]), .ZN(n6) );
  NAND2_X1 U11 ( .A1(addr[1]), .A2(n6), .ZN(n4) );
  INV_X1 U12 ( .A(n4), .ZN(n39) );
  MUX2_X1 U13 ( .A(n39), .B(n21), .S(addr[2]), .Z(n1) );
  INV_X1 U14 ( .A(n1), .ZN(n24) );
  INV_X1 U15 ( .A(addr[1]), .ZN(n3) );
  NAND2_X1 U16 ( .A1(n42), .A2(n3), .ZN(n41) );
  OAI21_X1 U17 ( .B1(n20), .B2(n42), .A(n41), .ZN(n25) );
  MUX2_X1 U18 ( .A(n4), .B(n19), .S(addr[2]), .Z(n5) );
  OAI21_X1 U19 ( .B1(n6), .B2(n41), .A(n5), .ZN(n26) );
  OAI21_X1 U20 ( .B1(n18), .B2(n42), .A(n41), .ZN(n27) );
  MUX2_X1 U21 ( .A(n39), .B(n17), .S(addr[2]), .Z(n40) );
  INV_X1 U22 ( .A(n40), .ZN(n28) );
  OAI22_X1 U23 ( .A1(addr[0]), .A2(n41), .B1(n16), .B2(n42), .ZN(n29) );
  OAI21_X1 U24 ( .B1(n15), .B2(n42), .A(n2), .ZN(n30) );
  OAI21_X1 U25 ( .B1(n14), .B2(n42), .A(n2), .ZN(n31) );
  OAI21_X1 U26 ( .B1(n13), .B2(n42), .A(n2), .ZN(n32) );
  OAI21_X1 U27 ( .B1(n12), .B2(n42), .A(n2), .ZN(n33) );
  OAI21_X1 U28 ( .B1(n11), .B2(n42), .A(n2), .ZN(n34) );
endmodule


module layer1_8_4_8_16_B_rom_2 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b1;
  assign z[14] = 1'b1;
  assign z[13] = 1'b1;
  assign z[12] = 1'b1;
  assign z[11] = 1'b1;
  assign z[10] = 1'b1;
  assign z[9] = 1'b1;
  assign z[8] = 1'b1;
  assign z[7] = 1'b1;
  assign z[6] = 1'b0;
  assign z[5] = 1'b0;
  assign z[4] = 1'b1;
  assign z[3] = 1'b1;
  assign z[2] = 1'b0;
  assign z[1] = 1'b1;
  assign z[0] = 1'b0;

endmodule


module layer1_8_4_8_16_W_rom_3 ( clk, addr, z );
  input [2:0] addr;
  output [15:0] z;
  input clk;
  wire   N17, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n1, n2,
         n3, n4, n17;
  assign z[15] = 1'b1;
  assign z[14] = 1'b1;
  assign z[13] = 1'b1;
  assign z[12] = 1'b1;
  assign z[11] = 1'b1;
  assign z[10] = 1'b1;
  assign z[9] = 1'b1;
  assign z[8] = 1'b1;
  assign z[7] = 1'b1;
  assign z[1] = 1'b0;
  assign N17 = addr[0];

  DFF_X1 \z_reg[6]  ( .D(n16), .CK(clk), .Q(z[6]), .QN(n5) );
  DFF_X1 \z_reg[5]  ( .D(n15), .CK(clk), .Q(z[5]), .QN(n6) );
  DFF_X1 \z_reg[4]  ( .D(n14), .CK(clk), .Q(z[4]), .QN(n7) );
  DFF_X1 \z_reg[3]  ( .D(n13), .CK(clk), .Q(z[3]), .QN(n8) );
  DFF_X1 \z_reg[2]  ( .D(n12), .CK(clk), .Q(z[2]), .QN(n9) );
  DFF_X1 \z_reg[0]  ( .D(n11), .CK(clk), .Q(z[0]), .QN(n10) );
  INV_X1 U3 ( .A(addr[2]), .ZN(n17) );
  NAND2_X1 U4 ( .A1(N17), .A2(n17), .ZN(n3) );
  INV_X1 U5 ( .A(addr[1]), .ZN(n2) );
  OAI22_X1 U6 ( .A1(n3), .A2(n2), .B1(n10), .B2(n17), .ZN(n11) );
  MUX2_X1 U7 ( .A(N17), .B(n9), .S(addr[2]), .Z(n1) );
  INV_X1 U8 ( .A(n1), .ZN(n12) );
  NAND2_X1 U9 ( .A1(n17), .A2(n2), .ZN(n4) );
  OAI21_X1 U10 ( .B1(n8), .B2(n17), .A(n4), .ZN(n13) );
  OAI211_X1 U11 ( .C1(n7), .C2(n17), .A(n3), .B(n4), .ZN(n14) );
  OAI21_X1 U12 ( .B1(n6), .B2(n17), .A(n3), .ZN(n15) );
  OAI21_X1 U23 ( .B1(n5), .B2(n17), .A(n4), .ZN(n16) );
endmodule


module layer1_8_4_8_16_B_rom_3 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b1;
  assign z[14] = 1'b1;
  assign z[13] = 1'b1;
  assign z[12] = 1'b1;
  assign z[11] = 1'b1;
  assign z[10] = 1'b1;
  assign z[9] = 1'b1;
  assign z[8] = 1'b1;
  assign z[7] = 1'b1;
  assign z[6] = 1'b0;
  assign z[5] = 1'b0;
  assign z[4] = 1'b0;
  assign z[3] = 1'b1;
  assign z[2] = 1'b0;
  assign z[1] = 1'b1;
  assign z[0] = 1'b0;

endmodule


module layer1_8_4_8_16_W_rom_4 ( clk, addr, z );
  input [2:0] addr;
  output [15:0] z;
  input clk;
  wire   n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n1, n2, n3, n4, n5, n6, n7;

  DFF_X1 \z_reg[15]  ( .D(n40), .CK(clk), .Q(z[15]), .QN(n9) );
  DFF_X1 \z_reg[13]  ( .D(n38), .CK(clk), .Q(z[13]), .QN(n11) );
  DFF_X1 \z_reg[12]  ( .D(n37), .CK(clk), .Q(z[12]), .QN(n12) );
  DFF_X1 \z_reg[11]  ( .D(n36), .CK(clk), .Q(z[11]), .QN(n13) );
  DFF_X1 \z_reg[10]  ( .D(n35), .CK(clk), .Q(z[10]), .QN(n14) );
  DFF_X1 \z_reg[9]  ( .D(n34), .CK(clk), .Q(z[9]), .QN(n15) );
  DFF_X1 \z_reg[8]  ( .D(n33), .CK(clk), .Q(z[8]), .QN(n16) );
  DFF_X1 \z_reg[7]  ( .D(n32), .CK(clk), .Q(z[7]), .QN(n17) );
  DFF_X1 \z_reg[6]  ( .D(n31), .CK(clk), .Q(z[6]), .QN(n18) );
  DFF_X1 \z_reg[5]  ( .D(n30), .CK(clk), .Q(z[5]), .QN(n19) );
  DFF_X1 \z_reg[4]  ( .D(n29), .CK(clk), .Q(z[4]), .QN(n20) );
  DFF_X1 \z_reg[3]  ( .D(n28), .CK(clk), .Q(z[3]), .QN(n21) );
  DFF_X1 \z_reg[2]  ( .D(n27), .CK(clk), .Q(z[2]), .QN(n22) );
  DFF_X1 \z_reg[1]  ( .D(n26), .CK(clk), .Q(z[1]), .QN(n23) );
  DFF_X1 \z_reg[0]  ( .D(n25), .CK(clk), .Q(z[0]), .QN(n24) );
  NAND3_X1 U22 ( .A1(addr[0]), .A2(n7), .A3(addr[1]), .ZN(n8) );
  DFF_X1 \z_reg[14]  ( .D(n39), .CK(clk), .Q(z[14]), .QN(n10) );
  AND2_X1 U3 ( .A1(n8), .A2(n4), .ZN(n1) );
  INV_X1 U4 ( .A(addr[2]), .ZN(n7) );
  OAI21_X1 U5 ( .B1(n7), .B2(n12), .A(n1), .ZN(n37) );
  OAI21_X1 U6 ( .B1(n7), .B2(n11), .A(n1), .ZN(n38) );
  OAI21_X1 U7 ( .B1(n7), .B2(n10), .A(n1), .ZN(n39) );
  OAI21_X1 U8 ( .B1(n7), .B2(n9), .A(n1), .ZN(n40) );
  INV_X1 U9 ( .A(addr[1]), .ZN(n2) );
  INV_X1 U10 ( .A(addr[0]), .ZN(n3) );
  NAND3_X1 U11 ( .A1(n7), .A2(n2), .A3(n3), .ZN(n4) );
  NAND3_X1 U12 ( .A1(addr[0]), .A2(n7), .A3(n2), .ZN(n5) );
  NAND3_X1 U13 ( .A1(addr[1]), .A2(n7), .A3(n3), .ZN(n6) );
  OAI211_X1 U14 ( .C1(n24), .C2(n7), .A(n5), .B(n6), .ZN(n25) );
  OAI21_X1 U15 ( .B1(n23), .B2(n7), .A(n4), .ZN(n26) );
  OAI21_X1 U16 ( .B1(n22), .B2(n7), .A(n5), .ZN(n27) );
  OAI21_X1 U17 ( .B1(n21), .B2(n7), .A(n4), .ZN(n28) );
  OAI21_X1 U18 ( .B1(n20), .B2(n7), .A(n5), .ZN(n29) );
  OAI21_X1 U19 ( .B1(n19), .B2(n7), .A(n6), .ZN(n30) );
  OAI21_X1 U20 ( .B1(n18), .B2(n7), .A(n6), .ZN(n31) );
  OAI21_X1 U21 ( .B1(n17), .B2(n7), .A(n1), .ZN(n32) );
  OAI21_X1 U23 ( .B1(n16), .B2(n7), .A(n1), .ZN(n33) );
  OAI21_X1 U24 ( .B1(n15), .B2(n7), .A(n1), .ZN(n34) );
  OAI21_X1 U25 ( .B1(n14), .B2(n7), .A(n1), .ZN(n35) );
  OAI21_X1 U26 ( .B1(n13), .B2(n7), .A(n1), .ZN(n36) );
endmodule


module layer1_8_4_8_16_B_rom_4 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b1;
  assign z[14] = 1'b1;
  assign z[13] = 1'b1;
  assign z[12] = 1'b1;
  assign z[11] = 1'b1;
  assign z[10] = 1'b1;
  assign z[9] = 1'b1;
  assign z[8] = 1'b1;
  assign z[7] = 1'b1;
  assign z[6] = 1'b0;
  assign z[5] = 1'b1;
  assign z[4] = 1'b1;
  assign z[3] = 1'b1;
  assign z[2] = 1'b0;
  assign z[1] = 1'b0;
  assign z[0] = 1'b0;

endmodule


module layer1_8_4_8_16_W_rom_5 ( clk, addr, z );
  input [2:0] addr;
  output [15:0] z;
  input clk;
  wire   N16, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n1, n2, n3, n33, n34, n35, n36;
  assign z[3] = 1'b0;
  assign z[2] = 1'b1;
  assign N16 = addr[1];

  DFF_X1 \z_reg[15]  ( .D(n32), .CK(clk), .Q(z[15]), .QN(n5) );
  DFF_X1 \z_reg[14]  ( .D(n31), .CK(clk), .Q(z[14]), .QN(n6) );
  DFF_X1 \z_reg[13]  ( .D(n30), .CK(clk), .Q(z[13]), .QN(n7) );
  DFF_X1 \z_reg[12]  ( .D(n29), .CK(clk), .Q(z[12]), .QN(n8) );
  DFF_X1 \z_reg[11]  ( .D(n28), .CK(clk), .Q(z[11]), .QN(n9) );
  DFF_X1 \z_reg[10]  ( .D(n27), .CK(clk), .Q(z[10]), .QN(n10) );
  DFF_X1 \z_reg[9]  ( .D(n26), .CK(clk), .Q(z[9]), .QN(n11) );
  DFF_X1 \z_reg[8]  ( .D(n25), .CK(clk), .Q(z[8]), .QN(n12) );
  DFF_X1 \z_reg[7]  ( .D(n24), .CK(clk), .Q(z[7]), .QN(n13) );
  DFF_X1 \z_reg[6]  ( .D(n23), .CK(clk), .Q(z[6]), .QN(n14) );
  DFF_X1 \z_reg[5]  ( .D(n22), .CK(clk), .Q(z[5]), .QN(n15) );
  DFF_X1 \z_reg[4]  ( .D(n21), .CK(clk), .Q(z[4]), .QN(n16) );
  DFF_X1 \z_reg[1]  ( .D(n20), .CK(clk), .Q(z[1]), .QN(n17) );
  DFF_X1 \z_reg[0]  ( .D(n19), .CK(clk), .Q(z[0]), .QN(n18) );
  INV_X1 U3 ( .A(addr[2]), .ZN(n36) );
  OAI21_X1 U4 ( .B1(n36), .B2(n8), .A(n4), .ZN(n29) );
  OAI21_X1 U5 ( .B1(n36), .B2(n7), .A(n4), .ZN(n30) );
  OAI21_X1 U6 ( .B1(n36), .B2(n6), .A(n4), .ZN(n31) );
  OAI21_X1 U7 ( .B1(n36), .B2(n5), .A(n4), .ZN(n32) );
  INV_X1 U8 ( .A(N16), .ZN(n1) );
  NAND2_X1 U9 ( .A1(n36), .A2(n1), .ZN(n4) );
  NAND2_X1 U10 ( .A1(N16), .A2(n36), .ZN(n35) );
  INV_X1 U11 ( .A(addr[0]), .ZN(n33) );
  OAI22_X1 U12 ( .A1(n35), .A2(n33), .B1(n18), .B2(n36), .ZN(n19) );
  OAI21_X1 U13 ( .B1(addr[2]), .B2(n33), .A(n4), .ZN(n2) );
  INV_X1 U14 ( .A(n2), .ZN(n3) );
  OAI21_X1 U15 ( .B1(n17), .B2(n36), .A(n3), .ZN(n20) );
  OAI21_X1 U16 ( .B1(n16), .B2(n36), .A(n3), .ZN(n21) );
  MUX2_X1 U17 ( .A(n33), .B(n15), .S(addr[2]), .Z(n34) );
  NAND2_X1 U18 ( .A1(n35), .A2(n34), .ZN(n22) );
  OAI21_X1 U19 ( .B1(n14), .B2(n36), .A(n35), .ZN(n23) );
  OAI21_X1 U20 ( .B1(n13), .B2(n36), .A(n4), .ZN(n24) );
  OAI21_X1 U23 ( .B1(n12), .B2(n36), .A(n4), .ZN(n25) );
  OAI21_X1 U24 ( .B1(n11), .B2(n36), .A(n4), .ZN(n26) );
  OAI21_X1 U25 ( .B1(n10), .B2(n36), .A(n4), .ZN(n27) );
  OAI21_X1 U26 ( .B1(n9), .B2(n36), .A(n4), .ZN(n28) );
endmodule


module layer1_8_4_8_16_B_rom_5 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b1;
  assign z[14] = 1'b1;
  assign z[13] = 1'b1;
  assign z[12] = 1'b1;
  assign z[11] = 1'b1;
  assign z[10] = 1'b1;
  assign z[9] = 1'b1;
  assign z[8] = 1'b1;
  assign z[7] = 1'b1;
  assign z[6] = 1'b1;
  assign z[5] = 1'b1;
  assign z[4] = 1'b1;
  assign z[3] = 1'b0;
  assign z[2] = 1'b0;
  assign z[1] = 1'b1;
  assign z[0] = 1'b1;

endmodule


module layer1_8_4_8_16_W_rom_6 ( clk, addr, z );
  input [2:0] addr;
  output [15:0] z;
  input clk;
  wire   N17, n2, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n1, n3, n4, n5, n38, n39, n40, n41, n42, n43,
         n44;
  assign N17 = addr[0];

  DFF_X1 \z_reg[15]  ( .D(n37), .CK(clk), .Q(z[15]), .QN(n6) );
  DFF_X1 \z_reg[14]  ( .D(n36), .CK(clk), .Q(z[14]), .QN(n7) );
  DFF_X1 \z_reg[13]  ( .D(n35), .CK(clk), .Q(z[13]), .QN(n8) );
  DFF_X1 \z_reg[12]  ( .D(n34), .CK(clk), .Q(z[12]), .QN(n9) );
  DFF_X1 \z_reg[11]  ( .D(n33), .CK(clk), .Q(z[11]), .QN(n10) );
  DFF_X1 \z_reg[10]  ( .D(n32), .CK(clk), .Q(z[10]), .QN(n11) );
  DFF_X1 \z_reg[9]  ( .D(n31), .CK(clk), .Q(z[9]), .QN(n12) );
  DFF_X1 \z_reg[8]  ( .D(n30), .CK(clk), .Q(z[8]), .QN(n13) );
  DFF_X1 \z_reg[7]  ( .D(n29), .CK(clk), .Q(z[7]), .QN(n14) );
  DFF_X1 \z_reg[6]  ( .D(n28), .CK(clk), .Q(z[6]), .QN(n15) );
  DFF_X1 \z_reg[5]  ( .D(n27), .CK(clk), .Q(z[5]), .QN(n16) );
  DFF_X1 \z_reg[4]  ( .D(n26), .CK(clk), .Q(z[4]), .QN(n17) );
  DFF_X1 \z_reg[3]  ( .D(n25), .CK(clk), .Q(z[3]), .QN(n18) );
  DFF_X1 \z_reg[2]  ( .D(n24), .CK(clk), .Q(z[2]), .QN(n19) );
  DFF_X1 \z_reg[1]  ( .D(n23), .CK(clk), .Q(z[1]), .QN(n20) );
  DFF_X1 \z_reg[0]  ( .D(n22), .CK(clk), .Q(z[0]), .QN(n21) );
  AND2_X1 U3 ( .A1(N17), .A2(addr[1]), .ZN(n1) );
  INV_X1 U4 ( .A(addr[2]), .ZN(n44) );
  OAI21_X1 U5 ( .B1(n44), .B2(n9), .A(n2), .ZN(n34) );
  OAI21_X1 U6 ( .B1(n44), .B2(n8), .A(n2), .ZN(n35) );
  OAI21_X1 U7 ( .B1(n44), .B2(n7), .A(n2), .ZN(n36) );
  OAI21_X1 U8 ( .B1(n44), .B2(n6), .A(n2), .ZN(n37) );
  NAND2_X1 U9 ( .A1(n1), .A2(n44), .ZN(n2) );
  OAI21_X1 U10 ( .B1(n21), .B2(n44), .A(n2), .ZN(n22) );
  INV_X1 U11 ( .A(addr[1]), .ZN(n3) );
  INV_X1 U12 ( .A(N17), .ZN(n41) );
  NAND2_X1 U13 ( .A1(n3), .A2(n41), .ZN(n39) );
  INV_X1 U14 ( .A(n39), .ZN(n4) );
  MUX2_X1 U15 ( .A(n4), .B(n20), .S(addr[2]), .Z(n5) );
  INV_X1 U16 ( .A(n5), .ZN(n23) );
  MUX2_X1 U17 ( .A(n1), .B(n19), .S(addr[2]), .Z(n38) );
  INV_X1 U18 ( .A(n38), .ZN(n24) );
  MUX2_X1 U19 ( .A(n39), .B(n18), .S(addr[2]), .Z(n40) );
  NAND2_X1 U20 ( .A1(n2), .A2(n40), .ZN(n25) );
  MUX2_X1 U21 ( .A(n41), .B(n17), .S(addr[2]), .Z(n42) );
  INV_X1 U22 ( .A(n42), .ZN(n26) );
  OAI21_X1 U23 ( .B1(n16), .B2(n44), .A(n2), .ZN(n27) );
  MUX2_X1 U24 ( .A(N17), .B(n15), .S(addr[2]), .Z(n43) );
  INV_X1 U25 ( .A(n43), .ZN(n28) );
  OAI21_X1 U26 ( .B1(n14), .B2(n44), .A(n2), .ZN(n29) );
  OAI21_X1 U27 ( .B1(n13), .B2(n44), .A(n2), .ZN(n30) );
  OAI21_X1 U28 ( .B1(n12), .B2(n44), .A(n2), .ZN(n31) );
  OAI21_X1 U29 ( .B1(n11), .B2(n44), .A(n2), .ZN(n32) );
  OAI21_X1 U30 ( .B1(n10), .B2(n44), .A(n2), .ZN(n33) );
endmodule


module layer1_8_4_8_16_B_rom_6 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b1;
  assign z[14] = 1'b1;
  assign z[13] = 1'b1;
  assign z[12] = 1'b1;
  assign z[11] = 1'b1;
  assign z[10] = 1'b1;
  assign z[9] = 1'b1;
  assign z[8] = 1'b1;
  assign z[7] = 1'b1;
  assign z[6] = 1'b0;
  assign z[5] = 1'b0;
  assign z[4] = 1'b0;
  assign z[3] = 1'b1;
  assign z[2] = 1'b0;
  assign z[1] = 1'b1;
  assign z[0] = 1'b1;

endmodule


module layer1_8_4_8_16_W_rom_7 ( clk, addr, z );
  input [2:0] addr;
  output [15:0] z;
  input clk;
  wire   N14, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n1, n2, n3, n4, n5, n6, n7, n39, n40, n41, n42,
         n43;
  assign z[2] = 1'b1;
  assign N14 = addr[0];

  DFF_X1 \z_reg[15]  ( .D(n38), .CK(clk), .Q(z[15]), .QN(n9) );
  DFF_X1 \z_reg[14]  ( .D(n37), .CK(clk), .Q(z[14]), .QN(n10) );
  DFF_X1 \z_reg[13]  ( .D(n36), .CK(clk), .Q(z[13]), .QN(n11) );
  DFF_X1 \z_reg[12]  ( .D(n35), .CK(clk), .Q(z[12]), .QN(n12) );
  DFF_X1 \z_reg[11]  ( .D(n34), .CK(clk), .Q(z[11]), .QN(n13) );
  DFF_X1 \z_reg[10]  ( .D(n33), .CK(clk), .Q(z[10]), .QN(n14) );
  DFF_X1 \z_reg[9]  ( .D(n32), .CK(clk), .Q(z[9]), .QN(n15) );
  DFF_X1 \z_reg[8]  ( .D(n31), .CK(clk), .Q(z[8]), .QN(n16) );
  DFF_X1 \z_reg[7]  ( .D(n30), .CK(clk), .Q(z[7]), .QN(n17) );
  DFF_X1 \z_reg[6]  ( .D(n29), .CK(clk), .Q(z[6]), .QN(n18) );
  DFF_X1 \z_reg[5]  ( .D(n28), .CK(clk), .Q(z[5]), .QN(n19) );
  DFF_X1 \z_reg[4]  ( .D(n27), .CK(clk), .Q(z[4]), .QN(n20) );
  DFF_X1 \z_reg[3]  ( .D(n26), .CK(clk), .Q(z[3]), .QN(n21) );
  DFF_X1 \z_reg[1]  ( .D(n25), .CK(clk), .Q(z[1]), .QN(n22) );
  DFF_X1 \z_reg[0]  ( .D(n24), .CK(clk), .Q(z[0]), .QN(n23) );
  NAND3_X1 U22 ( .A1(n43), .A2(n42), .A3(addr[1]), .ZN(n8) );
  AND2_X1 U3 ( .A1(addr[1]), .A2(N14), .ZN(n1) );
  INV_X1 U4 ( .A(addr[2]), .ZN(n42) );
  INV_X1 U5 ( .A(n2), .ZN(n41) );
  OAI21_X1 U6 ( .B1(n42), .B2(n12), .A(n41), .ZN(n35) );
  OAI21_X1 U7 ( .B1(n42), .B2(n11), .A(n41), .ZN(n36) );
  OAI21_X1 U8 ( .B1(n42), .B2(n10), .A(n41), .ZN(n37) );
  OAI21_X1 U9 ( .B1(n42), .B2(n9), .A(n41), .ZN(n38) );
  NAND2_X1 U10 ( .A1(N14), .A2(n42), .ZN(n7) );
  OAI21_X1 U11 ( .B1(addr[1]), .B2(n7), .A(n8), .ZN(n2) );
  MUX2_X1 U12 ( .A(n1), .B(n23), .S(addr[2]), .Z(n3) );
  INV_X1 U13 ( .A(n3), .ZN(n24) );
  OAI21_X1 U14 ( .B1(n22), .B2(n42), .A(n7), .ZN(n25) );
  INV_X1 U15 ( .A(addr[1]), .ZN(n4) );
  MUX2_X1 U16 ( .A(n4), .B(n21), .S(addr[2]), .Z(n5) );
  NAND2_X1 U17 ( .A1(n7), .A2(n5), .ZN(n26) );
  MUX2_X1 U18 ( .A(addr[1]), .B(n20), .S(addr[2]), .Z(n6) );
  NAND2_X1 U19 ( .A1(n7), .A2(n6), .ZN(n27) );
  MUX2_X1 U20 ( .A(N14), .B(n19), .S(addr[2]), .Z(n39) );
  INV_X1 U21 ( .A(n39), .ZN(n28) );
  MUX2_X1 U23 ( .A(n1), .B(n18), .S(addr[2]), .Z(n40) );
  INV_X1 U24 ( .A(n40), .ZN(n29) );
  OAI21_X1 U25 ( .B1(n17), .B2(n42), .A(n41), .ZN(n30) );
  OAI21_X1 U27 ( .B1(n16), .B2(n42), .A(n41), .ZN(n31) );
  OAI21_X1 U28 ( .B1(n15), .B2(n42), .A(n41), .ZN(n32) );
  OAI21_X1 U29 ( .B1(n14), .B2(n42), .A(n41), .ZN(n33) );
  OAI21_X1 U30 ( .B1(n13), .B2(n42), .A(n41), .ZN(n34) );
  INV_X1 U31 ( .A(N14), .ZN(n43) );
endmodule


module layer1_8_4_8_16_B_rom_7 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b1;
  assign z[14] = 1'b1;
  assign z[13] = 1'b1;
  assign z[12] = 1'b1;
  assign z[11] = 1'b1;
  assign z[10] = 1'b1;
  assign z[9] = 1'b1;
  assign z[8] = 1'b1;
  assign z[7] = 1'b1;
  assign z[6] = 1'b0;
  assign z[5] = 1'b1;
  assign z[4] = 1'b0;
  assign z[3] = 1'b1;
  assign z[2] = 1'b1;
  assign z[1] = 1'b1;
  assign z[0] = 1'b1;

endmodule


module layer1_8_4_8_16_datapath_M8_N4_T16_P8_0_DW_mult_tc_1 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n9, n12, n13, n16, n18, n19, n21, n23, n25, n27, n29, n31,
         n32, n34, n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n62, n63, n64, n65, n67,
         n69, n70, n72, n73, n74, n75, n76, n77, n78, n79, n80, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n93, n95, n96, n97, n98, n99, n101,
         n103, n104, n105, n106, n107, n109, n111, n112, n113, n114, n115,
         n117, n119, n120, n122, n125, n127, n131, n135, n139, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n237, n241, n247, n249, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n418, n419, n420, n421, n422, n423, n424, n426, n427, n429,
         n432, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U148 ( .A(n265), .B(n144), .Z(n145) );
  XOR2_X1 U150 ( .A(n271), .B(n146), .Z(n147) );
  XOR2_X1 U152 ( .A(n301), .B(n148), .Z(n149) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n263), .CI(n291), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n317), .B(n252), .CO(n173), .S(n174) );
  FA_X1 U167 ( .A(n180), .B(n187), .CI(n178), .CO(n175), .S(n176) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U169 ( .A(n193), .B(n282), .CI(n191), .CO(n179), .S(n180) );
  FA_X1 U170 ( .A(n268), .B(n292), .CI(n274), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U172 ( .A(n197), .B(n190), .CI(n188), .CO(n185), .S(n186) );
  FA_X1 U173 ( .A(n199), .B(n201), .CI(n192), .CO(n187), .S(n188) );
  FA_X1 U174 ( .A(n275), .B(n293), .CI(n194), .CO(n189), .S(n190) );
  FA_X1 U175 ( .A(n305), .B(n253), .CI(n283), .CO(n191), .S(n192) );
  HA_X1 U176 ( .A(n319), .B(n269), .CO(n193), .S(n194) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U179 ( .A(n294), .B(n284), .CI(n276), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n320), .B(n270), .CI(n306), .CO(n201), .S(n202) );
  FA_X1 U181 ( .A(n208), .B(n213), .CI(n206), .CO(n203), .S(n204) );
  FA_X1 U182 ( .A(n215), .B(n307), .CI(n210), .CO(n205), .S(n206) );
  FA_X1 U183 ( .A(n285), .B(n254), .CI(n295), .CO(n207), .S(n208) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U185 ( .A(n216), .B(n219), .CI(n214), .CO(n211), .S(n212) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n322), .B(n278), .CI(n308), .CO(n215), .S(n216) );
  FA_X1 U188 ( .A(n225), .B(n222), .CI(n220), .CO(n217), .S(n218) );
  HA_X1 U190 ( .A(n287), .B(n323), .CO(n221), .S(n222) );
  FA_X1 U192 ( .A(n324), .B(n288), .CI(n310), .CO(n225), .S(n226) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  HA_X1 U194 ( .A(n311), .B(n325), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n312), .B(n300), .CI(n326), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  OAI21_X2 U414 ( .B1(n113), .B2(n115), .A(n114), .ZN(n112) );
  BUF_X2 U415 ( .A(n578), .Z(n498) );
  XNOR2_X1 U416 ( .A(n590), .B(a[12]), .ZN(n37) );
  BUF_X2 U417 ( .A(n578), .Z(n528) );
  NOR2_X1 U418 ( .A1(n218), .A2(n223), .ZN(n97) );
  INV_X1 U419 ( .A(n554), .ZN(n32) );
  OR2_X1 U420 ( .A1(n228), .A2(n231), .ZN(n490) );
  OR2_X1 U421 ( .A1(n329), .A2(n258), .ZN(n491) );
  BUF_X1 U422 ( .A(n255), .Z(n492) );
  OR2_X2 U423 ( .A1(n552), .A2(n249), .ZN(n493) );
  OR2_X1 U424 ( .A1(n552), .A2(n249), .ZN(n6) );
  CLKBUF_X1 U425 ( .A(n95), .Z(n494) );
  INV_X1 U426 ( .A(n577), .ZN(n495) );
  OR2_X2 U427 ( .A1(n534), .A2(n562), .ZN(n23) );
  CLKBUF_X1 U428 ( .A(n31), .Z(n496) );
  XNOR2_X1 U429 ( .A(n582), .B(a[4]), .ZN(n497) );
  CLKBUF_X1 U430 ( .A(n542), .Z(n501) );
  CLKBUF_X3 U431 ( .A(n578), .Z(n499) );
  INV_X1 U432 ( .A(n509), .ZN(n500) );
  INV_X1 U433 ( .A(n509), .ZN(n21) );
  OR2_X1 U434 ( .A1(n196), .A2(n203), .ZN(n502) );
  BUF_X1 U435 ( .A(n309), .Z(n503) );
  XNOR2_X1 U436 ( .A(n45), .B(n504), .ZN(product[12]) );
  AND2_X1 U437 ( .A1(n524), .A2(n79), .ZN(n504) );
  INV_X1 U438 ( .A(n241), .ZN(n505) );
  OR2_X2 U439 ( .A1(n534), .A2(n562), .ZN(n506) );
  AOI21_X1 U440 ( .B1(n104), .B2(n575), .A(n101), .ZN(n507) );
  XOR2_X1 U441 ( .A(n592), .B(a[14]), .Z(n508) );
  INV_X2 U442 ( .A(n593), .ZN(n592) );
  XNOR2_X1 U443 ( .A(n585), .B(a[6]), .ZN(n509) );
  OAI21_X1 U444 ( .B1(n99), .B2(n97), .A(n98), .ZN(n510) );
  XNOR2_X1 U445 ( .A(n589), .B(a[8]), .ZN(n429) );
  INV_X1 U446 ( .A(n589), .ZN(n588) );
  XOR2_X1 U447 ( .A(n170), .B(n172), .Z(n511) );
  XOR2_X1 U448 ( .A(n511), .B(n179), .Z(n166) );
  XOR2_X1 U449 ( .A(n177), .B(n168), .Z(n512) );
  XOR2_X1 U450 ( .A(n512), .B(n166), .Z(n164) );
  NAND2_X1 U451 ( .A1(n170), .A2(n172), .ZN(n513) );
  NAND2_X1 U452 ( .A1(n170), .A2(n179), .ZN(n514) );
  NAND2_X1 U453 ( .A1(n172), .A2(n179), .ZN(n515) );
  NAND3_X1 U454 ( .A1(n513), .A2(n514), .A3(n515), .ZN(n165) );
  NAND2_X1 U455 ( .A1(n177), .A2(n168), .ZN(n516) );
  NAND2_X1 U456 ( .A1(n177), .A2(n166), .ZN(n517) );
  NAND2_X1 U457 ( .A1(n168), .A2(n166), .ZN(n518) );
  NAND3_X1 U458 ( .A1(n516), .A2(n517), .A3(n518), .ZN(n163) );
  INV_X2 U459 ( .A(n582), .ZN(n581) );
  AOI21_X1 U460 ( .B1(n567), .B2(n112), .A(n109), .ZN(n519) );
  XOR2_X1 U461 ( .A(n205), .B(n200), .Z(n520) );
  XOR2_X1 U462 ( .A(n198), .B(n520), .Z(n196) );
  NAND2_X1 U463 ( .A1(n198), .A2(n205), .ZN(n521) );
  NAND2_X1 U464 ( .A1(n198), .A2(n200), .ZN(n522) );
  NAND2_X1 U465 ( .A1(n205), .A2(n200), .ZN(n523) );
  NAND3_X1 U466 ( .A1(n521), .A2(n522), .A3(n523), .ZN(n195) );
  OR2_X1 U467 ( .A1(n176), .A2(n185), .ZN(n524) );
  INV_X1 U468 ( .A(n585), .ZN(n583) );
  BUF_X1 U469 ( .A(n9), .Z(n572) );
  OR2_X1 U470 ( .A1(n550), .A2(n78), .ZN(n525) );
  BUF_X2 U471 ( .A(n9), .Z(n573) );
  OR2_X2 U472 ( .A1(n526), .A2(n554), .ZN(n34) );
  XNOR2_X1 U473 ( .A(n496), .B(a[10]), .ZN(n526) );
  CLKBUF_X1 U474 ( .A(n578), .Z(n527) );
  INV_X1 U475 ( .A(n579), .ZN(n578) );
  NOR2_X1 U476 ( .A1(n186), .A2(n195), .ZN(n529) );
  NOR2_X1 U477 ( .A1(n186), .A2(n195), .ZN(n82) );
  XNOR2_X1 U478 ( .A(n582), .B(a[2]), .ZN(n432) );
  XNOR2_X1 U479 ( .A(n586), .B(a[8]), .ZN(n530) );
  XOR2_X1 U480 ( .A(n585), .B(a[4]), .Z(n537) );
  BUF_X2 U481 ( .A(n588), .Z(n533) );
  INV_X1 U482 ( .A(n583), .ZN(n531) );
  XOR2_X1 U483 ( .A(n579), .B(a[2]), .Z(n9) );
  OAI21_X1 U484 ( .B1(n82), .B2(n86), .A(n83), .ZN(n532) );
  XOR2_X1 U485 ( .A(n587), .B(a[6]), .Z(n534) );
  AOI21_X1 U486 ( .B1(n510), .B2(n564), .A(n93), .ZN(n535) );
  OR2_X1 U487 ( .A1(n204), .A2(n211), .ZN(n536) );
  OR2_X1 U488 ( .A1(n537), .A2(n497), .ZN(n18) );
  OR2_X1 U489 ( .A1(n537), .A2(n497), .ZN(n538) );
  OR2_X1 U490 ( .A1(n537), .A2(n497), .ZN(n539) );
  OAI21_X1 U491 ( .B1(n91), .B2(n89), .A(n90), .ZN(n540) );
  INV_X1 U492 ( .A(n524), .ZN(n541) );
  XNOR2_X1 U493 ( .A(n586), .B(a[8]), .ZN(n27) );
  AOI21_X1 U494 ( .B1(n540), .B2(n80), .A(n532), .ZN(n542) );
  AOI21_X1 U495 ( .B1(n80), .B2(n88), .A(n532), .ZN(n45) );
  INV_X1 U496 ( .A(n587), .ZN(n555) );
  BUF_X2 U497 ( .A(n27), .Z(n543) );
  INV_X2 U498 ( .A(n551), .ZN(n16) );
  NAND2_X1 U499 ( .A1(n432), .A2(n572), .ZN(n544) );
  NAND2_X1 U500 ( .A1(n432), .A2(n572), .ZN(n545) );
  NAND2_X1 U501 ( .A1(n432), .A2(n572), .ZN(n12) );
  XOR2_X1 U502 ( .A(n229), .B(n298), .Z(n546) );
  XOR2_X1 U503 ( .A(n226), .B(n546), .Z(n224) );
  NAND2_X1 U504 ( .A1(n226), .A2(n229), .ZN(n547) );
  NAND2_X1 U505 ( .A1(n226), .A2(n298), .ZN(n548) );
  NAND2_X1 U506 ( .A1(n229), .A2(n298), .ZN(n549) );
  NAND3_X1 U507 ( .A1(n547), .A2(n548), .A3(n549), .ZN(n223) );
  NOR2_X1 U508 ( .A1(n164), .A2(n175), .ZN(n550) );
  NOR2_X1 U509 ( .A1(n164), .A2(n175), .ZN(n75) );
  INV_X1 U510 ( .A(n582), .ZN(n580) );
  XNOR2_X1 U511 ( .A(n582), .B(a[4]), .ZN(n551) );
  XNOR2_X1 U512 ( .A(n577), .B(n249), .ZN(n552) );
  CLKBUF_X1 U513 ( .A(n510), .Z(n553) );
  XNOR2_X1 U514 ( .A(n589), .B(a[10]), .ZN(n554) );
  OAI21_X1 U515 ( .B1(n89), .B2(n535), .A(n90), .ZN(n88) );
  INV_X1 U516 ( .A(n587), .ZN(n556) );
  INV_X1 U517 ( .A(n587), .ZN(n586) );
  NAND2_X2 U518 ( .A1(n429), .A2(n530), .ZN(n29) );
  INV_X2 U519 ( .A(n249), .ZN(n557) );
  XNOR2_X1 U520 ( .A(n297), .B(n558), .ZN(n220) );
  XNOR2_X1 U521 ( .A(n255), .B(n309), .ZN(n558) );
  INV_X1 U522 ( .A(n579), .ZN(n577) );
  NAND2_X1 U523 ( .A1(n297), .A2(n492), .ZN(n559) );
  NAND2_X1 U524 ( .A1(n297), .A2(n503), .ZN(n560) );
  NAND2_X1 U525 ( .A1(n492), .A2(n503), .ZN(n561) );
  NAND3_X1 U526 ( .A1(n559), .A2(n560), .A3(n561), .ZN(n219) );
  XNOR2_X1 U527 ( .A(n88), .B(n51), .ZN(product[10]) );
  XNOR2_X1 U528 ( .A(n585), .B(a[6]), .ZN(n562) );
  XNOR2_X1 U529 ( .A(n70), .B(n47), .ZN(product[14]) );
  NAND2_X1 U530 ( .A1(n563), .A2(n69), .ZN(n47) );
  AOI21_X1 U531 ( .B1(n563), .B2(n74), .A(n67), .ZN(n65) );
  INV_X1 U532 ( .A(n69), .ZN(n67) );
  INV_X1 U533 ( .A(n74), .ZN(n72) );
  AOI21_X1 U534 ( .B1(n96), .B2(n564), .A(n93), .ZN(n91) );
  INV_X1 U535 ( .A(n95), .ZN(n93) );
  NAND2_X1 U536 ( .A1(n502), .A2(n86), .ZN(n51) );
  NAND2_X1 U537 ( .A1(n536), .A2(n90), .ZN(n52) );
  OR2_X1 U538 ( .A1(n152), .A2(n163), .ZN(n563) );
  NAND2_X1 U539 ( .A1(n125), .A2(n76), .ZN(n48) );
  INV_X1 U540 ( .A(n550), .ZN(n125) );
  OAI21_X1 U541 ( .B1(n75), .B2(n79), .A(n76), .ZN(n74) );
  NAND2_X1 U542 ( .A1(n127), .A2(n83), .ZN(n50) );
  NOR2_X1 U543 ( .A1(n78), .A2(n550), .ZN(n73) );
  NAND2_X1 U544 ( .A1(n152), .A2(n163), .ZN(n69) );
  NAND2_X1 U545 ( .A1(n564), .A2(n494), .ZN(n53) );
  NOR2_X1 U546 ( .A1(n196), .A2(n203), .ZN(n85) );
  NAND2_X1 U547 ( .A1(n131), .A2(n98), .ZN(n54) );
  INV_X1 U548 ( .A(n97), .ZN(n131) );
  OAI21_X1 U549 ( .B1(n507), .B2(n97), .A(n98), .ZN(n96) );
  AOI21_X1 U550 ( .B1(n565), .B2(n120), .A(n117), .ZN(n115) );
  INV_X1 U551 ( .A(n119), .ZN(n117) );
  NOR2_X1 U552 ( .A1(n176), .A2(n185), .ZN(n78) );
  XOR2_X1 U553 ( .A(n58), .B(n115), .Z(product[3]) );
  NAND2_X1 U554 ( .A1(n135), .A2(n114), .ZN(n58) );
  INV_X1 U555 ( .A(n113), .ZN(n135) );
  INV_X1 U556 ( .A(n122), .ZN(n120) );
  XNOR2_X1 U557 ( .A(n57), .B(n112), .ZN(product[4]) );
  XNOR2_X1 U558 ( .A(n59), .B(n120), .ZN(product[2]) );
  NAND2_X1 U559 ( .A1(n565), .A2(n119), .ZN(n59) );
  NAND2_X1 U560 ( .A1(n176), .A2(n185), .ZN(n79) );
  NAND2_X1 U561 ( .A1(n164), .A2(n175), .ZN(n76) );
  OR2_X1 U562 ( .A1(n212), .A2(n217), .ZN(n564) );
  NAND2_X1 U563 ( .A1(n196), .A2(n203), .ZN(n86) );
  NAND2_X1 U564 ( .A1(n212), .A2(n217), .ZN(n95) );
  NAND2_X1 U565 ( .A1(n204), .A2(n211), .ZN(n90) );
  NAND2_X1 U566 ( .A1(n186), .A2(n195), .ZN(n83) );
  XNOR2_X1 U567 ( .A(n63), .B(n46), .ZN(product[15]) );
  NAND2_X1 U568 ( .A1(n566), .A2(n62), .ZN(n46) );
  NAND2_X1 U569 ( .A1(n73), .A2(n563), .ZN(n64) );
  OR2_X1 U570 ( .A1(n328), .A2(n314), .ZN(n565) );
  OR2_X1 U571 ( .A1(n151), .A2(n139), .ZN(n566) );
  NAND2_X1 U572 ( .A1(n228), .A2(n231), .ZN(n106) );
  OR2_X1 U573 ( .A1(n232), .A2(n233), .ZN(n567) );
  AND2_X1 U574 ( .A1(n491), .A2(n122), .ZN(product[1]) );
  OR2_X1 U575 ( .A1(n43), .A2(n495), .ZN(n409) );
  OR2_X1 U576 ( .A1(n576), .A2(n582), .ZN(n392) );
  AND2_X1 U577 ( .A1(n576), .A2(n241), .ZN(n278) );
  OAI22_X1 U578 ( .A1(n39), .A2(n593), .B1(n337), .B2(n37), .ZN(n252) );
  OR2_X1 U579 ( .A1(n576), .A2(n593), .ZN(n337) );
  XNOR2_X1 U580 ( .A(n533), .B(n43), .ZN(n352) );
  XNOR2_X1 U581 ( .A(n155), .B(n569), .ZN(n139) );
  XNOR2_X1 U582 ( .A(n153), .B(n141), .ZN(n569) );
  XNOR2_X1 U583 ( .A(n157), .B(n570), .ZN(n141) );
  XNOR2_X1 U584 ( .A(n145), .B(n143), .ZN(n570) );
  OAI22_X1 U585 ( .A1(n42), .A2(n594), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U586 ( .A1(n43), .A2(n594), .ZN(n332) );
  OAI22_X1 U587 ( .A1(n34), .A2(n343), .B1(n342), .B2(n32), .ZN(n269) );
  XNOR2_X1 U588 ( .A(n31), .B(n43), .ZN(n343) );
  XNOR2_X1 U589 ( .A(n159), .B(n571), .ZN(n142) );
  XNOR2_X1 U590 ( .A(n315), .B(n261), .ZN(n571) );
  OR2_X1 U591 ( .A1(n576), .A2(n531), .ZN(n377) );
  INV_X1 U592 ( .A(n37), .ZN(n237) );
  XNOR2_X1 U593 ( .A(n592), .B(n43), .ZN(n336) );
  XNOR2_X1 U594 ( .A(n584), .B(n43), .ZN(n376) );
  OAI22_X1 U595 ( .A1(n34), .A2(n342), .B1(n341), .B2(n32), .ZN(n268) );
  OAI22_X1 U596 ( .A1(n34), .A2(n341), .B1(n340), .B2(n32), .ZN(n267) );
  OAI22_X1 U597 ( .A1(n39), .A2(n336), .B1(n37), .B2(n335), .ZN(n263) );
  AND2_X1 U598 ( .A1(n576), .A2(n497), .ZN(n300) );
  INV_X1 U599 ( .A(n19), .ZN(n587) );
  INV_X1 U600 ( .A(n25), .ZN(n589) );
  AND2_X1 U601 ( .A1(n576), .A2(n237), .ZN(n264) );
  AND2_X1 U602 ( .A1(n509), .A2(n576), .ZN(n288) );
  AND2_X1 U603 ( .A1(n576), .A2(n554), .ZN(n270) );
  AND2_X1 U604 ( .A1(n576), .A2(n508), .ZN(n260) );
  OAI22_X1 U605 ( .A1(n39), .A2(n335), .B1(n37), .B2(n334), .ZN(n262) );
  OAI22_X1 U606 ( .A1(n34), .A2(n591), .B1(n344), .B2(n32), .ZN(n253) );
  INV_X1 U607 ( .A(n7), .ZN(n582) );
  INV_X1 U608 ( .A(n13), .ZN(n585) );
  OAI22_X1 U609 ( .A1(n34), .A2(n340), .B1(n339), .B2(n32), .ZN(n266) );
  AND2_X1 U610 ( .A1(n576), .A2(n247), .ZN(n314) );
  OR2_X1 U611 ( .A1(n43), .A2(n591), .ZN(n344) );
  AND2_X1 U612 ( .A1(n576), .A2(n249), .ZN(product[0]) );
  OR2_X1 U613 ( .A1(n43), .A2(n587), .ZN(n364) );
  OR2_X1 U614 ( .A1(n576), .A2(n589), .ZN(n353) );
  XNOR2_X1 U615 ( .A(n592), .B(a[14]), .ZN(n41) );
  OAI22_X1 U616 ( .A1(n39), .A2(n334), .B1(n37), .B2(n333), .ZN(n261) );
  XNOR2_X1 U617 ( .A(n592), .B(n422), .ZN(n333) );
  XNOR2_X1 U618 ( .A(n584), .B(b[11]), .ZN(n365) );
  OAI22_X1 U619 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U620 ( .A(n40), .B(n424), .ZN(n330) );
  XNOR2_X1 U621 ( .A(n40), .B(n43), .ZN(n331) );
  XNOR2_X1 U622 ( .A(n496), .B(n422), .ZN(n340) );
  XNOR2_X1 U623 ( .A(n590), .B(n423), .ZN(n341) );
  XNOR2_X1 U624 ( .A(n590), .B(n421), .ZN(n339) );
  XNOR2_X1 U625 ( .A(n31), .B(n424), .ZN(n342) );
  XNOR2_X1 U626 ( .A(n592), .B(n423), .ZN(n334) );
  XNOR2_X1 U627 ( .A(n592), .B(n424), .ZN(n335) );
  XNOR2_X1 U628 ( .A(n533), .B(n418), .ZN(n345) );
  OAI22_X1 U629 ( .A1(n34), .A2(n339), .B1(n338), .B2(n32), .ZN(n265) );
  XNOR2_X1 U630 ( .A(n496), .B(n420), .ZN(n338) );
  XNOR2_X1 U631 ( .A(n581), .B(b[13]), .ZN(n378) );
  NAND2_X1 U632 ( .A1(n427), .A2(n37), .ZN(n39) );
  XNOR2_X1 U633 ( .A(n581), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U634 ( .A(n581), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U635 ( .A(n581), .B(n418), .ZN(n384) );
  XNOR2_X1 U636 ( .A(n581), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U637 ( .A(n581), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U638 ( .A(n581), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U639 ( .A(n581), .B(n419), .ZN(n385) );
  XNOR2_X1 U640 ( .A(n584), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U641 ( .A(n584), .B(n418), .ZN(n369) );
  XNOR2_X1 U642 ( .A(n584), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U643 ( .A(n584), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U644 ( .A(n533), .B(n422), .ZN(n349) );
  XNOR2_X1 U645 ( .A(n588), .B(n423), .ZN(n350) );
  XNOR2_X1 U646 ( .A(n588), .B(n421), .ZN(n348) );
  XNOR2_X1 U647 ( .A(n588), .B(n420), .ZN(n347) );
  XNOR2_X1 U648 ( .A(n533), .B(n419), .ZN(n346) );
  XNOR2_X1 U649 ( .A(n528), .B(b[11]), .ZN(n397) );
  XNOR2_X1 U650 ( .A(n499), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U651 ( .A(n499), .B(b[13]), .ZN(n395) );
  XNOR2_X1 U652 ( .A(n498), .B(b[14]), .ZN(n394) );
  XNOR2_X1 U653 ( .A(n588), .B(n424), .ZN(n351) );
  NAND2_X1 U654 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U655 ( .A(n40), .B(a[14]), .Z(n426) );
  BUF_X1 U656 ( .A(n43), .Z(n576) );
  XNOR2_X1 U657 ( .A(n528), .B(b[15]), .ZN(n393) );
  NAND2_X1 U658 ( .A1(n328), .A2(n314), .ZN(n119) );
  XOR2_X1 U659 ( .A(n592), .B(a[12]), .Z(n427) );
  XNOR2_X1 U660 ( .A(n553), .B(n53), .ZN(product[8]) );
  XOR2_X1 U661 ( .A(n91), .B(n52), .Z(product[9]) );
  CLKBUF_X1 U662 ( .A(n507), .Z(n574) );
  INV_X1 U663 ( .A(n529), .ZN(n127) );
  NOR2_X1 U664 ( .A1(n529), .A2(n85), .ZN(n80) );
  NAND2_X1 U665 ( .A1(n218), .A2(n223), .ZN(n98) );
  AOI21_X1 U666 ( .B1(n575), .B2(n104), .A(n101), .ZN(n99) );
  OR2_X1 U667 ( .A1(n224), .A2(n227), .ZN(n575) );
  OAI21_X1 U668 ( .B1(n105), .B2(n107), .A(n106), .ZN(n104) );
  NAND2_X1 U669 ( .A1(n567), .A2(n111), .ZN(n57) );
  NAND2_X1 U670 ( .A1(n232), .A2(n233), .ZN(n111) );
  XNOR2_X1 U671 ( .A(n84), .B(n50), .ZN(product[11]) );
  NAND2_X1 U672 ( .A1(n329), .A2(n258), .ZN(n122) );
  NOR2_X1 U673 ( .A1(n204), .A2(n211), .ZN(n89) );
  OAI22_X1 U674 ( .A1(n29), .A2(n346), .B1(n345), .B2(n543), .ZN(n271) );
  OAI22_X1 U675 ( .A1(n29), .A2(n350), .B1(n349), .B2(n543), .ZN(n275) );
  OAI22_X1 U676 ( .A1(n29), .A2(n347), .B1(n346), .B2(n543), .ZN(n272) );
  OAI22_X1 U677 ( .A1(n29), .A2(n348), .B1(n347), .B2(n543), .ZN(n273) );
  OAI22_X1 U678 ( .A1(n29), .A2(n351), .B1(n350), .B2(n543), .ZN(n276) );
  OAI22_X1 U679 ( .A1(n29), .A2(n349), .B1(n348), .B2(n543), .ZN(n274) );
  OAI22_X1 U680 ( .A1(n29), .A2(n589), .B1(n353), .B2(n543), .ZN(n254) );
  XNOR2_X1 U681 ( .A(n555), .B(n419), .ZN(n357) );
  INV_X1 U682 ( .A(n27), .ZN(n241) );
  XNOR2_X1 U683 ( .A(n556), .B(n418), .ZN(n356) );
  OAI22_X1 U684 ( .A1(n29), .A2(n352), .B1(n351), .B2(n505), .ZN(n277) );
  XNOR2_X1 U685 ( .A(n555), .B(n43), .ZN(n363) );
  XNOR2_X1 U686 ( .A(n555), .B(b[9]), .ZN(n354) );
  XNOR2_X1 U687 ( .A(n556), .B(n422), .ZN(n360) );
  XNOR2_X1 U688 ( .A(n555), .B(n423), .ZN(n361) );
  XNOR2_X1 U689 ( .A(n556), .B(b[8]), .ZN(n355) );
  XNOR2_X1 U690 ( .A(n556), .B(n424), .ZN(n362) );
  XNOR2_X1 U691 ( .A(n555), .B(n420), .ZN(n358) );
  XNOR2_X1 U692 ( .A(n556), .B(n421), .ZN(n359) );
  OAI22_X1 U693 ( .A1(n493), .A2(n395), .B1(n394), .B2(n557), .ZN(n316) );
  OAI22_X1 U694 ( .A1(n493), .A2(n394), .B1(n393), .B2(n557), .ZN(n315) );
  OAI22_X1 U695 ( .A1(n493), .A2(n397), .B1(n396), .B2(n557), .ZN(n318) );
  OAI22_X1 U696 ( .A1(n493), .A2(n396), .B1(n395), .B2(n557), .ZN(n317) );
  OAI22_X1 U697 ( .A1(n493), .A2(n398), .B1(n397), .B2(n557), .ZN(n319) );
  OAI22_X1 U698 ( .A1(n6), .A2(n402), .B1(n401), .B2(n557), .ZN(n323) );
  OAI22_X1 U699 ( .A1(n6), .A2(n406), .B1(n405), .B2(n557), .ZN(n327) );
  OAI22_X1 U700 ( .A1(n399), .A2(n493), .B1(n398), .B2(n557), .ZN(n320) );
  OAI22_X1 U701 ( .A1(n6), .A2(n401), .B1(n400), .B2(n557), .ZN(n322) );
  OAI22_X1 U702 ( .A1(n493), .A2(n403), .B1(n402), .B2(n557), .ZN(n324) );
  OAI22_X1 U703 ( .A1(n6), .A2(n404), .B1(n403), .B2(n557), .ZN(n325) );
  OAI22_X1 U704 ( .A1(n493), .A2(n400), .B1(n399), .B2(n557), .ZN(n321) );
  OAI22_X1 U705 ( .A1(n493), .A2(n405), .B1(n404), .B2(n557), .ZN(n326) );
  OAI22_X1 U706 ( .A1(n493), .A2(n407), .B1(n406), .B2(n557), .ZN(n328) );
  OAI22_X1 U707 ( .A1(n493), .A2(n408), .B1(n407), .B2(n557), .ZN(n329) );
  OAI22_X1 U708 ( .A1(n6), .A2(n495), .B1(n409), .B2(n557), .ZN(n258) );
  NOR2_X1 U709 ( .A1(n228), .A2(n231), .ZN(n105) );
  NAND2_X1 U710 ( .A1(n490), .A2(n106), .ZN(n56) );
  OAI21_X1 U711 ( .B1(n87), .B2(n85), .A(n86), .ZN(n84) );
  INV_X1 U712 ( .A(n540), .ZN(n87) );
  NAND2_X1 U713 ( .A1(n151), .A2(n139), .ZN(n62) );
  OAI22_X1 U714 ( .A1(n506), .A2(n358), .B1(n357), .B2(n500), .ZN(n282) );
  OAI22_X1 U715 ( .A1(n506), .A2(n356), .B1(n355), .B2(n500), .ZN(n280) );
  OAI22_X1 U716 ( .A1(n506), .A2(n362), .B1(n361), .B2(n500), .ZN(n286) );
  OAI22_X1 U717 ( .A1(n506), .A2(n360), .B1(n359), .B2(n500), .ZN(n284) );
  OAI22_X1 U718 ( .A1(n506), .A2(n357), .B1(n356), .B2(n500), .ZN(n281) );
  OAI22_X1 U719 ( .A1(n506), .A2(n361), .B1(n360), .B2(n500), .ZN(n285) );
  OAI22_X1 U720 ( .A1(n23), .A2(n363), .B1(n362), .B2(n21), .ZN(n287) );
  OAI22_X1 U721 ( .A1(n23), .A2(n587), .B1(n364), .B2(n21), .ZN(n255) );
  OAI22_X1 U722 ( .A1(n359), .A2(n23), .B1(n358), .B2(n21), .ZN(n283) );
  XNOR2_X1 U723 ( .A(n583), .B(n421), .ZN(n372) );
  XNOR2_X1 U724 ( .A(n583), .B(n424), .ZN(n375) );
  XNOR2_X1 U725 ( .A(n583), .B(n419), .ZN(n370) );
  XNOR2_X1 U726 ( .A(n583), .B(n420), .ZN(n371) );
  OAI22_X1 U727 ( .A1(n506), .A2(n355), .B1(n354), .B2(n500), .ZN(n279) );
  XNOR2_X1 U728 ( .A(n583), .B(n423), .ZN(n374) );
  XNOR2_X1 U729 ( .A(n583), .B(n422), .ZN(n373) );
  XNOR2_X1 U730 ( .A(n77), .B(n48), .ZN(product[13]) );
  NOR2_X1 U731 ( .A1(n234), .A2(n257), .ZN(n113) );
  NAND2_X1 U732 ( .A1(n224), .A2(n227), .ZN(n103) );
  INV_X1 U733 ( .A(n103), .ZN(n101) );
  NAND2_X1 U734 ( .A1(n575), .A2(n103), .ZN(n55) );
  INV_X1 U735 ( .A(n1), .ZN(n579) );
  OAI22_X1 U736 ( .A1(n539), .A2(n370), .B1(n369), .B2(n16), .ZN(n293) );
  OAI22_X1 U737 ( .A1(n538), .A2(n367), .B1(n366), .B2(n16), .ZN(n290) );
  OAI22_X1 U738 ( .A1(n538), .A2(n368), .B1(n367), .B2(n16), .ZN(n291) );
  OAI22_X1 U739 ( .A1(n539), .A2(n375), .B1(n374), .B2(n16), .ZN(n298) );
  OAI22_X1 U740 ( .A1(n18), .A2(n371), .B1(n370), .B2(n16), .ZN(n294) );
  OAI22_X1 U741 ( .A1(n539), .A2(n372), .B1(n371), .B2(n16), .ZN(n295) );
  OAI22_X1 U742 ( .A1(n539), .A2(n369), .B1(n368), .B2(n16), .ZN(n292) );
  OAI22_X1 U743 ( .A1(n539), .A2(n531), .B1(n377), .B2(n16), .ZN(n256) );
  OAI22_X1 U744 ( .A1(n538), .A2(n376), .B1(n375), .B2(n16), .ZN(n299) );
  OAI22_X1 U745 ( .A1(n538), .A2(n373), .B1(n372), .B2(n16), .ZN(n296) );
  OAI22_X1 U746 ( .A1(n538), .A2(n374), .B1(n373), .B2(n16), .ZN(n297) );
  OAI22_X1 U747 ( .A1(n18), .A2(n366), .B1(n365), .B2(n16), .ZN(n289) );
  XNOR2_X1 U748 ( .A(n580), .B(n420), .ZN(n386) );
  XNOR2_X1 U749 ( .A(n580), .B(n43), .ZN(n391) );
  XNOR2_X1 U750 ( .A(n580), .B(n423), .ZN(n389) );
  XNOR2_X1 U751 ( .A(n580), .B(n422), .ZN(n388) );
  XNOR2_X1 U752 ( .A(n580), .B(n424), .ZN(n390) );
  XNOR2_X1 U753 ( .A(n580), .B(n421), .ZN(n387) );
  XOR2_X1 U754 ( .A(n574), .B(n54), .Z(product[7]) );
  XNOR2_X1 U755 ( .A(n498), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U756 ( .A(n498), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U757 ( .A(n528), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U758 ( .A(n528), .B(n418), .ZN(n401) );
  XNOR2_X1 U759 ( .A(n498), .B(n419), .ZN(n402) );
  XNOR2_X1 U760 ( .A(n499), .B(n43), .ZN(n408) );
  XNOR2_X1 U761 ( .A(n528), .B(n422), .ZN(n405) );
  XNOR2_X1 U762 ( .A(n499), .B(n423), .ZN(n406) );
  XNOR2_X1 U763 ( .A(n527), .B(n420), .ZN(n403) );
  XNOR2_X1 U764 ( .A(n527), .B(n421), .ZN(n404) );
  XNOR2_X1 U765 ( .A(n499), .B(n424), .ZN(n407) );
  OAI21_X1 U766 ( .B1(n64), .B2(n501), .A(n65), .ZN(n63) );
  OAI21_X1 U767 ( .B1(n542), .B2(n525), .A(n72), .ZN(n70) );
  OAI21_X1 U768 ( .B1(n45), .B2(n541), .A(n79), .ZN(n77) );
  XNOR2_X1 U769 ( .A(n104), .B(n55), .ZN(product[6]) );
  XOR2_X1 U770 ( .A(n56), .B(n519), .Z(product[5]) );
  AOI21_X1 U771 ( .B1(n567), .B2(n112), .A(n109), .ZN(n107) );
  INV_X1 U772 ( .A(n111), .ZN(n109) );
  OAI22_X1 U773 ( .A1(n544), .A2(n379), .B1(n378), .B2(n573), .ZN(n301) );
  OAI22_X1 U774 ( .A1(n545), .A2(n380), .B1(n379), .B2(n573), .ZN(n302) );
  OAI22_X1 U775 ( .A1(n544), .A2(n385), .B1(n384), .B2(n573), .ZN(n307) );
  OAI22_X1 U776 ( .A1(n544), .A2(n382), .B1(n381), .B2(n573), .ZN(n304) );
  OAI22_X1 U777 ( .A1(n545), .A2(n381), .B1(n380), .B2(n573), .ZN(n303) );
  NAND2_X1 U778 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U779 ( .A1(n12), .A2(n383), .B1(n382), .B2(n573), .ZN(n305) );
  OAI22_X1 U780 ( .A1(n545), .A2(n384), .B1(n383), .B2(n573), .ZN(n306) );
  OAI22_X1 U781 ( .A1(n544), .A2(n386), .B1(n385), .B2(n573), .ZN(n308) );
  OAI22_X1 U782 ( .A1(n544), .A2(n387), .B1(n386), .B2(n573), .ZN(n309) );
  OAI22_X1 U783 ( .A1(n545), .A2(n582), .B1(n392), .B2(n573), .ZN(n257) );
  OAI22_X1 U784 ( .A1(n12), .A2(n389), .B1(n573), .B2(n388), .ZN(n311) );
  OAI22_X1 U785 ( .A1(n544), .A2(n388), .B1(n387), .B2(n573), .ZN(n310) );
  OAI22_X1 U786 ( .A1(n12), .A2(n390), .B1(n573), .B2(n389), .ZN(n312) );
  INV_X1 U787 ( .A(n573), .ZN(n247) );
  OAI22_X1 U788 ( .A1(n545), .A2(n391), .B1(n390), .B2(n573), .ZN(n313) );
  INV_X1 U789 ( .A(n585), .ZN(n584) );
  INV_X1 U790 ( .A(n591), .ZN(n590) );
  INV_X1 U791 ( .A(n31), .ZN(n591) );
  INV_X1 U792 ( .A(n36), .ZN(n593) );
  INV_X1 U793 ( .A(n40), .ZN(n594) );
  XOR2_X1 U794 ( .A(n259), .B(n251), .Z(n148) );
  XOR2_X1 U795 ( .A(n289), .B(n279), .Z(n146) );
  XOR2_X1 U796 ( .A(n149), .B(n147), .Z(n144) );
endmodule


module layer1_8_4_8_16_datapath_M8_N4_T16_P8_0_DW01_add_2 ( A, B, CI, SUM, CO
 );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n18,
         n19, n20, n21, n25, n26, n27, n28, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n46, n48, n49, n51, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n71, n72, n73,
         n74, n75, n77, n79, n80, n81, n82, n83, n85, n87, n88, n90, n98, n99,
         n100, n102, n104, n161, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186;

  OR2_X1 U126 ( .A1(A[11]), .A2(B[11]), .ZN(n161) );
  AND2_X1 U127 ( .A1(n178), .A2(n90), .ZN(SUM[0]) );
  NOR2_X1 U128 ( .A1(A[8]), .A2(B[8]), .ZN(n163) );
  NOR2_X1 U129 ( .A1(A[8]), .A2(B[8]), .ZN(n164) );
  NOR2_X1 U130 ( .A1(A[8]), .A2(B[8]), .ZN(n58) );
  XNOR2_X1 U131 ( .A(n41), .B(n165), .ZN(SUM[11]) );
  AND2_X1 U132 ( .A1(n161), .A2(n40), .ZN(n165) );
  OR2_X1 U133 ( .A1(A[15]), .A2(B[15]), .ZN(n166) );
  NOR2_X1 U134 ( .A1(n164), .A2(n61), .ZN(n167) );
  OR2_X1 U135 ( .A1(A[13]), .A2(B[13]), .ZN(n168) );
  OAI21_X1 U136 ( .B1(n163), .B2(n62), .A(n59), .ZN(n169) );
  OAI21_X1 U137 ( .B1(n164), .B2(n62), .A(n59), .ZN(n170) );
  AOI21_X1 U138 ( .B1(n183), .B2(n51), .A(n46), .ZN(n171) );
  AND2_X1 U139 ( .A1(A[13]), .A2(B[13]), .ZN(n172) );
  OR2_X2 U140 ( .A1(A[14]), .A2(B[14]), .ZN(n184) );
  AOI21_X1 U141 ( .B1(n167), .B2(n64), .A(n169), .ZN(n173) );
  AOI21_X1 U142 ( .B1(n56), .B2(n64), .A(n170), .ZN(n174) );
  OAI21_X1 U143 ( .B1(n43), .B2(n173), .A(n171), .ZN(n175) );
  NOR2_X1 U144 ( .A1(A[12]), .A2(B[12]), .ZN(n176) );
  AOI21_X1 U145 ( .B1(n175), .B2(n34), .A(n35), .ZN(n177) );
  OR2_X1 U146 ( .A1(A[0]), .A2(B[0]), .ZN(n178) );
  INV_X1 U147 ( .A(n64), .ZN(n63) );
  INV_X1 U148 ( .A(n174), .ZN(n54) );
  INV_X1 U149 ( .A(n42), .ZN(n41) );
  OAI21_X1 U150 ( .B1(n75), .B2(n73), .A(n74), .ZN(n72) );
  AOI21_X1 U151 ( .B1(n181), .B2(n88), .A(n85), .ZN(n83) );
  INV_X1 U152 ( .A(n87), .ZN(n85) );
  OAI21_X1 U153 ( .B1(n83), .B2(n81), .A(n82), .ZN(n80) );
  AOI21_X1 U154 ( .B1(n182), .B2(n80), .A(n77), .ZN(n75) );
  INV_X1 U155 ( .A(n79), .ZN(n77) );
  AOI21_X1 U156 ( .B1(n56), .B2(n64), .A(n57), .ZN(n55) );
  AOI21_X1 U157 ( .B1(n179), .B2(n72), .A(n69), .ZN(n67) );
  INV_X1 U158 ( .A(n71), .ZN(n69) );
  AOI21_X1 U159 ( .B1(n54), .B2(n180), .A(n51), .ZN(n49) );
  INV_X1 U160 ( .A(n90), .ZN(n88) );
  OAI21_X1 U161 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  INV_X1 U162 ( .A(n53), .ZN(n51) );
  NAND2_X1 U163 ( .A1(n99), .A2(n62), .ZN(n9) );
  INV_X1 U164 ( .A(n61), .ZN(n99) );
  NAND2_X1 U165 ( .A1(n180), .A2(n53), .ZN(n7) );
  NAND2_X1 U166 ( .A1(n182), .A2(n79), .ZN(n13) );
  NAND2_X1 U167 ( .A1(n179), .A2(n71), .ZN(n11) );
  NAND2_X1 U168 ( .A1(n104), .A2(n82), .ZN(n14) );
  INV_X1 U169 ( .A(n81), .ZN(n104) );
  NAND2_X1 U170 ( .A1(n98), .A2(n59), .ZN(n8) );
  NAND2_X1 U171 ( .A1(n181), .A2(n87), .ZN(n15) );
  NAND2_X1 U172 ( .A1(n102), .A2(n74), .ZN(n12) );
  INV_X1 U173 ( .A(n73), .ZN(n102) );
  NAND2_X1 U174 ( .A1(n100), .A2(n66), .ZN(n10) );
  INV_X1 U175 ( .A(n65), .ZN(n100) );
  XNOR2_X1 U176 ( .A(n11), .B(n72), .ZN(SUM[5]) );
  XNOR2_X1 U177 ( .A(n13), .B(n80), .ZN(SUM[3]) );
  XOR2_X1 U178 ( .A(n14), .B(n83), .Z(SUM[2]) );
  NAND2_X1 U179 ( .A1(n168), .A2(n28), .ZN(n3) );
  NAND2_X1 U180 ( .A1(n185), .A2(n37), .ZN(n4) );
  AOI21_X1 U181 ( .B1(n42), .B2(n34), .A(n35), .ZN(n33) );
  NOR2_X1 U182 ( .A1(A[11]), .A2(B[11]), .ZN(n39) );
  OR2_X1 U183 ( .A1(A[5]), .A2(B[5]), .ZN(n179) );
  NOR2_X1 U184 ( .A1(A[7]), .A2(B[7]), .ZN(n61) );
  OR2_X1 U185 ( .A1(B[9]), .A2(A[9]), .ZN(n180) );
  NOR2_X1 U186 ( .A1(A[2]), .A2(B[2]), .ZN(n81) );
  XOR2_X1 U187 ( .A(n49), .B(n6), .Z(SUM[10]) );
  NAND2_X1 U188 ( .A1(A[11]), .A2(B[11]), .ZN(n40) );
  OR2_X1 U189 ( .A1(A[1]), .A2(B[1]), .ZN(n181) );
  OR2_X1 U190 ( .A1(A[3]), .A2(B[3]), .ZN(n182) );
  OR2_X1 U191 ( .A1(A[10]), .A2(B[10]), .ZN(n183) );
  NAND2_X1 U192 ( .A1(n166), .A2(n18), .ZN(n1) );
  NOR2_X1 U193 ( .A1(A[4]), .A2(B[4]), .ZN(n73) );
  XNOR2_X1 U194 ( .A(n60), .B(n8), .ZN(SUM[8]) );
  XNOR2_X1 U195 ( .A(n54), .B(n7), .ZN(SUM[9]) );
  NOR2_X1 U196 ( .A1(A[6]), .A2(B[6]), .ZN(n65) );
  NAND2_X1 U197 ( .A1(A[7]), .A2(B[7]), .ZN(n62) );
  NAND2_X1 U198 ( .A1(A[2]), .A2(B[2]), .ZN(n82) );
  NAND2_X1 U199 ( .A1(A[1]), .A2(B[1]), .ZN(n87) );
  NAND2_X1 U200 ( .A1(A[0]), .A2(B[0]), .ZN(n90) );
  NAND2_X1 U201 ( .A1(A[4]), .A2(B[4]), .ZN(n74) );
  NAND2_X1 U202 ( .A1(A[6]), .A2(B[6]), .ZN(n66) );
  NAND2_X1 U203 ( .A1(A[8]), .A2(B[8]), .ZN(n59) );
  XOR2_X1 U204 ( .A(n63), .B(n9), .Z(SUM[7]) );
  XNOR2_X1 U205 ( .A(n15), .B(n88), .ZN(SUM[1]) );
  NAND2_X1 U206 ( .A1(A[5]), .A2(B[5]), .ZN(n71) );
  NAND2_X1 U207 ( .A1(A[12]), .A2(B[12]), .ZN(n37) );
  OR2_X1 U208 ( .A1(A[12]), .A2(B[12]), .ZN(n185) );
  AND2_X1 U209 ( .A1(A[14]), .A2(B[14]), .ZN(n186) );
  NAND2_X1 U210 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  NOR2_X1 U211 ( .A1(A[13]), .A2(B[13]), .ZN(n27) );
  NAND2_X1 U212 ( .A1(n183), .A2(n48), .ZN(n6) );
  NAND2_X1 U213 ( .A1(A[9]), .A2(B[9]), .ZN(n53) );
  OAI21_X1 U214 ( .B1(n41), .B2(n39), .A(n40), .ZN(n38) );
  AOI21_X1 U215 ( .B1(n184), .B2(n172), .A(n186), .ZN(n21) );
  NAND2_X1 U216 ( .A1(n168), .A2(n184), .ZN(n20) );
  NAND2_X1 U217 ( .A1(n184), .A2(n25), .ZN(n2) );
  INV_X1 U218 ( .A(n163), .ZN(n98) );
  NOR2_X1 U219 ( .A1(n58), .A2(n61), .ZN(n56) );
  OAI21_X1 U220 ( .B1(n58), .B2(n62), .A(n59), .ZN(n57) );
  XOR2_X1 U221 ( .A(n10), .B(n67), .Z(SUM[6]) );
  XOR2_X1 U222 ( .A(n12), .B(n75), .Z(SUM[4]) );
  OAI21_X1 U223 ( .B1(n67), .B2(n65), .A(n66), .ZN(n64) );
  NAND2_X1 U224 ( .A1(A[3]), .A2(B[3]), .ZN(n79) );
  NOR2_X1 U225 ( .A1(n176), .A2(n39), .ZN(n34) );
  OAI21_X1 U226 ( .B1(n40), .B2(n36), .A(n37), .ZN(n35) );
  NOR2_X1 U227 ( .A1(A[12]), .A2(B[12]), .ZN(n36) );
  NAND2_X1 U228 ( .A1(A[15]), .A2(B[15]), .ZN(n18) );
  INV_X1 U229 ( .A(n48), .ZN(n46) );
  NAND2_X1 U230 ( .A1(n183), .A2(n180), .ZN(n43) );
  AOI21_X1 U231 ( .B1(n183), .B2(n51), .A(n46), .ZN(n44) );
  XNOR2_X1 U232 ( .A(n38), .B(n4), .ZN(SUM[12]) );
  XNOR2_X1 U233 ( .A(n26), .B(n2), .ZN(SUM[14]) );
  XNOR2_X1 U234 ( .A(n19), .B(n1), .ZN(SUM[15]) );
  NAND2_X1 U235 ( .A1(A[14]), .A2(B[14]), .ZN(n25) );
  XOR2_X1 U236 ( .A(n33), .B(n3), .Z(SUM[13]) );
  OAI21_X1 U237 ( .B1(n177), .B2(n27), .A(n28), .ZN(n26) );
  NAND2_X1 U238 ( .A1(A[10]), .A2(B[10]), .ZN(n48) );
  OAI21_X1 U239 ( .B1(n177), .B2(n20), .A(n21), .ZN(n19) );
  OAI21_X1 U240 ( .B1(n43), .B2(n55), .A(n44), .ZN(n42) );
endmodule


module layer1_8_4_8_16_datapath_M8_N4_T16_P8_0 ( clk, clear_acc, data_out_x, 
        data_out, data_out_w, data_out_b, wr_en_y, m_valid, m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [3:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N27, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, n30, n31, n86, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n105,
         n106, n107, n108, n109, n110, n111, n112, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n12), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n103), .CK(clk), .Q(n16) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n102), .CK(clk), .Q(n17) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n101), .CK(clk), .Q(n18) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n100), .CK(clk), .Q(n19) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n96), .CK(clk), .Q(n23) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n95), .CK(clk), .Q(n24) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n94), .CK(clk), .Q(n25) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n93), .CK(clk), .Q(n26) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n92), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n91), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n90), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n89), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n88), .CK(clk), .Q(n33) );
  layer1_8_4_8_16_datapath_M8_N4_T16_P8_0_DW_mult_tc_1 mult_183 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer1_8_4_8_16_datapath_M8_N4_T16_P8_0_DW01_add_2 add_184 ( .A({n129, n130, 
        n131, n132, n133, n134, n120, n121, n122, n123, n124, n125, n126, n127, 
        n128, n135}), .B({f[15], n38, n39, n41, n43, n45, f[9:0]}), .CI(1'b0), 
        .SUM(adder) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n98), .CK(clk), .Q(n21) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n97), .CK(clk), .Q(n22) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n99), .CK(clk), .Q(n20) );
  DFF_X1 \data_out_reg[15]  ( .D(n167), .CK(clk), .Q(data_out[15]), .QN(n136)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n166), .CK(clk), .Q(data_out[14]), .QN(n137)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n165), .CK(clk), .Q(data_out[13]), .QN(n138)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n164), .CK(clk), .Q(data_out[12]), .QN(n139)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n163), .CK(clk), .Q(data_out[11]), .QN(n140)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n162), .CK(clk), .Q(data_out[10]), .QN(n141)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n161), .CK(clk), .Q(data_out[9]), .QN(n142) );
  DFF_X1 \data_out_reg[8]  ( .D(n160), .CK(clk), .Q(data_out[8]), .QN(n143) );
  DFF_X1 \data_out_reg[7]  ( .D(n159), .CK(clk), .Q(data_out[7]), .QN(n144) );
  DFF_X1 \data_out_reg[6]  ( .D(n158), .CK(clk), .Q(data_out[6]), .QN(n145) );
  DFF_X1 \data_out_reg[5]  ( .D(n157), .CK(clk), .Q(data_out[5]), .QN(n146) );
  DFF_X1 \data_out_reg[4]  ( .D(n156), .CK(clk), .Q(data_out[4]), .QN(n147) );
  DFF_X1 \data_out_reg[3]  ( .D(n155), .CK(clk), .Q(data_out[3]), .QN(n148) );
  DFF_X1 \data_out_reg[2]  ( .D(n154), .CK(clk), .Q(data_out[2]), .QN(n149) );
  DFF_X1 \data_out_reg[1]  ( .D(n153), .CK(clk), .Q(data_out[1]), .QN(n150) );
  DFF_X1 \data_out_reg[0]  ( .D(n152), .CK(clk), .Q(data_out[0]), .QN(n151) );
  DFF_X1 \f_reg[8]  ( .D(n73), .CK(clk), .Q(f[8]), .QN(n111) );
  DFF_X1 \f_reg[7]  ( .D(n74), .CK(clk), .Q(f[7]), .QN(n112) );
  DFF_X1 \f_reg[6]  ( .D(n75), .CK(clk), .Q(f[6]), .QN(n61) );
  DFF_X1 \f_reg[1]  ( .D(n80), .CK(clk), .Q(f[1]), .QN(n118) );
  DFF_X1 \f_reg[5]  ( .D(n76), .CK(clk), .Q(f[5]), .QN(n60) );
  DFF_X1 \f_reg[4]  ( .D(n77), .CK(clk), .Q(f[4]), .QN(n59) );
  DFF_X1 \f_reg[3]  ( .D(n78), .CK(clk), .Q(f[3]), .QN(n58) );
  DFF_X1 \f_reg[2]  ( .D(n79), .CK(clk), .Q(f[2]), .QN(n117) );
  DFF_X1 \f_reg[0]  ( .D(n81), .CK(clk), .Q(f[0]), .QN(n119) );
  DFF_X1 \f_reg[9]  ( .D(n72), .CK(clk), .Q(f[9]), .QN(n110) );
  DFF_X1 \f_reg[10]  ( .D(n71), .CK(clk), .Q(n45), .QN(n109) );
  DFF_X1 \f_reg[11]  ( .D(n70), .CK(clk), .Q(n43), .QN(n108) );
  DFF_X1 \f_reg[13]  ( .D(n68), .CK(clk), .Q(n39), .QN(n106) );
  DFF_X1 \f_reg[12]  ( .D(n69), .CK(clk), .Q(n41), .QN(n107) );
  DFF_X1 \f_reg[14]  ( .D(n2), .CK(clk), .Q(n38), .QN(n105) );
  DFF_X1 \f_reg[15]  ( .D(n4), .CK(clk), .Q(f[15]), .QN(n66) );
  DFF_X2 delay_reg ( .D(N27), .CK(clk), .Q(n35), .QN(n86) );
  AND2_X1 U3 ( .A1(clear_acc_delay), .A2(n86), .ZN(n1) );
  MUX2_X2 U4 ( .A(n16), .B(N44), .S(n86), .Z(n129) );
  MUX2_X2 U5 ( .A(n23), .B(N37), .S(n86), .Z(n121) );
  NAND3_X1 U6 ( .A1(n9), .A2(n8), .A3(n10), .ZN(n2) );
  MUX2_X1 U8 ( .A(N40), .B(n20), .S(n35), .Z(n133) );
  MUX2_X2 U9 ( .A(N43), .B(n17), .S(n35), .Z(n130) );
  NAND3_X1 U10 ( .A1(n6), .A2(n5), .A3(n7), .ZN(n4) );
  MUX2_X2 U11 ( .A(n18), .B(N42), .S(n86), .Z(n131) );
  NAND2_X1 U12 ( .A1(data_out_b[15]), .A2(n12), .ZN(n5) );
  NAND2_X1 U13 ( .A1(adder[15]), .A2(n11), .ZN(n6) );
  NAND2_X1 U14 ( .A1(n56), .A2(f[15]), .ZN(n7) );
  NAND2_X1 U15 ( .A1(data_out_b[14]), .A2(n12), .ZN(n8) );
  NAND2_X1 U16 ( .A1(adder[14]), .A2(n11), .ZN(n9) );
  NAND2_X1 U17 ( .A1(n56), .A2(n38), .ZN(n10) );
  AND2_X2 U18 ( .A1(n37), .A2(n13), .ZN(n11) );
  MUX2_X2 U19 ( .A(n19), .B(N41), .S(n86), .Z(n132) );
  INV_X1 U20 ( .A(n37), .ZN(n56) );
  INV_X1 U21 ( .A(clear_acc), .ZN(n13) );
  NAND2_X1 U22 ( .A1(n82), .A2(N27), .ZN(n30) );
  INV_X1 U23 ( .A(wr_en_y), .ZN(n82) );
  OAI22_X1 U24 ( .A1(n148), .A2(n30), .B1(n58), .B2(n31), .ZN(n155) );
  OAI22_X1 U25 ( .A1(n147), .A2(n30), .B1(n59), .B2(n31), .ZN(n156) );
  OAI22_X1 U26 ( .A1(n146), .A2(n30), .B1(n60), .B2(n31), .ZN(n157) );
  OAI22_X1 U27 ( .A1(n145), .A2(n30), .B1(n61), .B2(n31), .ZN(n158) );
  OAI22_X1 U28 ( .A1(n144), .A2(n30), .B1(n112), .B2(n31), .ZN(n159) );
  OAI22_X1 U29 ( .A1(n143), .A2(n30), .B1(n111), .B2(n31), .ZN(n160) );
  OAI22_X1 U30 ( .A1(n142), .A2(n30), .B1(n110), .B2(n31), .ZN(n161) );
  MUX2_X1 U31 ( .A(n26), .B(N34), .S(n86), .Z(n124) );
  INV_X1 U32 ( .A(n13), .ZN(n12) );
  AND3_X1 U33 ( .A1(sel[1]), .A2(sel[2]), .A3(sel[0]), .ZN(n15) );
  INV_X1 U34 ( .A(m_ready), .ZN(n14) );
  NAND2_X1 U35 ( .A1(m_valid), .A2(n14), .ZN(n34) );
  OAI21_X1 U36 ( .B1(sel[3]), .B2(n15), .A(n34), .ZN(N27) );
  MUX2_X1 U37 ( .A(n16), .B(N44), .S(n1), .Z(n103) );
  MUX2_X1 U38 ( .A(n17), .B(N43), .S(n1), .Z(n102) );
  MUX2_X1 U39 ( .A(n18), .B(N42), .S(n1), .Z(n101) );
  MUX2_X1 U40 ( .A(n19), .B(N41), .S(n1), .Z(n100) );
  MUX2_X1 U41 ( .A(n20), .B(N40), .S(n1), .Z(n99) );
  MUX2_X1 U42 ( .A(n21), .B(N39), .S(n1), .Z(n98) );
  MUX2_X1 U43 ( .A(n21), .B(N39), .S(n86), .Z(n134) );
  MUX2_X1 U44 ( .A(n22), .B(N38), .S(n1), .Z(n97) );
  MUX2_X1 U45 ( .A(n22), .B(N38), .S(n86), .Z(n120) );
  MUX2_X1 U46 ( .A(n23), .B(N37), .S(n1), .Z(n96) );
  MUX2_X1 U47 ( .A(n24), .B(N36), .S(n1), .Z(n95) );
  MUX2_X1 U48 ( .A(n24), .B(N36), .S(n86), .Z(n122) );
  MUX2_X1 U49 ( .A(n25), .B(N35), .S(n1), .Z(n94) );
  MUX2_X1 U50 ( .A(n25), .B(N35), .S(n86), .Z(n123) );
  MUX2_X1 U51 ( .A(n26), .B(N34), .S(n1), .Z(n93) );
  MUX2_X1 U52 ( .A(n27), .B(N33), .S(n1), .Z(n92) );
  MUX2_X1 U53 ( .A(n27), .B(N33), .S(n86), .Z(n125) );
  MUX2_X1 U54 ( .A(n28), .B(N32), .S(n1), .Z(n91) );
  MUX2_X1 U55 ( .A(n28), .B(N32), .S(n86), .Z(n126) );
  MUX2_X1 U56 ( .A(n29), .B(N31), .S(n1), .Z(n90) );
  MUX2_X1 U57 ( .A(n29), .B(N31), .S(n86), .Z(n127) );
  MUX2_X1 U58 ( .A(n32), .B(N30), .S(n1), .Z(n89) );
  MUX2_X1 U59 ( .A(n32), .B(N30), .S(n86), .Z(n128) );
  MUX2_X1 U60 ( .A(n33), .B(N29), .S(n1), .Z(n88) );
  MUX2_X1 U61 ( .A(n33), .B(N29), .S(n86), .Z(n135) );
  INV_X1 U62 ( .A(n34), .ZN(n36) );
  OAI21_X1 U63 ( .B1(n36), .B2(n35), .A(n13), .ZN(n37) );
  AOI222_X1 U64 ( .A1(data_out_b[13]), .A2(n12), .B1(adder[13]), .B2(n11), 
        .C1(n56), .C2(n39), .ZN(n40) );
  INV_X1 U65 ( .A(n40), .ZN(n68) );
  AOI222_X1 U66 ( .A1(data_out_b[12]), .A2(n12), .B1(adder[12]), .B2(n11), 
        .C1(n56), .C2(n41), .ZN(n42) );
  INV_X1 U67 ( .A(n42), .ZN(n69) );
  AOI222_X1 U68 ( .A1(data_out_b[11]), .A2(n12), .B1(adder[11]), .B2(n11), 
        .C1(n56), .C2(n43), .ZN(n44) );
  INV_X1 U69 ( .A(n44), .ZN(n70) );
  AOI222_X1 U70 ( .A1(data_out_b[10]), .A2(n12), .B1(adder[10]), .B2(n11), 
        .C1(n56), .C2(n45), .ZN(n46) );
  INV_X1 U71 ( .A(n46), .ZN(n71) );
  AOI222_X1 U72 ( .A1(data_out_b[8]), .A2(n12), .B1(adder[8]), .B2(n11), .C1(
        n56), .C2(f[8]), .ZN(n47) );
  INV_X1 U73 ( .A(n47), .ZN(n73) );
  AOI222_X1 U74 ( .A1(data_out_b[7]), .A2(n12), .B1(adder[7]), .B2(n11), .C1(
        n56), .C2(f[7]), .ZN(n48) );
  INV_X1 U75 ( .A(n48), .ZN(n74) );
  AOI222_X1 U76 ( .A1(data_out_b[6]), .A2(n12), .B1(adder[6]), .B2(n11), .C1(
        n56), .C2(f[6]), .ZN(n49) );
  INV_X1 U77 ( .A(n49), .ZN(n75) );
  AOI222_X1 U78 ( .A1(data_out_b[5]), .A2(n12), .B1(adder[5]), .B2(n11), .C1(
        n56), .C2(f[5]), .ZN(n50) );
  INV_X1 U79 ( .A(n50), .ZN(n76) );
  AOI222_X1 U80 ( .A1(data_out_b[4]), .A2(n12), .B1(adder[4]), .B2(n11), .C1(
        n56), .C2(f[4]), .ZN(n51) );
  INV_X1 U81 ( .A(n51), .ZN(n77) );
  AOI222_X1 U82 ( .A1(data_out_b[3]), .A2(n12), .B1(adder[3]), .B2(n11), .C1(
        n56), .C2(f[3]), .ZN(n52) );
  INV_X1 U83 ( .A(n52), .ZN(n78) );
  AOI222_X1 U84 ( .A1(data_out_b[2]), .A2(n12), .B1(adder[2]), .B2(n11), .C1(
        n56), .C2(f[2]), .ZN(n53) );
  INV_X1 U85 ( .A(n53), .ZN(n79) );
  AOI222_X1 U86 ( .A1(data_out_b[1]), .A2(n12), .B1(adder[1]), .B2(n11), .C1(
        n56), .C2(f[1]), .ZN(n54) );
  INV_X1 U87 ( .A(n54), .ZN(n80) );
  AOI222_X1 U88 ( .A1(data_out_b[0]), .A2(n12), .B1(adder[0]), .B2(n11), .C1(
        n56), .C2(f[0]), .ZN(n55) );
  INV_X1 U89 ( .A(n55), .ZN(n81) );
  AOI222_X1 U90 ( .A1(data_out_b[9]), .A2(n12), .B1(adder[9]), .B2(n11), .C1(
        n56), .C2(f[9]), .ZN(n57) );
  INV_X1 U91 ( .A(n57), .ZN(n72) );
  NOR4_X1 U92 ( .A1(n43), .A2(n41), .A3(n39), .A4(n38), .ZN(n65) );
  NOR4_X1 U93 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n45), .ZN(n64) );
  NAND4_X1 U94 ( .A1(n61), .A2(n60), .A3(n59), .A4(n58), .ZN(n62) );
  NOR4_X1 U95 ( .A1(n62), .A2(f[0]), .A3(f[1]), .A4(f[2]), .ZN(n63) );
  NAND3_X1 U96 ( .A1(n65), .A2(n64), .A3(n63), .ZN(n67) );
  NAND3_X1 U97 ( .A1(wr_en_y), .A2(n67), .A3(n66), .ZN(n31) );
  OAI22_X1 U98 ( .A1(n151), .A2(n30), .B1(n119), .B2(n31), .ZN(n152) );
  OAI22_X1 U99 ( .A1(n150), .A2(n30), .B1(n118), .B2(n31), .ZN(n153) );
  OAI22_X1 U100 ( .A1(n149), .A2(n30), .B1(n117), .B2(n31), .ZN(n154) );
  OAI22_X1 U101 ( .A1(n141), .A2(n30), .B1(n109), .B2(n31), .ZN(n162) );
  OAI22_X1 U102 ( .A1(n140), .A2(n30), .B1(n108), .B2(n31), .ZN(n163) );
  OAI22_X1 U103 ( .A1(n139), .A2(n30), .B1(n107), .B2(n31), .ZN(n164) );
  OAI22_X1 U104 ( .A1(n138), .A2(n30), .B1(n106), .B2(n31), .ZN(n165) );
  OAI22_X1 U105 ( .A1(n137), .A2(n30), .B1(n105), .B2(n31), .ZN(n166) );
  OAI22_X1 U106 ( .A1(n136), .A2(n30), .B1(n66), .B2(n31), .ZN(n167) );
endmodule


module layer1_8_4_8_16_datapath_M8_N4_T16_P8_7_DW_mult_tc_1 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n12, n13, n16, n18, n19, n21, n23, n25, n27, n29, n31,
         n34, n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n50, n52,
         n53, n55, n56, n57, n58, n59, n62, n63, n64, n65, n67, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n95, n96, n97, n98, n99, n101, n103,
         n104, n105, n106, n107, n111, n112, n113, n114, n115, n117, n119,
         n120, n122, n125, n129, n131, n139, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n237, n243, n249, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n418, n419,
         n420, n421, n422, n423, n424, n426, n427, n428, n429, n433, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U148 ( .A(n265), .B(n144), .Z(n145) );
  XOR2_X1 U150 ( .A(n271), .B(n146), .Z(n147) );
  XOR2_X1 U152 ( .A(n148), .B(n301), .Z(n149) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U161 ( .A(n177), .B(n168), .CI(n166), .CO(n163), .S(n164) );
  FA_X1 U162 ( .A(n170), .B(n172), .CI(n179), .CO(n165), .S(n166) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n263), .CI(n291), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n317), .B(n252), .CO(n173), .S(n174) );
  FA_X1 U167 ( .A(n180), .B(n187), .CI(n178), .CO(n175), .S(n176) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U169 ( .A(n193), .B(n282), .CI(n191), .CO(n179), .S(n180) );
  FA_X1 U170 ( .A(n268), .B(n292), .CI(n274), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U172 ( .A(n197), .B(n190), .CI(n188), .CO(n185), .S(n186) );
  FA_X1 U173 ( .A(n199), .B(n201), .CI(n192), .CO(n187), .S(n188) );
  FA_X1 U174 ( .A(n275), .B(n293), .CI(n194), .CO(n189), .S(n190) );
  FA_X1 U175 ( .A(n283), .B(n253), .CI(n305), .CO(n191), .S(n192) );
  HA_X1 U176 ( .A(n319), .B(n269), .CO(n193), .S(n194) );
  FA_X1 U177 ( .A(n205), .B(n200), .CI(n198), .CO(n195), .S(n196) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U179 ( .A(n284), .B(n294), .CI(n276), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n320), .B(n270), .CI(n306), .CO(n201), .S(n202) );
  FA_X1 U182 ( .A(n215), .B(n307), .CI(n210), .CO(n205), .S(n206) );
  FA_X1 U183 ( .A(n295), .B(n285), .CI(n254), .CO(n207), .S(n208) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U185 ( .A(n216), .B(n219), .CI(n214), .CO(n211), .S(n212) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n322), .B(n278), .CI(n308), .CO(n215), .S(n216) );
  FA_X1 U188 ( .A(n225), .B(n222), .CI(n220), .CO(n217), .S(n218) );
  FA_X1 U189 ( .A(n255), .B(n309), .CI(n297), .CO(n219), .S(n220) );
  HA_X1 U190 ( .A(n323), .B(n287), .CO(n221), .S(n222) );
  FA_X1 U192 ( .A(n324), .B(n288), .CI(n310), .CO(n225), .S(n226) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  HA_X1 U194 ( .A(n325), .B(n311), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n326), .B(n300), .CI(n312), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  CLKBUF_X1 U414 ( .A(n556), .Z(n542) );
  CLKBUF_X1 U415 ( .A(n556), .Z(n543) );
  CLKBUF_X1 U416 ( .A(n96), .Z(n531) );
  OR2_X1 U417 ( .A1(n196), .A2(n203), .ZN(n490) );
  XOR2_X1 U418 ( .A(n587), .B(a[12]), .Z(n37) );
  NAND2_X1 U419 ( .A1(n429), .A2(n27), .ZN(n29) );
  INV_X1 U420 ( .A(n501), .ZN(n111) );
  OR2_X1 U421 ( .A1(n186), .A2(n195), .ZN(n491) );
  OR2_X1 U422 ( .A1(n329), .A2(n258), .ZN(n492) );
  CLKBUF_X1 U423 ( .A(n86), .Z(n493) );
  INV_X2 U424 ( .A(n578), .ZN(n577) );
  BUF_X1 U425 ( .A(n497), .Z(n525) );
  INV_X1 U426 ( .A(n497), .ZN(n552) );
  XOR2_X1 U427 ( .A(n585), .B(a[10]), .Z(n497) );
  CLKBUF_X1 U428 ( .A(n570), .Z(n494) );
  INV_X1 U429 ( .A(n578), .ZN(n576) );
  INV_X1 U430 ( .A(n494), .ZN(n495) );
  CLKBUF_X1 U431 ( .A(n574), .Z(n496) );
  INV_X1 U432 ( .A(n577), .ZN(n498) );
  CLKBUF_X1 U433 ( .A(n18), .Z(n499) );
  INV_X1 U434 ( .A(n507), .ZN(n500) );
  AND2_X2 U435 ( .A1(n232), .A2(n233), .ZN(n501) );
  AND2_X1 U436 ( .A1(n529), .A2(n528), .ZN(n502) );
  AND2_X1 U437 ( .A1(n528), .A2(n529), .ZN(n45) );
  OR2_X1 U438 ( .A1(n522), .A2(n570), .ZN(n508) );
  CLKBUF_X1 U439 ( .A(n228), .Z(n503) );
  INV_X1 U440 ( .A(n95), .ZN(n504) );
  INV_X1 U441 ( .A(n535), .ZN(n95) );
  AND2_X1 U442 ( .A1(n212), .A2(n217), .ZN(n535) );
  OR2_X2 U443 ( .A1(n522), .A2(n507), .ZN(n12) );
  OAI21_X1 U444 ( .B1(n91), .B2(n89), .A(n90), .ZN(n505) );
  INV_X1 U445 ( .A(n544), .ZN(n506) );
  INV_X1 U446 ( .A(n544), .ZN(n27) );
  INV_X1 U447 ( .A(n570), .ZN(n521) );
  XNOR2_X1 U448 ( .A(n575), .B(a[2]), .ZN(n507) );
  XNOR2_X1 U449 ( .A(n226), .B(n509), .ZN(n224) );
  XNOR2_X1 U450 ( .A(n229), .B(n298), .ZN(n509) );
  NOR2_X1 U451 ( .A1(n164), .A2(n175), .ZN(n510) );
  NOR2_X1 U452 ( .A1(n164), .A2(n175), .ZN(n75) );
  XNOR2_X1 U453 ( .A(n587), .B(a[10]), .ZN(n428) );
  CLKBUF_X1 U454 ( .A(n104), .Z(n511) );
  INV_X1 U455 ( .A(n581), .ZN(n512) );
  INV_X1 U456 ( .A(n581), .ZN(n513) );
  INV_X1 U457 ( .A(n581), .ZN(n580) );
  INV_X1 U458 ( .A(n582), .ZN(n514) );
  INV_X1 U459 ( .A(n237), .ZN(n515) );
  INV_X1 U460 ( .A(n585), .ZN(n516) );
  INV_X1 U461 ( .A(n585), .ZN(n584) );
  NAND2_X1 U462 ( .A1(n428), .A2(n497), .ZN(n517) );
  XOR2_X1 U463 ( .A(n579), .B(a[6]), .Z(n518) );
  OR2_X1 U464 ( .A1(n176), .A2(n185), .ZN(n519) );
  BUF_X2 U465 ( .A(n21), .Z(n520) );
  XNOR2_X1 U466 ( .A(n575), .B(n249), .ZN(n433) );
  XOR2_X1 U467 ( .A(n578), .B(a[2]), .Z(n522) );
  OR2_X1 U468 ( .A1(n196), .A2(n203), .ZN(n523) );
  BUF_X2 U469 ( .A(n569), .Z(n524) );
  INV_X1 U470 ( .A(n249), .ZN(n569) );
  INV_X2 U471 ( .A(n587), .ZN(n586) );
  INV_X1 U472 ( .A(n490), .ZN(n526) );
  XNOR2_X1 U473 ( .A(n579), .B(a[6]), .ZN(n21) );
  NOR2_X1 U474 ( .A1(n186), .A2(n195), .ZN(n527) );
  NOR2_X1 U475 ( .A1(n186), .A2(n195), .ZN(n82) );
  NAND2_X1 U476 ( .A1(n505), .A2(n80), .ZN(n528) );
  INV_X1 U477 ( .A(n81), .ZN(n529) );
  INV_X1 U478 ( .A(n575), .ZN(n530) );
  OR2_X1 U479 ( .A1(n503), .A2(n231), .ZN(n532) );
  OAI21_X1 U480 ( .B1(n99), .B2(n97), .A(n98), .ZN(n96) );
  OR2_X2 U481 ( .A1(n533), .A2(n518), .ZN(n23) );
  XOR2_X1 U482 ( .A(n583), .B(a[6]), .Z(n533) );
  INV_X1 U483 ( .A(n574), .ZN(n534) );
  INV_X1 U484 ( .A(n513), .ZN(n536) );
  OAI21_X1 U485 ( .B1(n115), .B2(n113), .A(n114), .ZN(n537) );
  OR2_X1 U486 ( .A1(n234), .A2(n257), .ZN(n538) );
  OAI21_X1 U487 ( .B1(n115), .B2(n113), .A(n114), .ZN(n112) );
  OR2_X2 U488 ( .A1(n539), .A2(n553), .ZN(n18) );
  XNOR2_X1 U489 ( .A(n580), .B(a[4]), .ZN(n539) );
  INV_X2 U490 ( .A(n553), .ZN(n16) );
  XNOR2_X1 U491 ( .A(n502), .B(n540), .ZN(product[12]) );
  AND2_X1 U492 ( .A1(n519), .A2(n79), .ZN(n540) );
  OAI21_X1 U493 ( .B1(n91), .B2(n89), .A(n90), .ZN(n88) );
  BUF_X1 U494 ( .A(n556), .Z(n541) );
  XNOR2_X1 U495 ( .A(n583), .B(a[8]), .ZN(n544) );
  INV_X2 U496 ( .A(n575), .ZN(n574) );
  XOR2_X1 U497 ( .A(n208), .B(n213), .Z(n545) );
  XOR2_X1 U498 ( .A(n206), .B(n545), .Z(n204) );
  NAND2_X1 U499 ( .A1(n206), .A2(n208), .ZN(n546) );
  NAND2_X1 U500 ( .A1(n206), .A2(n213), .ZN(n547) );
  NAND2_X1 U501 ( .A1(n208), .A2(n213), .ZN(n548) );
  NAND3_X1 U502 ( .A1(n546), .A2(n547), .A3(n548), .ZN(n203) );
  NAND2_X1 U503 ( .A1(n226), .A2(n229), .ZN(n549) );
  NAND2_X1 U504 ( .A1(n226), .A2(n298), .ZN(n550) );
  NAND2_X1 U505 ( .A1(n229), .A2(n298), .ZN(n551) );
  NAND3_X1 U506 ( .A1(n549), .A2(n550), .A3(n551), .ZN(n223) );
  XNOR2_X1 U507 ( .A(n578), .B(a[4]), .ZN(n553) );
  INV_X1 U508 ( .A(n97), .ZN(n131) );
  NOR2_X1 U509 ( .A1(n203), .A2(n196), .ZN(n85) );
  INV_X1 U510 ( .A(n581), .ZN(n579) );
  AOI21_X1 U511 ( .B1(n531), .B2(n558), .A(n504), .ZN(n554) );
  CLKBUF_X1 U512 ( .A(n99), .Z(n555) );
  NAND2_X1 U513 ( .A1(n433), .A2(n569), .ZN(n556) );
  NAND2_X1 U514 ( .A1(n433), .A2(n569), .ZN(n6) );
  XNOR2_X1 U515 ( .A(n557), .B(n87), .ZN(product[10]) );
  AND2_X1 U516 ( .A1(n523), .A2(n86), .ZN(n557) );
  OR2_X1 U517 ( .A1(n152), .A2(n163), .ZN(n560) );
  OR2_X1 U518 ( .A1(n212), .A2(n217), .ZN(n558) );
  XOR2_X1 U519 ( .A(n555), .B(n559), .Z(product[7]) );
  NAND2_X1 U520 ( .A1(n131), .A2(n98), .ZN(n559) );
  INV_X2 U521 ( .A(n583), .ZN(n582) );
  OR2_X1 U522 ( .A1(n233), .A2(n232), .ZN(n563) );
  OR2_X1 U523 ( .A1(n328), .A2(n314), .ZN(n561) );
  NAND2_X1 U524 ( .A1(n560), .A2(n69), .ZN(n47) );
  INV_X1 U525 ( .A(n73), .ZN(n71) );
  AOI21_X1 U526 ( .B1(n74), .B2(n560), .A(n67), .ZN(n65) );
  INV_X1 U527 ( .A(n69), .ZN(n67) );
  NAND2_X1 U528 ( .A1(n73), .A2(n560), .ZN(n64) );
  INV_X1 U529 ( .A(n74), .ZN(n72) );
  NAND2_X1 U530 ( .A1(n129), .A2(n90), .ZN(n52) );
  INV_X1 U531 ( .A(n89), .ZN(n129) );
  NAND2_X1 U532 ( .A1(n125), .A2(n76), .ZN(n48) );
  INV_X1 U533 ( .A(n75), .ZN(n125) );
  OAI21_X1 U534 ( .B1(n510), .B2(n79), .A(n76), .ZN(n74) );
  NAND2_X1 U535 ( .A1(n491), .A2(n83), .ZN(n50) );
  NOR2_X1 U536 ( .A1(n75), .A2(n78), .ZN(n73) );
  XNOR2_X1 U537 ( .A(n531), .B(n53), .ZN(product[8]) );
  NAND2_X1 U538 ( .A1(n558), .A2(n95), .ZN(n53) );
  NAND2_X1 U539 ( .A1(n152), .A2(n163), .ZN(n69) );
  NAND2_X1 U540 ( .A1(n532), .A2(n106), .ZN(n56) );
  NOR2_X1 U541 ( .A1(n176), .A2(n185), .ZN(n78) );
  NAND2_X1 U542 ( .A1(n563), .A2(n111), .ZN(n57) );
  AOI21_X1 U543 ( .B1(n561), .B2(n120), .A(n117), .ZN(n115) );
  INV_X1 U544 ( .A(n119), .ZN(n117) );
  INV_X1 U545 ( .A(n122), .ZN(n120) );
  NAND2_X1 U546 ( .A1(n176), .A2(n185), .ZN(n79) );
  NAND2_X1 U547 ( .A1(n164), .A2(n175), .ZN(n76) );
  NAND2_X1 U548 ( .A1(n204), .A2(n211), .ZN(n90) );
  NAND2_X1 U549 ( .A1(n196), .A2(n203), .ZN(n86) );
  NAND2_X1 U550 ( .A1(n538), .A2(n114), .ZN(n58) );
  XNOR2_X1 U551 ( .A(n59), .B(n120), .ZN(product[2]) );
  NAND2_X1 U552 ( .A1(n561), .A2(n119), .ZN(n59) );
  XNOR2_X1 U553 ( .A(n63), .B(n46), .ZN(product[15]) );
  NAND2_X1 U554 ( .A1(n562), .A2(n62), .ZN(n46) );
  NAND2_X1 U555 ( .A1(n328), .A2(n314), .ZN(n119) );
  NOR2_X1 U556 ( .A1(n218), .A2(n223), .ZN(n97) );
  OR2_X1 U557 ( .A1(n139), .A2(n151), .ZN(n562) );
  NOR2_X1 U558 ( .A1(n234), .A2(n257), .ZN(n113) );
  NAND2_X1 U559 ( .A1(n218), .A2(n223), .ZN(n98) );
  NAND2_X1 U560 ( .A1(n228), .A2(n231), .ZN(n106) );
  OR2_X1 U561 ( .A1(n224), .A2(n227), .ZN(n564) );
  AND2_X1 U562 ( .A1(n492), .A2(n122), .ZN(product[1]) );
  OR2_X1 U563 ( .A1(n572), .A2(n498), .ZN(n392) );
  OR2_X1 U564 ( .A1(n572), .A2(n534), .ZN(n409) );
  XNOR2_X1 U565 ( .A(n574), .B(n572), .ZN(n408) );
  XNOR2_X1 U566 ( .A(n516), .B(n572), .ZN(n352) );
  XNOR2_X1 U567 ( .A(n155), .B(n566), .ZN(n139) );
  XNOR2_X1 U568 ( .A(n153), .B(n141), .ZN(n566) );
  XNOR2_X1 U569 ( .A(n157), .B(n567), .ZN(n141) );
  XNOR2_X1 U570 ( .A(n145), .B(n143), .ZN(n567) );
  OAI22_X1 U571 ( .A1(n42), .A2(n591), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U572 ( .A1(n572), .A2(n591), .ZN(n332) );
  OAI22_X1 U573 ( .A1(n517), .A2(n343), .B1(n342), .B2(n497), .ZN(n269) );
  XNOR2_X1 U574 ( .A(n586), .B(n572), .ZN(n343) );
  XNOR2_X1 U575 ( .A(n159), .B(n568), .ZN(n142) );
  XNOR2_X1 U576 ( .A(n315), .B(n261), .ZN(n568) );
  XNOR2_X1 U577 ( .A(n580), .B(n572), .ZN(n376) );
  AND2_X1 U578 ( .A1(n573), .A2(n553), .ZN(n300) );
  INV_X1 U579 ( .A(n37), .ZN(n237) );
  XNOR2_X1 U580 ( .A(n588), .B(n572), .ZN(n336) );
  AND2_X1 U581 ( .A1(n573), .A2(n494), .ZN(n314) );
  OAI22_X1 U582 ( .A1(n517), .A2(n342), .B1(n341), .B2(n525), .ZN(n268) );
  OAI22_X1 U583 ( .A1(n34), .A2(n341), .B1(n340), .B2(n525), .ZN(n267) );
  OAI22_X1 U584 ( .A1(n39), .A2(n336), .B1(n515), .B2(n335), .ZN(n263) );
  INV_X1 U585 ( .A(n19), .ZN(n583) );
  INV_X1 U586 ( .A(n25), .ZN(n585) );
  AND2_X1 U587 ( .A1(n573), .A2(n237), .ZN(n264) );
  AND2_X1 U588 ( .A1(n573), .A2(n243), .ZN(n288) );
  AND2_X1 U589 ( .A1(n573), .A2(n552), .ZN(n270) );
  AND2_X1 U590 ( .A1(n573), .A2(n235), .ZN(n260) );
  OAI22_X1 U591 ( .A1(n39), .A2(n335), .B1(n515), .B2(n334), .ZN(n262) );
  AND2_X1 U592 ( .A1(n573), .A2(n544), .ZN(n278) );
  OAI22_X1 U593 ( .A1(n34), .A2(n587), .B1(n344), .B2(n497), .ZN(n253) );
  INV_X1 U594 ( .A(n7), .ZN(n578) );
  INV_X1 U595 ( .A(n13), .ZN(n581) );
  OAI22_X1 U596 ( .A1(n34), .A2(n340), .B1(n339), .B2(n525), .ZN(n266) );
  INV_X1 U597 ( .A(n41), .ZN(n235) );
  XNOR2_X1 U598 ( .A(n582), .B(n572), .ZN(n363) );
  OAI22_X1 U599 ( .A1(n39), .A2(n589), .B1(n337), .B2(n515), .ZN(n252) );
  OR2_X1 U600 ( .A1(n572), .A2(n589), .ZN(n337) );
  OR2_X1 U601 ( .A1(n572), .A2(n587), .ZN(n344) );
  AND2_X1 U602 ( .A1(n573), .A2(n249), .ZN(product[0]) );
  OR2_X1 U603 ( .A1(n572), .A2(n536), .ZN(n377) );
  OR2_X1 U604 ( .A1(n572), .A2(n514), .ZN(n364) );
  OR2_X1 U605 ( .A1(n572), .A2(n585), .ZN(n353) );
  XNOR2_X1 U606 ( .A(n588), .B(a[14]), .ZN(n41) );
  OAI22_X1 U607 ( .A1(n39), .A2(n334), .B1(n515), .B2(n333), .ZN(n261) );
  XNOR2_X1 U608 ( .A(n588), .B(n422), .ZN(n333) );
  XNOR2_X1 U609 ( .A(n513), .B(b[11]), .ZN(n365) );
  XNOR2_X1 U610 ( .A(n582), .B(b[9]), .ZN(n354) );
  OAI22_X1 U611 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U612 ( .A(n590), .B(n424), .ZN(n330) );
  XNOR2_X1 U613 ( .A(n590), .B(n572), .ZN(n331) );
  XNOR2_X1 U614 ( .A(n586), .B(n423), .ZN(n341) );
  XNOR2_X1 U615 ( .A(n586), .B(n424), .ZN(n342) );
  XNOR2_X1 U616 ( .A(n586), .B(n422), .ZN(n340) );
  XNOR2_X1 U617 ( .A(n586), .B(n421), .ZN(n339) );
  XNOR2_X1 U618 ( .A(n588), .B(n424), .ZN(n335) );
  XNOR2_X1 U619 ( .A(n588), .B(n423), .ZN(n334) );
  XOR2_X1 U620 ( .A(n584), .B(a[8]), .Z(n429) );
  XNOR2_X1 U621 ( .A(n516), .B(n418), .ZN(n345) );
  OAI22_X1 U622 ( .A1(n517), .A2(n339), .B1(n338), .B2(n525), .ZN(n265) );
  XNOR2_X1 U623 ( .A(n586), .B(n420), .ZN(n338) );
  XNOR2_X1 U624 ( .A(n577), .B(b[13]), .ZN(n378) );
  XNOR2_X1 U625 ( .A(n574), .B(n424), .ZN(n407) );
  XNOR2_X1 U626 ( .A(n582), .B(n424), .ZN(n362) );
  XNOR2_X1 U627 ( .A(n584), .B(n424), .ZN(n351) );
  NAND2_X1 U628 ( .A1(n428), .A2(n497), .ZN(n34) );
  NAND2_X1 U629 ( .A1(n427), .A2(n37), .ZN(n39) );
  XNOR2_X1 U630 ( .A(n577), .B(n419), .ZN(n385) );
  XNOR2_X1 U631 ( .A(n574), .B(n423), .ZN(n406) );
  XNOR2_X1 U632 ( .A(n582), .B(n423), .ZN(n361) );
  XNOR2_X1 U633 ( .A(n582), .B(n422), .ZN(n360) );
  XNOR2_X1 U634 ( .A(n584), .B(n423), .ZN(n350) );
  XNOR2_X1 U635 ( .A(n516), .B(n422), .ZN(n349) );
  XNOR2_X1 U636 ( .A(n574), .B(n422), .ZN(n405) );
  XNOR2_X1 U637 ( .A(n582), .B(n420), .ZN(n358) );
  XNOR2_X1 U638 ( .A(n582), .B(n421), .ZN(n359) );
  XNOR2_X1 U639 ( .A(n516), .B(n421), .ZN(n348) );
  XNOR2_X1 U640 ( .A(n584), .B(n420), .ZN(n347) );
  XNOR2_X1 U641 ( .A(n530), .B(n421), .ZN(n404) );
  XNOR2_X1 U642 ( .A(n530), .B(n420), .ZN(n403) );
  XNOR2_X1 U643 ( .A(n582), .B(n419), .ZN(n357) );
  XNOR2_X1 U644 ( .A(n516), .B(n419), .ZN(n346) );
  XNOR2_X1 U645 ( .A(n574), .B(n419), .ZN(n402) );
  NAND2_X1 U646 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U647 ( .A(n590), .B(a[14]), .Z(n426) );
  BUF_X1 U648 ( .A(n43), .Z(n573) );
  XNOR2_X1 U649 ( .A(n576), .B(n418), .ZN(n384) );
  XNOR2_X1 U650 ( .A(n577), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U651 ( .A(n577), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U652 ( .A(n576), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U653 ( .A(n577), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U654 ( .A(n577), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U655 ( .A(n512), .B(n418), .ZN(n369) );
  XNOR2_X1 U656 ( .A(n513), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U657 ( .A(n512), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U658 ( .A(n580), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U659 ( .A(n574), .B(b[11]), .ZN(n397) );
  XNOR2_X1 U660 ( .A(n574), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U661 ( .A(n574), .B(b[13]), .ZN(n395) );
  XNOR2_X1 U662 ( .A(n496), .B(b[14]), .ZN(n394) );
  XNOR2_X1 U663 ( .A(n582), .B(n418), .ZN(n356) );
  XNOR2_X1 U664 ( .A(n582), .B(b[8]), .ZN(n355) );
  XNOR2_X1 U665 ( .A(n530), .B(n418), .ZN(n401) );
  XNOR2_X1 U666 ( .A(n530), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U667 ( .A(n530), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U668 ( .A(n574), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U669 ( .A(n496), .B(b[15]), .ZN(n393) );
  XOR2_X1 U670 ( .A(n588), .B(a[12]), .Z(n427) );
  XNOR2_X1 U671 ( .A(n575), .B(a[2]), .ZN(n570) );
  INV_X1 U672 ( .A(n1), .ZN(n575) );
  OAI22_X1 U673 ( .A1(n543), .A2(n395), .B1(n394), .B2(n524), .ZN(n316) );
  NAND2_X1 U674 ( .A1(n329), .A2(n258), .ZN(n122) );
  OAI22_X1 U675 ( .A1(n542), .A2(n394), .B1(n393), .B2(n524), .ZN(n315) );
  OAI22_X1 U676 ( .A1(n6), .A2(n399), .B1(n398), .B2(n569), .ZN(n320) );
  OAI22_X1 U677 ( .A1(n542), .A2(n401), .B1(n400), .B2(n524), .ZN(n322) );
  OAI22_X1 U678 ( .A1(n542), .A2(n396), .B1(n395), .B2(n524), .ZN(n317) );
  OAI22_X1 U679 ( .A1(n542), .A2(n397), .B1(n396), .B2(n524), .ZN(n318) );
  OAI22_X1 U680 ( .A1(n543), .A2(n400), .B1(n399), .B2(n524), .ZN(n321) );
  OAI22_X1 U681 ( .A1(n404), .A2(n6), .B1(n403), .B2(n524), .ZN(n325) );
  OAI22_X1 U682 ( .A1(n6), .A2(n406), .B1(n405), .B2(n524), .ZN(n327) );
  OAI22_X1 U683 ( .A1(n6), .A2(n405), .B1(n404), .B2(n524), .ZN(n326) );
  OAI22_X1 U684 ( .A1(n543), .A2(n398), .B1(n397), .B2(n524), .ZN(n319) );
  OAI22_X1 U685 ( .A1(n541), .A2(n402), .B1(n401), .B2(n524), .ZN(n323) );
  OAI22_X1 U686 ( .A1(n6), .A2(n403), .B1(n402), .B2(n524), .ZN(n324) );
  OAI22_X1 U687 ( .A1(n542), .A2(n407), .B1(n406), .B2(n524), .ZN(n328) );
  OAI22_X1 U688 ( .A1(n541), .A2(n408), .B1(n407), .B2(n524), .ZN(n329) );
  OAI22_X1 U689 ( .A1(n543), .A2(n534), .B1(n409), .B2(n524), .ZN(n258) );
  OAI21_X1 U690 ( .B1(n86), .B2(n527), .A(n83), .ZN(n81) );
  NOR2_X1 U691 ( .A1(n82), .A2(n85), .ZN(n80) );
  AOI21_X1 U692 ( .B1(n563), .B2(n537), .A(n501), .ZN(n571) );
  NAND2_X1 U693 ( .A1(n186), .A2(n195), .ZN(n83) );
  NAND2_X1 U694 ( .A1(n564), .A2(n103), .ZN(n55) );
  NAND2_X1 U695 ( .A1(n224), .A2(n227), .ZN(n103) );
  XNOR2_X1 U696 ( .A(n84), .B(n50), .ZN(product[11]) );
  XOR2_X1 U697 ( .A(n58), .B(n115), .Z(product[3]) );
  AOI21_X1 U698 ( .B1(n563), .B2(n112), .A(n501), .ZN(n107) );
  NOR2_X1 U699 ( .A1(n228), .A2(n231), .ZN(n105) );
  NOR2_X1 U700 ( .A1(n204), .A2(n211), .ZN(n89) );
  OAI22_X1 U701 ( .A1(n29), .A2(n346), .B1(n345), .B2(n506), .ZN(n271) );
  OAI22_X1 U702 ( .A1(n29), .A2(n350), .B1(n349), .B2(n506), .ZN(n275) );
  OAI22_X1 U703 ( .A1(n29), .A2(n347), .B1(n346), .B2(n506), .ZN(n272) );
  OAI22_X1 U704 ( .A1(n29), .A2(n348), .B1(n347), .B2(n506), .ZN(n273) );
  OAI22_X1 U705 ( .A1(n29), .A2(n349), .B1(n348), .B2(n506), .ZN(n274) );
  OAI22_X1 U706 ( .A1(n29), .A2(n585), .B1(n353), .B2(n506), .ZN(n254) );
  OAI22_X1 U707 ( .A1(n29), .A2(n351), .B1(n350), .B2(n506), .ZN(n276) );
  OAI22_X1 U708 ( .A1(n29), .A2(n352), .B1(n351), .B2(n506), .ZN(n277) );
  XNOR2_X1 U709 ( .A(n512), .B(n424), .ZN(n375) );
  XNOR2_X1 U710 ( .A(n580), .B(n419), .ZN(n370) );
  XNOR2_X1 U711 ( .A(n512), .B(n420), .ZN(n371) );
  XNOR2_X1 U712 ( .A(n580), .B(n423), .ZN(n374) );
  XNOR2_X1 U713 ( .A(n513), .B(n422), .ZN(n373) );
  XNOR2_X1 U714 ( .A(n513), .B(n421), .ZN(n372) );
  XNOR2_X1 U715 ( .A(n577), .B(n572), .ZN(n391) );
  XNOR2_X1 U716 ( .A(n577), .B(n420), .ZN(n386) );
  XNOR2_X1 U717 ( .A(n577), .B(n424), .ZN(n390) );
  XNOR2_X1 U718 ( .A(n576), .B(n423), .ZN(n389) );
  XNOR2_X1 U719 ( .A(n576), .B(n422), .ZN(n388) );
  XNOR2_X1 U720 ( .A(n577), .B(n421), .ZN(n387) );
  XNOR2_X1 U721 ( .A(n77), .B(n48), .ZN(product[13]) );
  OAI21_X1 U722 ( .B1(n87), .B2(n526), .A(n493), .ZN(n84) );
  INV_X1 U723 ( .A(n88), .ZN(n87) );
  OAI22_X1 U724 ( .A1(n23), .A2(n358), .B1(n357), .B2(n520), .ZN(n282) );
  OAI22_X1 U725 ( .A1(n23), .A2(n356), .B1(n355), .B2(n520), .ZN(n280) );
  OAI22_X1 U726 ( .A1(n23), .A2(n362), .B1(n361), .B2(n520), .ZN(n286) );
  OAI22_X1 U727 ( .A1(n23), .A2(n357), .B1(n356), .B2(n520), .ZN(n281) );
  OAI22_X1 U728 ( .A1(n23), .A2(n360), .B1(n359), .B2(n520), .ZN(n284) );
  OAI22_X1 U729 ( .A1(n23), .A2(n514), .B1(n364), .B2(n520), .ZN(n255) );
  OAI22_X1 U730 ( .A1(n23), .A2(n361), .B1(n360), .B2(n520), .ZN(n285) );
  OAI22_X1 U731 ( .A1(n23), .A2(n355), .B1(n354), .B2(n520), .ZN(n279) );
  OAI22_X1 U732 ( .A1(n23), .A2(n363), .B1(n362), .B2(n520), .ZN(n287) );
  OAI22_X1 U733 ( .A1(n23), .A2(n359), .B1(n358), .B2(n520), .ZN(n283) );
  INV_X1 U734 ( .A(n520), .ZN(n243) );
  AOI21_X1 U735 ( .B1(n96), .B2(n558), .A(n535), .ZN(n91) );
  OAI21_X1 U736 ( .B1(n105), .B2(n107), .A(n106), .ZN(n104) );
  INV_X1 U737 ( .A(n103), .ZN(n101) );
  NAND2_X1 U738 ( .A1(n151), .A2(n139), .ZN(n62) );
  OAI22_X1 U739 ( .A1(n499), .A2(n370), .B1(n369), .B2(n16), .ZN(n293) );
  OAI22_X1 U740 ( .A1(n499), .A2(n367), .B1(n366), .B2(n16), .ZN(n290) );
  OAI22_X1 U741 ( .A1(n18), .A2(n375), .B1(n374), .B2(n16), .ZN(n298) );
  OAI22_X1 U742 ( .A1(n18), .A2(n368), .B1(n367), .B2(n16), .ZN(n291) );
  OAI22_X1 U743 ( .A1(n18), .A2(n373), .B1(n372), .B2(n16), .ZN(n296) );
  OAI22_X1 U744 ( .A1(n18), .A2(n372), .B1(n371), .B2(n16), .ZN(n295) );
  OAI22_X1 U745 ( .A1(n18), .A2(n376), .B1(n375), .B2(n16), .ZN(n299) );
  OAI22_X1 U746 ( .A1(n18), .A2(n536), .B1(n377), .B2(n16), .ZN(n256) );
  OAI22_X1 U747 ( .A1(n18), .A2(n369), .B1(n368), .B2(n16), .ZN(n292) );
  OAI22_X1 U748 ( .A1(n18), .A2(n371), .B1(n370), .B2(n16), .ZN(n294) );
  OAI22_X1 U749 ( .A1(n18), .A2(n374), .B1(n373), .B2(n16), .ZN(n297) );
  OAI22_X1 U750 ( .A1(n18), .A2(n366), .B1(n365), .B2(n16), .ZN(n289) );
  XNOR2_X1 U751 ( .A(n511), .B(n55), .ZN(product[6]) );
  XNOR2_X1 U752 ( .A(n57), .B(n537), .ZN(product[4]) );
  AOI21_X1 U753 ( .B1(n104), .B2(n564), .A(n101), .ZN(n99) );
  XOR2_X1 U754 ( .A(n554), .B(n52), .Z(product[9]) );
  XOR2_X1 U755 ( .A(n56), .B(n571), .Z(product[5]) );
  OAI21_X1 U756 ( .B1(n45), .B2(n78), .A(n79), .ZN(n77) );
  OAI21_X1 U757 ( .B1(n45), .B2(n71), .A(n72), .ZN(n70) );
  OAI21_X1 U758 ( .B1(n64), .B2(n502), .A(n65), .ZN(n63) );
  XNOR2_X1 U759 ( .A(n70), .B(n47), .ZN(product[14]) );
  OAI22_X1 U760 ( .A1(n12), .A2(n379), .B1(n378), .B2(n495), .ZN(n301) );
  OAI22_X1 U761 ( .A1(n12), .A2(n380), .B1(n379), .B2(n500), .ZN(n302) );
  OAI22_X1 U762 ( .A1(n12), .A2(n385), .B1(n384), .B2(n500), .ZN(n307) );
  OAI22_X1 U763 ( .A1(n12), .A2(n382), .B1(n381), .B2(n500), .ZN(n304) );
  OAI22_X1 U764 ( .A1(n12), .A2(n381), .B1(n380), .B2(n521), .ZN(n303) );
  NAND2_X1 U765 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U766 ( .A1(n508), .A2(n383), .B1(n382), .B2(n500), .ZN(n305) );
  OAI22_X1 U767 ( .A1(n508), .A2(n384), .B1(n383), .B2(n521), .ZN(n306) );
  OAI22_X1 U768 ( .A1(n12), .A2(n386), .B1(n385), .B2(n495), .ZN(n308) );
  OAI22_X1 U769 ( .A1(n12), .A2(n387), .B1(n386), .B2(n521), .ZN(n309) );
  OAI22_X1 U770 ( .A1(n12), .A2(n498), .B1(n392), .B2(n495), .ZN(n257) );
  OAI22_X1 U771 ( .A1(n508), .A2(n389), .B1(n388), .B2(n500), .ZN(n311) );
  OAI22_X1 U772 ( .A1(n12), .A2(n388), .B1(n387), .B2(n521), .ZN(n310) );
  OAI22_X1 U773 ( .A1(n12), .A2(n390), .B1(n389), .B2(n521), .ZN(n312) );
  OAI22_X1 U774 ( .A1(n12), .A2(n391), .B1(n390), .B2(n500), .ZN(n313) );
  BUF_X4 U775 ( .A(n43), .Z(n572) );
  INV_X1 U776 ( .A(n31), .ZN(n587) );
  INV_X1 U777 ( .A(n589), .ZN(n588) );
  INV_X1 U778 ( .A(n36), .ZN(n589) );
  INV_X1 U779 ( .A(n591), .ZN(n590) );
  INV_X1 U780 ( .A(n40), .ZN(n591) );
  XOR2_X1 U781 ( .A(n259), .B(n251), .Z(n148) );
  XOR2_X1 U782 ( .A(n289), .B(n279), .Z(n146) );
  XOR2_X1 U783 ( .A(n149), .B(n147), .Z(n144) );
endmodule


module layer1_8_4_8_16_datapath_M8_N4_T16_P8_7_DW01_add_2 ( A, B, CI, SUM, CO
 );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n4, n6, n8, n9, n10, n11, n12, n13, n14, n15, n18, n19, n20,
         n21, n25, n26, n27, n28, n30, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n48, n49, n51, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n69, n71, n72, n73, n74, n75, n77,
         n79, n80, n81, n82, n83, n85, n87, n88, n90, n94, n95, n99, n100,
         n102, n104, n161, n162, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185;

  CLKBUF_X1 U126 ( .A(n182), .Z(n174) );
  XNOR2_X1 U127 ( .A(n169), .B(n161), .ZN(SUM[11]) );
  AND2_X1 U128 ( .A1(n95), .A2(n40), .ZN(n161) );
  OR2_X1 U129 ( .A1(A[8]), .A2(B[8]), .ZN(n162) );
  AND2_X1 U130 ( .A1(n178), .A2(n90), .ZN(SUM[0]) );
  OR2_X1 U131 ( .A1(A[15]), .A2(B[15]), .ZN(n164) );
  NOR2_X1 U132 ( .A1(A[8]), .A2(B[8]), .ZN(n165) );
  XNOR2_X1 U133 ( .A(n171), .B(n166), .ZN(SUM[9]) );
  AND2_X1 U134 ( .A1(n180), .A2(n53), .ZN(n166) );
  NOR2_X1 U135 ( .A1(A[8]), .A2(B[8]), .ZN(n58) );
  XNOR2_X1 U136 ( .A(n176), .B(n167), .ZN(SUM[13]) );
  AND2_X1 U137 ( .A1(n173), .A2(n28), .ZN(n167) );
  AOI21_X1 U138 ( .B1(n182), .B2(n51), .A(n175), .ZN(n168) );
  CLKBUF_X1 U139 ( .A(n41), .Z(n169) );
  OAI21_X1 U140 ( .B1(n55), .B2(n43), .A(n44), .ZN(n170) );
  INV_X1 U141 ( .A(n175), .ZN(n48) );
  AOI21_X1 U142 ( .B1(n56), .B2(n64), .A(n57), .ZN(n171) );
  NOR2_X1 U143 ( .A1(A[12]), .A2(B[12]), .ZN(n172) );
  NOR2_X1 U144 ( .A1(A[12]), .A2(B[12]), .ZN(n36) );
  OR2_X1 U145 ( .A1(A[13]), .A2(B[13]), .ZN(n173) );
  NOR2_X2 U146 ( .A1(A[11]), .A2(B[11]), .ZN(n39) );
  OR2_X2 U147 ( .A1(A[10]), .A2(B[10]), .ZN(n182) );
  AND2_X1 U148 ( .A1(A[10]), .A2(B[10]), .ZN(n175) );
  OR2_X2 U149 ( .A1(A[14]), .A2(B[14]), .ZN(n181) );
  AOI21_X1 U150 ( .B1(n42), .B2(n34), .A(n35), .ZN(n176) );
  AOI21_X1 U151 ( .B1(n42), .B2(n34), .A(n35), .ZN(n177) );
  NOR2_X1 U152 ( .A1(A[7]), .A2(B[7]), .ZN(n61) );
  OR2_X1 U153 ( .A1(A[9]), .A2(B[9]), .ZN(n180) );
  OR2_X1 U154 ( .A1(A[0]), .A2(B[0]), .ZN(n178) );
  INV_X1 U155 ( .A(n171), .ZN(n54) );
  INV_X1 U156 ( .A(n71), .ZN(n69) );
  OAI21_X1 U157 ( .B1(n83), .B2(n81), .A(n82), .ZN(n80) );
  AOI21_X1 U158 ( .B1(n179), .B2(n80), .A(n77), .ZN(n75) );
  INV_X1 U159 ( .A(n79), .ZN(n77) );
  AOI21_X1 U160 ( .B1(n54), .B2(n180), .A(n51), .ZN(n49) );
  NAND2_X1 U161 ( .A1(n162), .A2(n59), .ZN(n8) );
  INV_X1 U162 ( .A(n90), .ZN(n88) );
  OAI21_X1 U163 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  INV_X1 U164 ( .A(n53), .ZN(n51) );
  AOI21_X1 U165 ( .B1(n183), .B2(n88), .A(n85), .ZN(n83) );
  INV_X1 U166 ( .A(n87), .ZN(n85) );
  NAND2_X1 U167 ( .A1(n104), .A2(n82), .ZN(n14) );
  INV_X1 U168 ( .A(n81), .ZN(n104) );
  INV_X1 U169 ( .A(n39), .ZN(n95) );
  NAND2_X1 U170 ( .A1(n179), .A2(n79), .ZN(n13) );
  NAND2_X1 U171 ( .A1(n99), .A2(n62), .ZN(n9) );
  INV_X1 U172 ( .A(n61), .ZN(n99) );
  NAND2_X1 U173 ( .A1(n183), .A2(n87), .ZN(n15) );
  NAND2_X1 U174 ( .A1(n184), .A2(n71), .ZN(n11) );
  NAND2_X1 U175 ( .A1(n100), .A2(n66), .ZN(n10) );
  INV_X1 U176 ( .A(n65), .ZN(n100) );
  NAND2_X1 U177 ( .A1(n102), .A2(n74), .ZN(n12) );
  INV_X1 U178 ( .A(n73), .ZN(n102) );
  XNOR2_X1 U179 ( .A(n13), .B(n80), .ZN(SUM[3]) );
  XOR2_X1 U180 ( .A(n14), .B(n83), .Z(SUM[2]) );
  XNOR2_X1 U181 ( .A(n15), .B(n88), .ZN(SUM[1]) );
  XNOR2_X1 U182 ( .A(n38), .B(n4), .ZN(SUM[12]) );
  OR2_X1 U183 ( .A1(A[3]), .A2(B[3]), .ZN(n179) );
  NOR2_X1 U184 ( .A1(A[2]), .A2(B[2]), .ZN(n81) );
  XOR2_X1 U185 ( .A(n49), .B(n6), .Z(SUM[10]) );
  NAND2_X1 U186 ( .A1(A[11]), .A2(B[11]), .ZN(n40) );
  NAND2_X1 U187 ( .A1(n164), .A2(n18), .ZN(n1) );
  XNOR2_X1 U188 ( .A(n60), .B(n8), .ZN(SUM[8]) );
  NOR2_X1 U189 ( .A1(A[6]), .A2(B[6]), .ZN(n65) );
  NOR2_X1 U190 ( .A1(A[4]), .A2(B[4]), .ZN(n73) );
  NAND2_X1 U191 ( .A1(A[7]), .A2(B[7]), .ZN(n62) );
  NAND2_X1 U192 ( .A1(A[2]), .A2(B[2]), .ZN(n82) );
  OR2_X1 U193 ( .A1(A[1]), .A2(B[1]), .ZN(n183) );
  NAND2_X1 U194 ( .A1(A[9]), .A2(B[9]), .ZN(n53) );
  NAND2_X1 U195 ( .A1(A[5]), .A2(B[5]), .ZN(n71) );
  NAND2_X1 U196 ( .A1(A[1]), .A2(B[1]), .ZN(n87) );
  NAND2_X1 U197 ( .A1(A[0]), .A2(B[0]), .ZN(n90) );
  NAND2_X1 U198 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  OR2_X1 U199 ( .A1(A[5]), .A2(B[5]), .ZN(n184) );
  NAND2_X1 U200 ( .A1(A[6]), .A2(B[6]), .ZN(n66) );
  NAND2_X1 U201 ( .A1(A[4]), .A2(B[4]), .ZN(n74) );
  XOR2_X1 U202 ( .A(n63), .B(n9), .Z(SUM[7]) );
  NAND2_X1 U203 ( .A1(n94), .A2(n37), .ZN(n4) );
  INV_X1 U204 ( .A(n64), .ZN(n63) );
  AOI21_X1 U205 ( .B1(n56), .B2(n64), .A(n57), .ZN(n55) );
  AND2_X1 U206 ( .A1(A[14]), .A2(B[14]), .ZN(n185) );
  INV_X1 U207 ( .A(n28), .ZN(n30) );
  NAND2_X1 U208 ( .A1(A[12]), .A2(B[12]), .ZN(n37) );
  NOR2_X1 U209 ( .A1(n58), .A2(n61), .ZN(n56) );
  OAI21_X1 U210 ( .B1(n165), .B2(n62), .A(n59), .ZN(n57) );
  NAND2_X1 U211 ( .A1(A[8]), .A2(B[8]), .ZN(n59) );
  NAND2_X1 U212 ( .A1(A[15]), .A2(B[15]), .ZN(n18) );
  INV_X1 U213 ( .A(n172), .ZN(n94) );
  NOR2_X1 U214 ( .A1(n172), .A2(n39), .ZN(n34) );
  XOR2_X1 U215 ( .A(n10), .B(n67), .Z(SUM[6]) );
  OAI21_X1 U216 ( .B1(n67), .B2(n65), .A(n66), .ZN(n64) );
  AOI21_X1 U217 ( .B1(n184), .B2(n72), .A(n69), .ZN(n67) );
  XNOR2_X1 U218 ( .A(n11), .B(n72), .ZN(SUM[5]) );
  OAI21_X1 U219 ( .B1(n75), .B2(n73), .A(n74), .ZN(n72) );
  NAND2_X1 U220 ( .A1(n181), .A2(n25), .ZN(n2) );
  NAND2_X1 U221 ( .A1(n181), .A2(n173), .ZN(n20) );
  AOI21_X1 U222 ( .B1(n181), .B2(n30), .A(n185), .ZN(n21) );
  OAI21_X1 U223 ( .B1(n36), .B2(n40), .A(n37), .ZN(n35) );
  NAND2_X1 U224 ( .A1(A[14]), .A2(B[14]), .ZN(n25) );
  NOR2_X1 U225 ( .A1(A[13]), .A2(B[13]), .ZN(n27) );
  XOR2_X1 U226 ( .A(n12), .B(n75), .Z(SUM[4]) );
  OAI21_X1 U227 ( .B1(n41), .B2(n39), .A(n40), .ZN(n38) );
  NAND2_X1 U228 ( .A1(A[3]), .A2(B[3]), .ZN(n79) );
  XNOR2_X1 U229 ( .A(n19), .B(n1), .ZN(SUM[15]) );
  NAND2_X1 U230 ( .A1(n174), .A2(n48), .ZN(n6) );
  INV_X1 U231 ( .A(n170), .ZN(n41) );
  NAND2_X1 U232 ( .A1(n182), .A2(n180), .ZN(n43) );
  OAI21_X1 U233 ( .B1(n55), .B2(n43), .A(n168), .ZN(n42) );
  AOI21_X1 U234 ( .B1(n182), .B2(n51), .A(n175), .ZN(n44) );
  XNOR2_X1 U235 ( .A(n26), .B(n2), .ZN(SUM[14]) );
  OAI21_X1 U236 ( .B1(n177), .B2(n27), .A(n28), .ZN(n26) );
  OAI21_X1 U237 ( .B1(n176), .B2(n20), .A(n21), .ZN(n19) );
endmodule


module layer1_8_4_8_16_datapath_M8_N4_T16_P8_7 ( clk, clear_acc, data_out_x, 
        data_out, data_out_w, data_out_b, wr_en_y, m_valid, m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [3:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N27, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, n1, n2, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n87, n104, n113, n114, n115, n116, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(clear_acc), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n223), .CK(clk), .Q(n21) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n224), .CK(clk), .Q(n22) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n225), .CK(clk), .Q(n23) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n226), .CK(clk), .Q(n24) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n227), .CK(clk), .Q(n25) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n228), .CK(clk), .Q(n26) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n229), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n230), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n231), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n232), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n233), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n234), .CK(clk), .Q(n34) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n235), .CK(clk), .Q(n35) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n236), .CK(clk), .Q(n36) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n237), .CK(clk), .Q(n37) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n238), .CK(clk), .Q(n39) );
  DFF_X1 \f_reg[0]  ( .D(n113), .CK(clk), .Q(n61), .QN(n212) );
  DFF_X1 \f_reg[1]  ( .D(n104), .CK(clk), .Q(n59), .QN(n213) );
  DFF_X1 \f_reg[2]  ( .D(n87), .CK(clk), .Q(n57), .QN(n214) );
  DFF_X1 \f_reg[3]  ( .D(n85), .CK(clk), .Q(f[3]), .QN(n65) );
  DFF_X1 \f_reg[4]  ( .D(n84), .CK(clk), .Q(f[4]), .QN(n66) );
  DFF_X1 \f_reg[5]  ( .D(n83), .CK(clk), .Q(f[5]), .QN(n67) );
  DFF_X1 \f_reg[6]  ( .D(n82), .CK(clk), .Q(f[6]), .QN(n68) );
  DFF_X1 \f_reg[7]  ( .D(n81), .CK(clk), .Q(f[7]), .QN(n215) );
  DFF_X1 \f_reg[8]  ( .D(n80), .CK(clk), .Q(f[8]), .QN(n216) );
  DFF_X1 \f_reg[9]  ( .D(n79), .CK(clk), .Q(f[9]), .QN(n217) );
  DFF_X1 \f_reg[10]  ( .D(n78), .CK(clk), .Q(n49), .QN(n218) );
  DFF_X1 \f_reg[11]  ( .D(n1), .CK(clk), .Q(n48), .QN(n219) );
  DFF_X1 \f_reg[12]  ( .D(n77), .CK(clk), .Q(n46), .QN(n220) );
  DFF_X1 \f_reg[13]  ( .D(n76), .CK(clk), .Q(n44), .QN(n221) );
  DFF_X1 \f_reg[14]  ( .D(n2), .CK(clk), .Q(n43), .QN(n222) );
  DFF_X1 \f_reg[15]  ( .D(n75), .CK(clk), .Q(f[15]), .QN(n73) );
  DFF_X1 \data_out_reg[15]  ( .D(n115), .CK(clk), .Q(data_out[15]), .QN(n195)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n116), .CK(clk), .Q(data_out[14]), .QN(n194)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n166), .CK(clk), .Q(data_out[13]), .QN(n193)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n167), .CK(clk), .Q(data_out[12]), .QN(n192)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n168), .CK(clk), .Q(data_out[11]), .QN(n191)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n169), .CK(clk), .Q(data_out[10]), .QN(n190)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n170), .CK(clk), .Q(data_out[9]), .QN(n189) );
  DFF_X1 \data_out_reg[8]  ( .D(n171), .CK(clk), .Q(data_out[8]), .QN(n188) );
  DFF_X1 \data_out_reg[7]  ( .D(n172), .CK(clk), .Q(data_out[7]), .QN(n187) );
  DFF_X1 \data_out_reg[6]  ( .D(n173), .CK(clk), .Q(data_out[6]), .QN(n186) );
  DFF_X1 \data_out_reg[5]  ( .D(n174), .CK(clk), .Q(data_out[5]), .QN(n185) );
  DFF_X1 \data_out_reg[4]  ( .D(n175), .CK(clk), .Q(data_out[4]), .QN(n184) );
  DFF_X1 \data_out_reg[3]  ( .D(n176), .CK(clk), .Q(data_out[3]), .QN(n183) );
  DFF_X1 \data_out_reg[2]  ( .D(n177), .CK(clk), .Q(data_out[2]), .QN(n182) );
  DFF_X1 \data_out_reg[1]  ( .D(n178), .CK(clk), .Q(data_out[1]), .QN(n181) );
  DFF_X1 \data_out_reg[0]  ( .D(n179), .CK(clk), .Q(data_out[0]), .QN(n180) );
  layer1_8_4_8_16_datapath_M8_N4_T16_P8_7_DW_mult_tc_1 mult_183 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer1_8_4_8_16_datapath_M8_N4_T16_P8_7_DW01_add_2 add_184 ( .A({n202, n201, 
        n200, n199, n198, n197, n211, n210, n209, n208, n207, n206, n205, n204, 
        n203, n196}), .B({f[15], n43, n44, n46, n48, n49, f[9:3], n57, n59, 
        n61}), .CI(1'b0), .SUM(adder) );
  DFF_X2 delay_reg ( .D(N27), .CK(clk), .Q(n11), .QN(n239) );
  NAND3_X1 U3 ( .A1(n5), .A2(n4), .A3(n6), .ZN(n1) );
  NAND3_X1 U4 ( .A1(n14), .A2(n13), .A3(n15), .ZN(n2) );
  NAND2_X1 U5 ( .A1(data_out_b[11]), .A2(clear_acc), .ZN(n4) );
  NAND2_X1 U6 ( .A1(adder[11]), .A2(n16), .ZN(n5) );
  NAND2_X1 U8 ( .A1(n63), .A2(n48), .ZN(n6) );
  AND2_X1 U9 ( .A1(n10), .A2(n8), .ZN(n7) );
  NAND2_X1 U10 ( .A1(n9), .A2(n7), .ZN(n75) );
  NAND2_X1 U11 ( .A1(data_out_b[15]), .A2(clear_acc), .ZN(n8) );
  NAND2_X1 U12 ( .A1(adder[15]), .A2(n16), .ZN(n9) );
  NAND2_X1 U13 ( .A1(n63), .A2(f[15]), .ZN(n10) );
  MUX2_X2 U14 ( .A(N39), .B(n26), .S(n11), .Z(n197) );
  CLKBUF_X1 U15 ( .A(N39), .Z(n12) );
  MUX2_X2 U16 ( .A(n23), .B(N42), .S(n239), .Z(n200) );
  MUX2_X2 U17 ( .A(n25), .B(N40), .S(n239), .Z(n198) );
  NAND2_X1 U18 ( .A1(data_out_b[14]), .A2(clear_acc), .ZN(n13) );
  NAND2_X1 U19 ( .A1(adder[14]), .A2(n16), .ZN(n14) );
  NAND2_X1 U20 ( .A1(n63), .A2(n43), .ZN(n15) );
  MUX2_X2 U21 ( .A(n24), .B(N41), .S(n239), .Z(n199) );
  MUX2_X2 U22 ( .A(n28), .B(N37), .S(n239), .Z(n210) );
  MUX2_X2 U23 ( .A(n22), .B(N43), .S(n239), .Z(n201) );
  AND2_X2 U24 ( .A1(n42), .A2(n17), .ZN(n16) );
  INV_X1 U25 ( .A(n42), .ZN(n63) );
  INV_X1 U26 ( .A(clear_acc), .ZN(n17) );
  NAND2_X1 U27 ( .A1(n114), .A2(N27), .ZN(n241) );
  INV_X1 U28 ( .A(wr_en_y), .ZN(n114) );
  INV_X1 U29 ( .A(n20), .ZN(n38) );
  OAI22_X1 U30 ( .A1(n183), .A2(n241), .B1(n65), .B2(n240), .ZN(n176) );
  OAI22_X1 U31 ( .A1(n184), .A2(n241), .B1(n66), .B2(n240), .ZN(n175) );
  OAI22_X1 U32 ( .A1(n185), .A2(n241), .B1(n67), .B2(n240), .ZN(n174) );
  OAI22_X1 U33 ( .A1(n186), .A2(n241), .B1(n68), .B2(n240), .ZN(n173) );
  OAI22_X1 U34 ( .A1(n187), .A2(n241), .B1(n215), .B2(n240), .ZN(n172) );
  OAI22_X1 U35 ( .A1(n188), .A2(n241), .B1(n216), .B2(n240), .ZN(n171) );
  OAI22_X1 U36 ( .A1(n189), .A2(n241), .B1(n217), .B2(n240), .ZN(n170) );
  AND3_X1 U37 ( .A1(sel[1]), .A2(sel[2]), .A3(sel[0]), .ZN(n19) );
  INV_X1 U38 ( .A(m_ready), .ZN(n18) );
  NAND2_X1 U39 ( .A1(m_valid), .A2(n18), .ZN(n40) );
  OAI21_X1 U40 ( .B1(sel[3]), .B2(n19), .A(n40), .ZN(N27) );
  NAND2_X1 U41 ( .A1(clear_acc_delay), .A2(n239), .ZN(n20) );
  MUX2_X1 U42 ( .A(n21), .B(N44), .S(n38), .Z(n223) );
  MUX2_X1 U43 ( .A(n21), .B(N44), .S(n239), .Z(n202) );
  MUX2_X1 U44 ( .A(n22), .B(N43), .S(n38), .Z(n224) );
  MUX2_X1 U45 ( .A(n23), .B(N42), .S(n38), .Z(n225) );
  MUX2_X1 U46 ( .A(n24), .B(N41), .S(n38), .Z(n226) );
  MUX2_X1 U47 ( .A(n25), .B(N40), .S(n38), .Z(n227) );
  MUX2_X1 U48 ( .A(n26), .B(n12), .S(n38), .Z(n228) );
  MUX2_X1 U49 ( .A(n27), .B(N38), .S(n38), .Z(n229) );
  MUX2_X1 U50 ( .A(n27), .B(N38), .S(n239), .Z(n211) );
  MUX2_X1 U51 ( .A(n28), .B(N37), .S(n38), .Z(n230) );
  MUX2_X1 U52 ( .A(n29), .B(N36), .S(n38), .Z(n231) );
  MUX2_X1 U53 ( .A(n29), .B(N36), .S(n239), .Z(n209) );
  MUX2_X1 U54 ( .A(n32), .B(N35), .S(n38), .Z(n232) );
  MUX2_X1 U55 ( .A(n32), .B(N35), .S(n239), .Z(n208) );
  MUX2_X1 U56 ( .A(n33), .B(N34), .S(n38), .Z(n233) );
  MUX2_X1 U57 ( .A(n33), .B(N34), .S(n239), .Z(n207) );
  MUX2_X1 U58 ( .A(n34), .B(N33), .S(n38), .Z(n234) );
  MUX2_X1 U59 ( .A(n34), .B(N33), .S(n239), .Z(n206) );
  MUX2_X1 U60 ( .A(n35), .B(N32), .S(n38), .Z(n235) );
  MUX2_X1 U61 ( .A(n35), .B(N32), .S(n239), .Z(n205) );
  MUX2_X1 U62 ( .A(n36), .B(N31), .S(n38), .Z(n236) );
  MUX2_X1 U63 ( .A(n36), .B(N31), .S(n239), .Z(n204) );
  MUX2_X1 U64 ( .A(n37), .B(N30), .S(n38), .Z(n237) );
  MUX2_X1 U65 ( .A(n37), .B(N30), .S(n239), .Z(n203) );
  MUX2_X1 U66 ( .A(n39), .B(N29), .S(n38), .Z(n238) );
  MUX2_X1 U67 ( .A(n39), .B(N29), .S(n239), .Z(n196) );
  INV_X1 U68 ( .A(n40), .ZN(n41) );
  OAI21_X1 U69 ( .B1(n41), .B2(n11), .A(n17), .ZN(n42) );
  AOI222_X1 U70 ( .A1(data_out_b[13]), .A2(clear_acc), .B1(adder[13]), .B2(n16), .C1(n63), .C2(n44), .ZN(n45) );
  INV_X1 U71 ( .A(n45), .ZN(n76) );
  AOI222_X1 U72 ( .A1(data_out_b[12]), .A2(clear_acc), .B1(adder[12]), .B2(n16), .C1(n63), .C2(n46), .ZN(n47) );
  INV_X1 U73 ( .A(n47), .ZN(n77) );
  AOI222_X1 U74 ( .A1(data_out_b[10]), .A2(clear_acc), .B1(adder[10]), .B2(n16), .C1(n63), .C2(n49), .ZN(n50) );
  INV_X1 U75 ( .A(n50), .ZN(n78) );
  AOI222_X1 U76 ( .A1(data_out_b[8]), .A2(clear_acc), .B1(adder[8]), .B2(n16), 
        .C1(n63), .C2(f[8]), .ZN(n51) );
  INV_X1 U77 ( .A(n51), .ZN(n80) );
  AOI222_X1 U78 ( .A1(data_out_b[7]), .A2(clear_acc), .B1(adder[7]), .B2(n16), 
        .C1(n63), .C2(f[7]), .ZN(n52) );
  INV_X1 U79 ( .A(n52), .ZN(n81) );
  AOI222_X1 U80 ( .A1(data_out_b[6]), .A2(clear_acc), .B1(adder[6]), .B2(n16), 
        .C1(n63), .C2(f[6]), .ZN(n53) );
  INV_X1 U81 ( .A(n53), .ZN(n82) );
  AOI222_X1 U82 ( .A1(data_out_b[5]), .A2(clear_acc), .B1(adder[5]), .B2(n16), 
        .C1(n63), .C2(f[5]), .ZN(n54) );
  INV_X1 U83 ( .A(n54), .ZN(n83) );
  AOI222_X1 U84 ( .A1(data_out_b[4]), .A2(clear_acc), .B1(adder[4]), .B2(n16), 
        .C1(n63), .C2(f[4]), .ZN(n55) );
  INV_X1 U85 ( .A(n55), .ZN(n84) );
  AOI222_X1 U86 ( .A1(data_out_b[3]), .A2(clear_acc), .B1(adder[3]), .B2(n16), 
        .C1(n63), .C2(f[3]), .ZN(n56) );
  INV_X1 U87 ( .A(n56), .ZN(n85) );
  AOI222_X1 U88 ( .A1(data_out_b[2]), .A2(clear_acc), .B1(adder[2]), .B2(n16), 
        .C1(n63), .C2(n57), .ZN(n58) );
  INV_X1 U89 ( .A(n58), .ZN(n87) );
  AOI222_X1 U90 ( .A1(data_out_b[1]), .A2(clear_acc), .B1(adder[1]), .B2(n16), 
        .C1(n63), .C2(n59), .ZN(n60) );
  INV_X1 U91 ( .A(n60), .ZN(n104) );
  AOI222_X1 U92 ( .A1(data_out_b[0]), .A2(clear_acc), .B1(adder[0]), .B2(n16), 
        .C1(n63), .C2(n61), .ZN(n62) );
  INV_X1 U93 ( .A(n62), .ZN(n113) );
  AOI222_X1 U94 ( .A1(data_out_b[9]), .A2(clear_acc), .B1(adder[9]), .B2(n16), 
        .C1(n63), .C2(f[9]), .ZN(n64) );
  INV_X1 U95 ( .A(n64), .ZN(n79) );
  NOR4_X1 U96 ( .A1(n48), .A2(n46), .A3(n44), .A4(n43), .ZN(n72) );
  NOR4_X1 U97 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n49), .ZN(n71) );
  NAND4_X1 U98 ( .A1(n68), .A2(n67), .A3(n66), .A4(n65), .ZN(n69) );
  NOR4_X1 U99 ( .A1(n69), .A2(n61), .A3(n59), .A4(n57), .ZN(n70) );
  NAND3_X1 U100 ( .A1(n72), .A2(n71), .A3(n70), .ZN(n74) );
  NAND3_X1 U101 ( .A1(wr_en_y), .A2(n74), .A3(n73), .ZN(n240) );
  OAI22_X1 U102 ( .A1(n180), .A2(n241), .B1(n212), .B2(n240), .ZN(n179) );
  OAI22_X1 U103 ( .A1(n181), .A2(n241), .B1(n213), .B2(n240), .ZN(n178) );
  OAI22_X1 U104 ( .A1(n182), .A2(n241), .B1(n214), .B2(n240), .ZN(n177) );
  OAI22_X1 U105 ( .A1(n190), .A2(n241), .B1(n218), .B2(n240), .ZN(n169) );
  OAI22_X1 U106 ( .A1(n191), .A2(n241), .B1(n219), .B2(n240), .ZN(n168) );
  OAI22_X1 U107 ( .A1(n192), .A2(n241), .B1(n220), .B2(n240), .ZN(n167) );
  OAI22_X1 U108 ( .A1(n193), .A2(n241), .B1(n221), .B2(n240), .ZN(n166) );
  OAI22_X1 U109 ( .A1(n194), .A2(n241), .B1(n222), .B2(n240), .ZN(n116) );
  OAI22_X1 U110 ( .A1(n195), .A2(n241), .B1(n73), .B2(n240), .ZN(n115) );
endmodule


module layer1_8_4_8_16_datapath_M8_N4_T16_P8_6_DW_mult_tc_1 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n9, n12, n13, n16, n18, n19, n21, n23, n25, n27, n29, n31,
         n32, n34, n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n50,
         n51, n53, n54, n55, n56, n57, n58, n59, n62, n63, n64, n65, n67, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n89, n90, n91, n93, n95, n96, n97, n98, n99, n103,
         n104, n105, n106, n107, n109, n111, n112, n113, n114, n115, n117,
         n119, n120, n122, n125, n127, n128, n131, n133, n135, n139, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n237, n245, n247, n249, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n418, n419, n420, n421, n422, n423, n424, n426,
         n427, n429, n430, n433, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U148 ( .A(n265), .B(n144), .Z(n145) );
  XOR2_X1 U150 ( .A(n271), .B(n146), .Z(n147) );
  XOR2_X1 U152 ( .A(n301), .B(n148), .Z(n149) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n263), .CI(n291), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n252), .B(n317), .CO(n173), .S(n174) );
  FA_X1 U167 ( .A(n180), .B(n187), .CI(n178), .CO(n175), .S(n176) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U169 ( .A(n193), .B(n282), .CI(n191), .CO(n179), .S(n180) );
  FA_X1 U170 ( .A(n268), .B(n292), .CI(n274), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U172 ( .A(n197), .B(n190), .CI(n188), .CO(n185), .S(n186) );
  FA_X1 U173 ( .A(n199), .B(n201), .CI(n192), .CO(n187), .S(n188) );
  FA_X1 U174 ( .A(n275), .B(n293), .CI(n194), .CO(n189), .S(n190) );
  FA_X1 U175 ( .A(n305), .B(n253), .CI(n283), .CO(n191), .S(n192) );
  HA_X1 U176 ( .A(n319), .B(n269), .CO(n193), .S(n194) );
  FA_X1 U177 ( .A(n205), .B(n200), .CI(n198), .CO(n195), .S(n196) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U179 ( .A(n284), .B(n276), .CI(n294), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n320), .B(n270), .CI(n306), .CO(n201), .S(n202) );
  FA_X1 U181 ( .A(n208), .B(n213), .CI(n206), .CO(n203), .S(n204) );
  FA_X1 U182 ( .A(n210), .B(n307), .CI(n215), .CO(n205), .S(n206) );
  FA_X1 U183 ( .A(n295), .B(n285), .CI(n254), .CO(n207), .S(n208) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U185 ( .A(n216), .B(n219), .CI(n214), .CO(n211), .S(n212) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n322), .B(n278), .CI(n308), .CO(n215), .S(n216) );
  FA_X1 U188 ( .A(n225), .B(n222), .CI(n220), .CO(n217), .S(n218) );
  FA_X1 U189 ( .A(n255), .B(n309), .CI(n297), .CO(n219), .S(n220) );
  HA_X1 U190 ( .A(n287), .B(n323), .CO(n221), .S(n222) );
  FA_X1 U191 ( .A(n229), .B(n298), .CI(n226), .CO(n223), .S(n224) );
  FA_X1 U192 ( .A(n310), .B(n288), .CI(n324), .CO(n225), .S(n226) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  HA_X1 U194 ( .A(n311), .B(n325), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n326), .B(n300), .CI(n312), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  CLKBUF_X1 U414 ( .A(n494), .Z(n535) );
  OAI21_X1 U415 ( .B1(n515), .B2(n89), .A(n90), .ZN(n490) );
  XOR2_X1 U416 ( .A(n578), .B(a[12]), .Z(n37) );
  AOI21_X1 U417 ( .B1(n556), .B2(n104), .A(n521), .ZN(n491) );
  CLKBUF_X3 U418 ( .A(n16), .Z(n561) );
  BUF_X1 U419 ( .A(n566), .Z(n518) );
  NAND2_X1 U420 ( .A1(n429), .A2(n27), .ZN(n29) );
  NOR2_X1 U421 ( .A1(n228), .A2(n231), .ZN(n105) );
  AND2_X1 U422 ( .A1(n224), .A2(n227), .ZN(n521) );
  BUF_X1 U423 ( .A(n567), .Z(n511) );
  OR2_X1 U424 ( .A1(n329), .A2(n258), .ZN(n492) );
  NOR2_X1 U425 ( .A1(n196), .A2(n203), .ZN(n85) );
  OAI21_X1 U426 ( .B1(n82), .B2(n86), .A(n83), .ZN(n493) );
  OAI21_X1 U427 ( .B1(n99), .B2(n97), .A(n98), .ZN(n494) );
  AOI21_X1 U428 ( .B1(n80), .B2(n490), .A(n493), .ZN(n495) );
  BUF_X2 U429 ( .A(n12), .Z(n545) );
  INV_X1 U430 ( .A(n569), .ZN(n496) );
  INV_X2 U431 ( .A(n570), .ZN(n569) );
  XOR2_X1 U432 ( .A(n511), .B(n419), .Z(n402) );
  INV_X1 U433 ( .A(n521), .ZN(n103) );
  OR2_X2 U434 ( .A1(n224), .A2(n227), .ZN(n556) );
  INV_X1 U435 ( .A(n27), .ZN(n497) );
  XNOR2_X1 U436 ( .A(n495), .B(n498), .ZN(product[12]) );
  AND2_X1 U437 ( .A1(n506), .A2(n79), .ZN(n498) );
  BUF_X1 U438 ( .A(n107), .Z(n512) );
  CLKBUF_X1 U439 ( .A(n74), .Z(n499) );
  CLKBUF_X1 U440 ( .A(n105), .Z(n500) );
  XNOR2_X1 U441 ( .A(n576), .B(a[8]), .ZN(n429) );
  BUF_X2 U442 ( .A(n516), .Z(n501) );
  CLKBUF_X1 U443 ( .A(n516), .Z(n562) );
  XNOR2_X1 U444 ( .A(n543), .B(n502), .ZN(product[9]) );
  AND2_X1 U445 ( .A1(n513), .A2(n90), .ZN(n502) );
  XOR2_X1 U446 ( .A(n511), .B(b[10]), .Z(n398) );
  BUF_X2 U447 ( .A(n566), .Z(n520) );
  OAI21_X1 U448 ( .B1(n515), .B2(n89), .A(n90), .ZN(n503) );
  CLKBUF_X1 U449 ( .A(n18), .Z(n504) );
  CLKBUF_X3 U450 ( .A(n18), .Z(n505) );
  OR2_X1 U451 ( .A1(n176), .A2(n185), .ZN(n506) );
  XNOR2_X1 U452 ( .A(n574), .B(a[6]), .ZN(n430) );
  OAI21_X1 U453 ( .B1(n512), .B2(n500), .A(n106), .ZN(n507) );
  BUF_X2 U454 ( .A(n12), .Z(n508) );
  OR2_X2 U455 ( .A1(n509), .A2(n542), .ZN(n34) );
  XNOR2_X1 U456 ( .A(n577), .B(a[10]), .ZN(n509) );
  INV_X1 U457 ( .A(n542), .ZN(n32) );
  XNOR2_X1 U458 ( .A(n510), .B(n166), .ZN(n164) );
  XNOR2_X1 U459 ( .A(n177), .B(n168), .ZN(n510) );
  XOR2_X1 U460 ( .A(n511), .B(b[9]), .Z(n399) );
  BUF_X1 U461 ( .A(n566), .Z(n519) );
  OR2_X1 U462 ( .A1(n204), .A2(n211), .ZN(n513) );
  XNOR2_X1 U463 ( .A(n573), .B(a[4]), .ZN(n550) );
  INV_X1 U464 ( .A(n548), .ZN(n514) );
  INV_X1 U465 ( .A(n548), .ZN(n21) );
  AOI21_X1 U466 ( .B1(n96), .B2(n552), .A(n93), .ZN(n515) );
  XOR2_X1 U467 ( .A(n567), .B(a[2]), .Z(n516) );
  NOR2_X1 U468 ( .A1(n186), .A2(n195), .ZN(n517) );
  NOR2_X1 U469 ( .A1(n186), .A2(n195), .ZN(n82) );
  INV_X2 U470 ( .A(n578), .ZN(n577) );
  INV_X1 U471 ( .A(n567), .ZN(n566) );
  INV_X2 U472 ( .A(n541), .ZN(n27) );
  CLKBUF_X3 U473 ( .A(n19), .Z(n522) );
  OR2_X1 U474 ( .A1(n23), .A2(n359), .ZN(n523) );
  OR2_X1 U475 ( .A1(n358), .A2(n21), .ZN(n524) );
  NAND2_X1 U476 ( .A1(n523), .A2(n524), .ZN(n283) );
  AOI21_X1 U477 ( .B1(n556), .B2(n507), .A(n521), .ZN(n525) );
  OAI21_X1 U478 ( .B1(n91), .B2(n89), .A(n90), .ZN(n526) );
  XOR2_X1 U479 ( .A(n567), .B(a[2]), .Z(n9) );
  XOR2_X1 U480 ( .A(n170), .B(n172), .Z(n527) );
  XOR2_X1 U481 ( .A(n527), .B(n179), .Z(n166) );
  NAND2_X1 U482 ( .A1(n170), .A2(n172), .ZN(n528) );
  NAND2_X1 U483 ( .A1(n170), .A2(n179), .ZN(n529) );
  NAND2_X1 U484 ( .A1(n172), .A2(n179), .ZN(n530) );
  NAND3_X1 U485 ( .A1(n528), .A2(n529), .A3(n530), .ZN(n165) );
  NAND2_X1 U486 ( .A1(n177), .A2(n168), .ZN(n531) );
  NAND2_X1 U487 ( .A1(n177), .A2(n166), .ZN(n532) );
  NAND2_X1 U488 ( .A1(n168), .A2(n166), .ZN(n533) );
  NAND3_X1 U489 ( .A1(n531), .A2(n532), .A3(n533), .ZN(n163) );
  AOI21_X1 U490 ( .B1(n503), .B2(n80), .A(n81), .ZN(n534) );
  NOR2_X2 U491 ( .A1(n164), .A2(n175), .ZN(n75) );
  XNOR2_X1 U492 ( .A(n526), .B(n51), .ZN(product[10]) );
  CLKBUF_X1 U493 ( .A(n534), .Z(n536) );
  INV_X1 U494 ( .A(n563), .ZN(n537) );
  INV_X1 U495 ( .A(n537), .ZN(n538) );
  INV_X1 U496 ( .A(n537), .ZN(n539) );
  INV_X1 U497 ( .A(n537), .ZN(n540) );
  XNOR2_X1 U498 ( .A(n574), .B(a[8]), .ZN(n541) );
  XNOR2_X1 U499 ( .A(n570), .B(a[2]), .ZN(n549) );
  INV_X1 U500 ( .A(n570), .ZN(n568) );
  XNOR2_X1 U501 ( .A(n576), .B(a[10]), .ZN(n542) );
  BUF_X1 U502 ( .A(n12), .Z(n544) );
  XNOR2_X1 U503 ( .A(n567), .B(n249), .ZN(n433) );
  NAND2_X2 U504 ( .A1(n430), .A2(n514), .ZN(n23) );
  CLKBUF_X1 U505 ( .A(n515), .Z(n543) );
  XOR2_X1 U506 ( .A(n570), .B(a[4]), .Z(n16) );
  INV_X2 U507 ( .A(n576), .ZN(n575) );
  NAND2_X1 U508 ( .A1(n433), .A2(n540), .ZN(n546) );
  NAND2_X1 U509 ( .A1(n433), .A2(n540), .ZN(n547) );
  AOI21_X1 U510 ( .B1(n490), .B2(n80), .A(n493), .ZN(n45) );
  XNOR2_X1 U511 ( .A(n573), .B(a[6]), .ZN(n548) );
  NAND2_X1 U512 ( .A1(n9), .A2(n549), .ZN(n12) );
  NAND2_X1 U513 ( .A1(n550), .A2(n16), .ZN(n18) );
  BUF_X1 U514 ( .A(n43), .Z(n564) );
  NAND2_X1 U515 ( .A1(n551), .A2(n69), .ZN(n47) );
  INV_X1 U516 ( .A(n73), .ZN(n71) );
  AOI21_X1 U517 ( .B1(n499), .B2(n551), .A(n67), .ZN(n65) );
  INV_X1 U518 ( .A(n69), .ZN(n67) );
  INV_X1 U519 ( .A(n74), .ZN(n72) );
  INV_X1 U520 ( .A(n95), .ZN(n93) );
  NAND2_X1 U521 ( .A1(n128), .A2(n86), .ZN(n51) );
  INV_X1 U522 ( .A(n85), .ZN(n128) );
  NAND2_X1 U523 ( .A1(n125), .A2(n76), .ZN(n48) );
  INV_X1 U524 ( .A(n75), .ZN(n125) );
  OR2_X1 U525 ( .A1(n152), .A2(n163), .ZN(n551) );
  OAI21_X1 U526 ( .B1(n75), .B2(n79), .A(n76), .ZN(n74) );
  NAND2_X1 U527 ( .A1(n127), .A2(n83), .ZN(n50) );
  NOR2_X1 U528 ( .A1(n75), .A2(n78), .ZN(n73) );
  NAND2_X1 U529 ( .A1(n152), .A2(n163), .ZN(n69) );
  NAND2_X1 U530 ( .A1(n552), .A2(n95), .ZN(n53) );
  AOI21_X1 U531 ( .B1(n555), .B2(n112), .A(n109), .ZN(n107) );
  OAI21_X1 U532 ( .B1(n113), .B2(n115), .A(n114), .ZN(n112) );
  AOI21_X1 U533 ( .B1(n554), .B2(n120), .A(n117), .ZN(n115) );
  INV_X1 U534 ( .A(n119), .ZN(n117) );
  NOR2_X1 U535 ( .A1(n176), .A2(n185), .ZN(n78) );
  OAI21_X1 U536 ( .B1(n107), .B2(n105), .A(n106), .ZN(n104) );
  INV_X1 U537 ( .A(n122), .ZN(n120) );
  XNOR2_X1 U538 ( .A(n59), .B(n120), .ZN(product[2]) );
  NAND2_X1 U539 ( .A1(n554), .A2(n119), .ZN(n59) );
  NAND2_X1 U540 ( .A1(n176), .A2(n185), .ZN(n79) );
  XOR2_X1 U541 ( .A(n58), .B(n115), .Z(product[3]) );
  NAND2_X1 U542 ( .A1(n164), .A2(n175), .ZN(n76) );
  NAND2_X1 U543 ( .A1(n196), .A2(n203), .ZN(n86) );
  NAND2_X1 U544 ( .A1(n212), .A2(n217), .ZN(n95) );
  OR2_X1 U545 ( .A1(n212), .A2(n217), .ZN(n552) );
  NAND2_X1 U546 ( .A1(n204), .A2(n211), .ZN(n90) );
  XNOR2_X1 U547 ( .A(n63), .B(n46), .ZN(product[15]) );
  NAND2_X1 U548 ( .A1(n553), .A2(n62), .ZN(n46) );
  NAND2_X1 U549 ( .A1(n73), .A2(n551), .ZN(n64) );
  NAND2_X1 U550 ( .A1(n131), .A2(n98), .ZN(n54) );
  INV_X1 U551 ( .A(n97), .ZN(n131) );
  NAND2_X1 U552 ( .A1(n133), .A2(n106), .ZN(n56) );
  INV_X1 U553 ( .A(n105), .ZN(n133) );
  OR2_X1 U554 ( .A1(n151), .A2(n139), .ZN(n553) );
  OR2_X1 U555 ( .A1(n328), .A2(n314), .ZN(n554) );
  NOR2_X1 U556 ( .A1(n218), .A2(n223), .ZN(n97) );
  NAND2_X1 U557 ( .A1(n218), .A2(n223), .ZN(n98) );
  NAND2_X1 U558 ( .A1(n228), .A2(n231), .ZN(n106) );
  OR2_X1 U559 ( .A1(n232), .A2(n233), .ZN(n555) );
  AND2_X1 U560 ( .A1(n492), .A2(n122), .ZN(product[1]) );
  NAND2_X1 U561 ( .A1(n433), .A2(n540), .ZN(n6) );
  OR2_X1 U562 ( .A1(n564), .A2(n496), .ZN(n392) );
  AND2_X1 U563 ( .A1(n565), .A2(n542), .ZN(n270) );
  AND2_X1 U564 ( .A1(n565), .A2(n548), .ZN(n288) );
  XNOR2_X1 U565 ( .A(n575), .B(n564), .ZN(n352) );
  XNOR2_X1 U566 ( .A(n155), .B(n558), .ZN(n139) );
  XNOR2_X1 U567 ( .A(n153), .B(n141), .ZN(n558) );
  XNOR2_X1 U568 ( .A(n157), .B(n559), .ZN(n141) );
  XNOR2_X1 U569 ( .A(n145), .B(n143), .ZN(n559) );
  OAI22_X1 U570 ( .A1(n42), .A2(n582), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U571 ( .A1(n564), .A2(n582), .ZN(n332) );
  XNOR2_X1 U572 ( .A(n577), .B(n564), .ZN(n343) );
  XNOR2_X1 U573 ( .A(n159), .B(n560), .ZN(n142) );
  XNOR2_X1 U574 ( .A(n315), .B(n261), .ZN(n560) );
  XNOR2_X1 U575 ( .A(n572), .B(n564), .ZN(n376) );
  INV_X1 U576 ( .A(n37), .ZN(n237) );
  XNOR2_X1 U577 ( .A(n579), .B(n564), .ZN(n336) );
  AND2_X1 U578 ( .A1(n565), .A2(n497), .ZN(n278) );
  OAI22_X1 U579 ( .A1(n39), .A2(n336), .B1(n37), .B2(n335), .ZN(n263) );
  AND2_X1 U580 ( .A1(n565), .A2(n237), .ZN(n264) );
  INV_X1 U581 ( .A(n19), .ZN(n574) );
  INV_X1 U582 ( .A(n25), .ZN(n576) );
  AND2_X1 U583 ( .A1(n565), .A2(n235), .ZN(n260) );
  OAI22_X1 U584 ( .A1(n39), .A2(n335), .B1(n37), .B2(n334), .ZN(n262) );
  INV_X1 U585 ( .A(n7), .ZN(n570) );
  INV_X1 U586 ( .A(n13), .ZN(n573) );
  INV_X1 U587 ( .A(n41), .ZN(n235) );
  XNOR2_X1 U588 ( .A(n522), .B(n564), .ZN(n363) );
  OAI22_X1 U589 ( .A1(n39), .A2(n580), .B1(n337), .B2(n37), .ZN(n252) );
  OR2_X1 U590 ( .A1(n564), .A2(n580), .ZN(n337) );
  AND2_X1 U591 ( .A1(n565), .A2(n247), .ZN(n314) );
  AND2_X1 U592 ( .A1(n565), .A2(n249), .ZN(product[0]) );
  OR2_X1 U593 ( .A1(n564), .A2(n574), .ZN(n364) );
  OR2_X1 U594 ( .A1(n564), .A2(n578), .ZN(n344) );
  OR2_X1 U595 ( .A1(n564), .A2(n576), .ZN(n353) );
  OR2_X1 U596 ( .A1(n564), .A2(n573), .ZN(n377) );
  XNOR2_X1 U597 ( .A(n579), .B(a[14]), .ZN(n41) );
  OAI22_X1 U598 ( .A1(n39), .A2(n334), .B1(n37), .B2(n333), .ZN(n261) );
  XNOR2_X1 U599 ( .A(n579), .B(n422), .ZN(n333) );
  XNOR2_X1 U600 ( .A(n522), .B(b[9]), .ZN(n354) );
  XNOR2_X1 U601 ( .A(n572), .B(b[11]), .ZN(n365) );
  OAI22_X1 U602 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U603 ( .A(n581), .B(n424), .ZN(n330) );
  XNOR2_X1 U604 ( .A(n581), .B(n564), .ZN(n331) );
  XNOR2_X1 U605 ( .A(n579), .B(n424), .ZN(n335) );
  XNOR2_X1 U606 ( .A(n579), .B(n423), .ZN(n334) );
  XNOR2_X1 U607 ( .A(n575), .B(n418), .ZN(n345) );
  XNOR2_X1 U608 ( .A(n577), .B(n420), .ZN(n338) );
  XNOR2_X1 U609 ( .A(n569), .B(b[13]), .ZN(n378) );
  NAND2_X1 U610 ( .A1(n427), .A2(n37), .ZN(n39) );
  XNOR2_X1 U611 ( .A(n522), .B(n424), .ZN(n362) );
  XNOR2_X1 U612 ( .A(n577), .B(n424), .ZN(n342) );
  XNOR2_X1 U613 ( .A(n575), .B(n424), .ZN(n351) );
  XNOR2_X1 U614 ( .A(n568), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U615 ( .A(n568), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U616 ( .A(n568), .B(n418), .ZN(n384) );
  XNOR2_X1 U617 ( .A(n569), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U618 ( .A(n569), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U619 ( .A(n569), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U620 ( .A(n569), .B(n419), .ZN(n385) );
  XNOR2_X1 U621 ( .A(n577), .B(n423), .ZN(n341) );
  XNOR2_X1 U622 ( .A(n577), .B(n422), .ZN(n340) );
  XNOR2_X1 U623 ( .A(n577), .B(n421), .ZN(n339) );
  XNOR2_X1 U624 ( .A(n572), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U625 ( .A(n572), .B(n418), .ZN(n369) );
  XNOR2_X1 U626 ( .A(n572), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U627 ( .A(n572), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U628 ( .A(n522), .B(n423), .ZN(n361) );
  XNOR2_X1 U629 ( .A(n522), .B(n422), .ZN(n360) );
  XNOR2_X1 U630 ( .A(n575), .B(n422), .ZN(n349) );
  XNOR2_X1 U631 ( .A(n575), .B(n423), .ZN(n350) );
  XNOR2_X1 U632 ( .A(n520), .B(b[11]), .ZN(n397) );
  XNOR2_X1 U633 ( .A(n519), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U634 ( .A(n519), .B(b[13]), .ZN(n395) );
  XNOR2_X1 U635 ( .A(n520), .B(b[14]), .ZN(n394) );
  XNOR2_X1 U636 ( .A(n522), .B(n421), .ZN(n359) );
  XNOR2_X1 U637 ( .A(n522), .B(n420), .ZN(n358) );
  XNOR2_X1 U638 ( .A(n575), .B(n421), .ZN(n348) );
  XNOR2_X1 U639 ( .A(n575), .B(n420), .ZN(n347) );
  XNOR2_X1 U640 ( .A(n522), .B(n418), .ZN(n356) );
  XNOR2_X1 U641 ( .A(n522), .B(n419), .ZN(n357) );
  XNOR2_X1 U642 ( .A(n575), .B(n419), .ZN(n346) );
  XNOR2_X1 U643 ( .A(n522), .B(b[8]), .ZN(n355) );
  NAND2_X1 U644 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U645 ( .A(n581), .B(a[14]), .Z(n426) );
  XNOR2_X1 U646 ( .A(n519), .B(b[15]), .ZN(n393) );
  BUF_X1 U647 ( .A(n43), .Z(n565) );
  XOR2_X1 U648 ( .A(n579), .B(a[12]), .Z(n427) );
  NAND2_X1 U649 ( .A1(n328), .A2(n314), .ZN(n119) );
  INV_X1 U650 ( .A(n249), .ZN(n563) );
  INV_X1 U651 ( .A(n113), .ZN(n135) );
  NOR2_X1 U652 ( .A1(n234), .A2(n257), .ZN(n113) );
  INV_X1 U653 ( .A(n517), .ZN(n127) );
  NOR2_X1 U654 ( .A1(n517), .A2(n85), .ZN(n80) );
  OAI21_X1 U655 ( .B1(n82), .B2(n86), .A(n83), .ZN(n81) );
  NAND2_X1 U656 ( .A1(n186), .A2(n195), .ZN(n83) );
  OAI22_X1 U657 ( .A1(n34), .A2(n339), .B1(n338), .B2(n32), .ZN(n265) );
  OAI22_X1 U658 ( .A1(n34), .A2(n340), .B1(n339), .B2(n32), .ZN(n266) );
  OAI22_X1 U659 ( .A1(n34), .A2(n342), .B1(n341), .B2(n32), .ZN(n268) );
  OAI22_X1 U660 ( .A1(n34), .A2(n341), .B1(n340), .B2(n32), .ZN(n267) );
  OAI22_X1 U661 ( .A1(n34), .A2(n343), .B1(n342), .B2(n32), .ZN(n269) );
  OAI22_X1 U662 ( .A1(n34), .A2(n578), .B1(n344), .B2(n32), .ZN(n253) );
  NAND2_X1 U663 ( .A1(n556), .A2(n103), .ZN(n55) );
  NAND2_X1 U664 ( .A1(n232), .A2(n233), .ZN(n111) );
  INV_X1 U665 ( .A(n111), .ZN(n109) );
  NAND2_X1 U666 ( .A1(n555), .A2(n111), .ZN(n57) );
  XNOR2_X1 U667 ( .A(n84), .B(n50), .ZN(product[11]) );
  XNOR2_X1 U668 ( .A(n571), .B(n424), .ZN(n375) );
  XNOR2_X1 U669 ( .A(n571), .B(n423), .ZN(n374) );
  XNOR2_X1 U670 ( .A(n571), .B(n422), .ZN(n373) );
  XNOR2_X1 U671 ( .A(n571), .B(n419), .ZN(n370) );
  XNOR2_X1 U672 ( .A(n571), .B(n420), .ZN(n371) );
  XNOR2_X1 U673 ( .A(n571), .B(n421), .ZN(n372) );
  NOR2_X1 U674 ( .A1(n204), .A2(n211), .ZN(n89) );
  OAI22_X1 U675 ( .A1(n29), .A2(n346), .B1(n345), .B2(n27), .ZN(n271) );
  OAI22_X1 U676 ( .A1(n29), .A2(n350), .B1(n349), .B2(n27), .ZN(n275) );
  OAI22_X1 U677 ( .A1(n29), .A2(n347), .B1(n346), .B2(n27), .ZN(n272) );
  OAI22_X1 U678 ( .A1(n29), .A2(n349), .B1(n348), .B2(n27), .ZN(n274) );
  OAI22_X1 U679 ( .A1(n29), .A2(n576), .B1(n353), .B2(n27), .ZN(n254) );
  OAI22_X1 U680 ( .A1(n29), .A2(n348), .B1(n347), .B2(n27), .ZN(n273) );
  OAI22_X1 U681 ( .A1(n29), .A2(n351), .B1(n350), .B2(n27), .ZN(n276) );
  OAI22_X1 U682 ( .A1(n29), .A2(n352), .B1(n351), .B2(n27), .ZN(n277) );
  INV_X1 U683 ( .A(n1), .ZN(n567) );
  OR2_X1 U684 ( .A1(n564), .A2(n511), .ZN(n409) );
  OAI21_X1 U685 ( .B1(n491), .B2(n97), .A(n98), .ZN(n96) );
  XNOR2_X1 U686 ( .A(n507), .B(n55), .ZN(product[6]) );
  AOI21_X1 U687 ( .B1(n556), .B2(n104), .A(n521), .ZN(n99) );
  OAI22_X1 U688 ( .A1(n6), .A2(n394), .B1(n393), .B2(n539), .ZN(n315) );
  OAI22_X1 U689 ( .A1(n547), .A2(n395), .B1(n394), .B2(n538), .ZN(n316) );
  NAND2_X1 U690 ( .A1(n329), .A2(n258), .ZN(n122) );
  OAI22_X1 U691 ( .A1(n6), .A2(n397), .B1(n396), .B2(n539), .ZN(n318) );
  OAI22_X1 U692 ( .A1(n547), .A2(n401), .B1(n400), .B2(n539), .ZN(n322) );
  OAI22_X1 U693 ( .A1(n546), .A2(n398), .B1(n397), .B2(n538), .ZN(n319) );
  OAI22_X1 U694 ( .A1(n546), .A2(n396), .B1(n395), .B2(n539), .ZN(n317) );
  OAI22_X1 U695 ( .A1(n547), .A2(n399), .B1(n398), .B2(n539), .ZN(n320) );
  OAI22_X1 U696 ( .A1(n6), .A2(n400), .B1(n399), .B2(n538), .ZN(n321) );
  OAI22_X1 U697 ( .A1(n6), .A2(n402), .B1(n401), .B2(n538), .ZN(n323) );
  OAI22_X1 U698 ( .A1(n547), .A2(n404), .B1(n403), .B2(n539), .ZN(n325) );
  OAI22_X1 U699 ( .A1(n403), .A2(n6), .B1(n402), .B2(n538), .ZN(n324) );
  OAI22_X1 U700 ( .A1(n546), .A2(n406), .B1(n405), .B2(n539), .ZN(n327) );
  OAI22_X1 U701 ( .A1(n546), .A2(n405), .B1(n404), .B2(n538), .ZN(n326) );
  OAI22_X1 U702 ( .A1(n546), .A2(n407), .B1(n406), .B2(n538), .ZN(n328) );
  OAI22_X1 U703 ( .A1(n547), .A2(n408), .B1(n407), .B2(n538), .ZN(n329) );
  OAI22_X1 U704 ( .A1(n6), .A2(n511), .B1(n409), .B2(n539), .ZN(n258) );
  OAI22_X1 U705 ( .A1(n23), .A2(n358), .B1(n357), .B2(n21), .ZN(n282) );
  OAI22_X1 U706 ( .A1(n23), .A2(n356), .B1(n355), .B2(n21), .ZN(n280) );
  OAI22_X1 U707 ( .A1(n23), .A2(n360), .B1(n359), .B2(n21), .ZN(n284) );
  OAI22_X1 U708 ( .A1(n23), .A2(n362), .B1(n361), .B2(n21), .ZN(n286) );
  OAI22_X1 U709 ( .A1(n23), .A2(n355), .B1(n354), .B2(n21), .ZN(n279) );
  OAI22_X1 U710 ( .A1(n23), .A2(n361), .B1(n360), .B2(n21), .ZN(n285) );
  OAI22_X1 U711 ( .A1(n23), .A2(n574), .B1(n364), .B2(n21), .ZN(n255) );
  OAI22_X1 U712 ( .A1(n23), .A2(n357), .B1(n356), .B2(n21), .ZN(n281) );
  OAI22_X1 U713 ( .A1(n23), .A2(n363), .B1(n362), .B2(n21), .ZN(n287) );
  XNOR2_X1 U714 ( .A(n77), .B(n48), .ZN(product[13]) );
  XOR2_X1 U715 ( .A(n56), .B(n512), .Z(product[5]) );
  XNOR2_X1 U716 ( .A(n70), .B(n47), .ZN(product[14]) );
  XNOR2_X1 U717 ( .A(n57), .B(n112), .ZN(product[4]) );
  OAI21_X1 U718 ( .B1(n87), .B2(n85), .A(n86), .ZN(n84) );
  NAND2_X1 U719 ( .A1(n151), .A2(n139), .ZN(n62) );
  OAI22_X1 U720 ( .A1(n505), .A2(n375), .B1(n374), .B2(n561), .ZN(n298) );
  OAI22_X1 U721 ( .A1(n505), .A2(n370), .B1(n369), .B2(n561), .ZN(n293) );
  OAI22_X1 U722 ( .A1(n505), .A2(n373), .B1(n372), .B2(n561), .ZN(n296) );
  OAI22_X1 U723 ( .A1(n505), .A2(n367), .B1(n366), .B2(n561), .ZN(n290) );
  OAI22_X1 U724 ( .A1(n504), .A2(n372), .B1(n371), .B2(n561), .ZN(n295) );
  OAI22_X1 U725 ( .A1(n505), .A2(n374), .B1(n373), .B2(n561), .ZN(n297) );
  OAI22_X1 U726 ( .A1(n505), .A2(n376), .B1(n375), .B2(n561), .ZN(n299) );
  OAI22_X1 U727 ( .A1(n505), .A2(n573), .B1(n377), .B2(n561), .ZN(n256) );
  OAI22_X1 U728 ( .A1(n505), .A2(n371), .B1(n370), .B2(n561), .ZN(n294) );
  OAI22_X1 U729 ( .A1(n505), .A2(n368), .B1(n367), .B2(n561), .ZN(n291) );
  OAI22_X1 U730 ( .A1(n504), .A2(n369), .B1(n368), .B2(n561), .ZN(n292) );
  XNOR2_X1 U731 ( .A(n569), .B(n420), .ZN(n386) );
  OAI22_X1 U732 ( .A1(n504), .A2(n366), .B1(n365), .B2(n561), .ZN(n289) );
  INV_X1 U733 ( .A(n561), .ZN(n245) );
  XNOR2_X1 U734 ( .A(n568), .B(n422), .ZN(n388) );
  XNOR2_X1 U735 ( .A(n568), .B(n421), .ZN(n387) );
  XNOR2_X1 U736 ( .A(n569), .B(n564), .ZN(n391) );
  XNOR2_X1 U737 ( .A(n569), .B(n423), .ZN(n389) );
  XNOR2_X1 U738 ( .A(n569), .B(n424), .ZN(n390) );
  INV_X1 U739 ( .A(n526), .ZN(n87) );
  AOI21_X1 U740 ( .B1(n494), .B2(n552), .A(n93), .ZN(n91) );
  AND2_X1 U741 ( .A1(n565), .A2(n245), .ZN(n300) );
  NAND2_X1 U742 ( .A1(n135), .A2(n114), .ZN(n58) );
  OAI21_X1 U743 ( .B1(n534), .B2(n78), .A(n79), .ZN(n77) );
  OAI21_X1 U744 ( .B1(n45), .B2(n71), .A(n72), .ZN(n70) );
  OAI21_X1 U745 ( .B1(n64), .B2(n536), .A(n65), .ZN(n63) );
  XNOR2_X1 U746 ( .A(n535), .B(n53), .ZN(product[8]) );
  XNOR2_X1 U747 ( .A(n520), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U748 ( .A(n520), .B(n418), .ZN(n401) );
  XNOR2_X1 U749 ( .A(n518), .B(n420), .ZN(n403) );
  XNOR2_X1 U750 ( .A(n518), .B(n421), .ZN(n404) );
  XNOR2_X1 U751 ( .A(n518), .B(n422), .ZN(n405) );
  XNOR2_X1 U752 ( .A(n520), .B(n564), .ZN(n408) );
  XNOR2_X1 U753 ( .A(n519), .B(n423), .ZN(n406) );
  XNOR2_X1 U754 ( .A(n519), .B(n424), .ZN(n407) );
  XOR2_X1 U755 ( .A(n525), .B(n54), .Z(product[7]) );
  OAI22_X1 U756 ( .A1(n545), .A2(n379), .B1(n378), .B2(n501), .ZN(n301) );
  OAI22_X1 U757 ( .A1(n508), .A2(n380), .B1(n379), .B2(n501), .ZN(n302) );
  OAI22_X1 U758 ( .A1(n545), .A2(n385), .B1(n384), .B2(n501), .ZN(n307) );
  OAI22_X1 U759 ( .A1(n508), .A2(n382), .B1(n381), .B2(n501), .ZN(n304) );
  OAI22_X1 U760 ( .A1(n508), .A2(n381), .B1(n380), .B2(n501), .ZN(n303) );
  NAND2_X1 U761 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U762 ( .A1(n544), .A2(n383), .B1(n382), .B2(n562), .ZN(n305) );
  OAI22_X1 U763 ( .A1(n545), .A2(n384), .B1(n383), .B2(n501), .ZN(n306) );
  OAI22_X1 U764 ( .A1(n545), .A2(n386), .B1(n385), .B2(n501), .ZN(n308) );
  OAI22_X1 U765 ( .A1(n545), .A2(n387), .B1(n386), .B2(n501), .ZN(n309) );
  OAI22_X1 U766 ( .A1(n508), .A2(n496), .B1(n392), .B2(n501), .ZN(n257) );
  OAI22_X1 U767 ( .A1(n508), .A2(n389), .B1(n388), .B2(n562), .ZN(n311) );
  OAI22_X1 U768 ( .A1(n544), .A2(n388), .B1(n562), .B2(n387), .ZN(n310) );
  OAI22_X1 U769 ( .A1(n508), .A2(n390), .B1(n389), .B2(n501), .ZN(n312) );
  INV_X1 U770 ( .A(n501), .ZN(n247) );
  OAI22_X1 U771 ( .A1(n545), .A2(n391), .B1(n390), .B2(n501), .ZN(n313) );
  INV_X1 U772 ( .A(n573), .ZN(n571) );
  INV_X1 U773 ( .A(n573), .ZN(n572) );
  INV_X1 U774 ( .A(n31), .ZN(n578) );
  INV_X1 U775 ( .A(n580), .ZN(n579) );
  INV_X1 U776 ( .A(n36), .ZN(n580) );
  INV_X1 U777 ( .A(n582), .ZN(n581) );
  INV_X1 U778 ( .A(n40), .ZN(n582) );
  XOR2_X1 U779 ( .A(n259), .B(n251), .Z(n148) );
  XOR2_X1 U780 ( .A(n289), .B(n279), .Z(n146) );
  XOR2_X1 U781 ( .A(n149), .B(n147), .Z(n144) );
endmodule


module layer1_8_4_8_16_datapath_M8_N4_T16_P8_6_DW01_add_2 ( A, B, CI, SUM, CO
 );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n4, n6, n8, n9, n10, n11, n12, n13, n14, n15, n18, n19, n20,
         n21, n23, n25, n26, n27, n28, n30, n34, n35, n36, n37, n38, n39, n40,
         n41, n43, n44, n48, n49, n51, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n69, n71, n72, n73, n74, n75, n77,
         n79, n80, n81, n82, n83, n85, n87, n88, n90, n93, n95, n98, n99, n100,
         n102, n104, n161, n162, n163, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185;

  XNOR2_X1 U126 ( .A(n162), .B(n161), .ZN(SUM[9]) );
  AND2_X1 U127 ( .A1(n180), .A2(n53), .ZN(n161) );
  AOI21_X1 U128 ( .B1(n56), .B2(n64), .A(n57), .ZN(n162) );
  BUF_X1 U129 ( .A(n40), .Z(n172) );
  OR2_X1 U130 ( .A1(A[12]), .A2(B[12]), .ZN(n163) );
  AND2_X1 U131 ( .A1(n179), .A2(n90), .ZN(SUM[0]) );
  OR2_X1 U132 ( .A1(A[15]), .A2(B[15]), .ZN(n165) );
  BUF_X1 U133 ( .A(n59), .Z(n166) );
  INV_X1 U134 ( .A(n170), .ZN(n48) );
  AND2_X1 U135 ( .A1(A[10]), .A2(B[10]), .ZN(n170) );
  CLKBUF_X1 U136 ( .A(n183), .Z(n167) );
  NOR2_X1 U137 ( .A1(A[12]), .A2(B[12]), .ZN(n168) );
  NOR2_X1 U138 ( .A1(A[12]), .A2(B[12]), .ZN(n36) );
  XNOR2_X1 U139 ( .A(n169), .B(n41), .ZN(SUM[11]) );
  AND2_X1 U140 ( .A1(n95), .A2(n172), .ZN(n169) );
  OR2_X2 U141 ( .A1(A[10]), .A2(B[10]), .ZN(n183) );
  XNOR2_X1 U142 ( .A(n177), .B(n171), .ZN(SUM[13]) );
  AND2_X1 U143 ( .A1(n93), .A2(n28), .ZN(n171) );
  INV_X1 U144 ( .A(n95), .ZN(n173) );
  NOR2_X1 U145 ( .A1(A[8]), .A2(B[8]), .ZN(n174) );
  OAI21_X1 U146 ( .B1(n43), .B2(n55), .A(n44), .ZN(n175) );
  OAI21_X1 U147 ( .B1(n36), .B2(n40), .A(n37), .ZN(n176) );
  AOI21_X1 U148 ( .B1(n175), .B2(n34), .A(n176), .ZN(n177) );
  AOI21_X1 U149 ( .B1(n175), .B2(n34), .A(n35), .ZN(n178) );
  OR2_X1 U150 ( .A1(A[0]), .A2(B[0]), .ZN(n179) );
  INV_X1 U151 ( .A(n162), .ZN(n54) );
  AOI21_X1 U152 ( .B1(n181), .B2(n80), .A(n77), .ZN(n75) );
  INV_X1 U153 ( .A(n79), .ZN(n77) );
  AOI21_X1 U154 ( .B1(n182), .B2(n88), .A(n85), .ZN(n83) );
  INV_X1 U155 ( .A(n87), .ZN(n85) );
  AOI21_X1 U156 ( .B1(n56), .B2(n64), .A(n57), .ZN(n55) );
  OAI21_X1 U157 ( .B1(n83), .B2(n81), .A(n82), .ZN(n80) );
  AOI21_X1 U158 ( .B1(n184), .B2(n72), .A(n69), .ZN(n67) );
  INV_X1 U159 ( .A(n71), .ZN(n69) );
  INV_X1 U160 ( .A(n28), .ZN(n30) );
  OAI21_X1 U161 ( .B1(n75), .B2(n73), .A(n74), .ZN(n72) );
  AOI21_X1 U162 ( .B1(n54), .B2(n180), .A(n51), .ZN(n49) );
  NAND2_X1 U163 ( .A1(n98), .A2(n166), .ZN(n8) );
  INV_X1 U164 ( .A(n90), .ZN(n88) );
  OAI21_X1 U165 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  INV_X1 U166 ( .A(n53), .ZN(n51) );
  INV_X1 U167 ( .A(n27), .ZN(n93) );
  NAND2_X1 U168 ( .A1(n102), .A2(n74), .ZN(n12) );
  INV_X1 U169 ( .A(n73), .ZN(n102) );
  INV_X1 U170 ( .A(n39), .ZN(n95) );
  NAND2_X1 U171 ( .A1(n99), .A2(n62), .ZN(n9) );
  INV_X1 U172 ( .A(n61), .ZN(n99) );
  NAND2_X1 U173 ( .A1(n104), .A2(n82), .ZN(n14) );
  INV_X1 U174 ( .A(n81), .ZN(n104) );
  NAND2_X1 U175 ( .A1(n184), .A2(n71), .ZN(n11) );
  NAND2_X1 U176 ( .A1(n181), .A2(n79), .ZN(n13) );
  NAND2_X1 U177 ( .A1(n182), .A2(n87), .ZN(n15) );
  NAND2_X1 U178 ( .A1(n100), .A2(n66), .ZN(n10) );
  INV_X1 U179 ( .A(n65), .ZN(n100) );
  INV_X1 U180 ( .A(n25), .ZN(n23) );
  XNOR2_X1 U181 ( .A(n38), .B(n4), .ZN(SUM[12]) );
  NAND2_X1 U182 ( .A1(n163), .A2(n37), .ZN(n4) );
  XOR2_X1 U183 ( .A(n12), .B(n75), .Z(SUM[4]) );
  XNOR2_X1 U184 ( .A(n13), .B(n80), .ZN(SUM[3]) );
  XNOR2_X1 U185 ( .A(n15), .B(n88), .ZN(SUM[1]) );
  NOR2_X1 U186 ( .A1(A[7]), .A2(B[7]), .ZN(n61) );
  OR2_X1 U187 ( .A1(A[9]), .A2(B[9]), .ZN(n180) );
  NOR2_X1 U188 ( .A1(A[2]), .A2(B[2]), .ZN(n81) );
  NOR2_X1 U189 ( .A1(A[4]), .A2(B[4]), .ZN(n73) );
  NAND2_X1 U190 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  XOR2_X1 U191 ( .A(n49), .B(n6), .Z(SUM[10]) );
  XOR2_X1 U192 ( .A(n63), .B(n9), .Z(SUM[7]) );
  NAND2_X1 U193 ( .A1(A[11]), .A2(B[11]), .ZN(n40) );
  OR2_X1 U194 ( .A1(A[3]), .A2(B[3]), .ZN(n181) );
  OR2_X1 U195 ( .A1(A[1]), .A2(B[1]), .ZN(n182) );
  NOR2_X1 U196 ( .A1(A[11]), .A2(B[11]), .ZN(n39) );
  NOR2_X1 U197 ( .A1(A[8]), .A2(B[8]), .ZN(n58) );
  XNOR2_X1 U198 ( .A(n60), .B(n8), .ZN(SUM[8]) );
  NOR2_X1 U199 ( .A1(A[6]), .A2(B[6]), .ZN(n65) );
  NAND2_X1 U200 ( .A1(A[7]), .A2(B[7]), .ZN(n62) );
  OR2_X1 U201 ( .A1(A[5]), .A2(B[5]), .ZN(n184) );
  NAND2_X1 U202 ( .A1(A[2]), .A2(B[2]), .ZN(n82) );
  NAND2_X1 U203 ( .A1(A[4]), .A2(B[4]), .ZN(n74) );
  NAND2_X1 U204 ( .A1(A[9]), .A2(B[9]), .ZN(n53) );
  NAND2_X1 U205 ( .A1(A[1]), .A2(B[1]), .ZN(n87) );
  NAND2_X1 U206 ( .A1(A[5]), .A2(B[5]), .ZN(n71) );
  NAND2_X1 U207 ( .A1(A[3]), .A2(B[3]), .ZN(n79) );
  NAND2_X1 U208 ( .A1(A[0]), .A2(B[0]), .ZN(n90) );
  NAND2_X1 U209 ( .A1(A[8]), .A2(B[8]), .ZN(n59) );
  NAND2_X1 U210 ( .A1(A[6]), .A2(B[6]), .ZN(n66) );
  NAND2_X1 U211 ( .A1(A[12]), .A2(B[12]), .ZN(n37) );
  XNOR2_X1 U212 ( .A(n11), .B(n72), .ZN(SUM[5]) );
  XOR2_X1 U213 ( .A(n14), .B(n83), .Z(SUM[2]) );
  NAND2_X1 U214 ( .A1(n165), .A2(n18), .ZN(n1) );
  OR2_X1 U215 ( .A1(A[14]), .A2(B[14]), .ZN(n185) );
  NAND2_X1 U216 ( .A1(A[14]), .A2(B[14]), .ZN(n25) );
  AOI21_X1 U217 ( .B1(n183), .B2(n51), .A(n170), .ZN(n44) );
  INV_X1 U218 ( .A(n174), .ZN(n98) );
  NOR2_X1 U219 ( .A1(n174), .A2(n61), .ZN(n56) );
  OAI21_X1 U220 ( .B1(n58), .B2(n62), .A(n59), .ZN(n57) );
  XNOR2_X1 U221 ( .A(n19), .B(n1), .ZN(SUM[15]) );
  INV_X1 U222 ( .A(n64), .ZN(n63) );
  OAI21_X1 U223 ( .B1(n67), .B2(n65), .A(n66), .ZN(n64) );
  XOR2_X1 U224 ( .A(n10), .B(n67), .Z(SUM[6]) );
  NAND2_X1 U225 ( .A1(n185), .A2(n25), .ZN(n2) );
  NAND2_X1 U226 ( .A1(n185), .A2(n93), .ZN(n20) );
  NOR2_X1 U227 ( .A1(A[13]), .A2(B[13]), .ZN(n27) );
  AOI21_X1 U228 ( .B1(n185), .B2(n30), .A(n23), .ZN(n21) );
  NAND2_X1 U229 ( .A1(A[15]), .A2(B[15]), .ZN(n18) );
  OAI21_X1 U230 ( .B1(n41), .B2(n173), .A(n172), .ZN(n38) );
  INV_X1 U231 ( .A(n175), .ZN(n41) );
  NOR2_X1 U232 ( .A1(n168), .A2(n39), .ZN(n34) );
  OAI21_X1 U233 ( .B1(n168), .B2(n40), .A(n37), .ZN(n35) );
  NAND2_X1 U234 ( .A1(n167), .A2(n48), .ZN(n6) );
  NAND2_X1 U235 ( .A1(n183), .A2(n180), .ZN(n43) );
  XNOR2_X1 U236 ( .A(n26), .B(n2), .ZN(SUM[14]) );
  OAI21_X1 U237 ( .B1(n177), .B2(n27), .A(n28), .ZN(n26) );
  OAI21_X1 U238 ( .B1(n178), .B2(n20), .A(n21), .ZN(n19) );
endmodule


module layer1_8_4_8_16_datapath_M8_N4_T16_P8_6 ( clk, clear_acc, data_out_x, 
        data_out, data_out_w, data_out_b, wr_en_y, m_valid, m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [3:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N27, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, n1, n2, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n87, n104, n113, n114, n115, n116, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n22), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n229), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n230), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n231), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n232), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n233), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n234), .CK(clk), .Q(n34) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n235), .CK(clk), .Q(n35) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n236), .CK(clk), .Q(n36) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n237), .CK(clk), .Q(n37) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n238), .CK(clk), .Q(n38) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n239), .CK(clk), .Q(n39) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n240), .CK(clk), .Q(n40) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n241), .CK(clk), .Q(n41) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n242), .CK(clk), .Q(n42) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n243), .CK(clk), .Q(n43) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n244), .CK(clk), .Q(n45) );
  DFF_X1 \f_reg[0]  ( .D(n168), .CK(clk), .Q(n66), .QN(n218) );
  DFF_X1 \f_reg[1]  ( .D(n116), .CK(clk), .Q(n64), .QN(n219) );
  DFF_X1 \f_reg[2]  ( .D(n115), .CK(clk), .Q(n62), .QN(n220) );
  DFF_X1 \f_reg[3]  ( .D(n114), .CK(clk), .Q(f[3]), .QN(n70) );
  DFF_X1 \f_reg[4]  ( .D(n113), .CK(clk), .Q(f[4]), .QN(n71) );
  DFF_X1 \f_reg[5]  ( .D(n104), .CK(clk), .Q(f[5]), .QN(n72) );
  DFF_X1 \f_reg[6]  ( .D(n87), .CK(clk), .Q(f[6]), .QN(n73) );
  DFF_X1 \f_reg[7]  ( .D(n85), .CK(clk), .Q(f[7]), .QN(n221) );
  DFF_X1 \f_reg[8]  ( .D(n84), .CK(clk), .Q(f[8]), .QN(n222) );
  DFF_X1 \f_reg[9]  ( .D(n83), .CK(clk), .Q(f[9]), .QN(n223) );
  DFF_X1 \f_reg[10]  ( .D(n82), .CK(clk), .Q(n54), .QN(n224) );
  DFF_X1 \f_reg[11]  ( .D(n81), .CK(clk), .Q(n52), .QN(n225) );
  DFF_X1 \f_reg[12]  ( .D(n7), .CK(clk), .Q(n51), .QN(n226) );
  DFF_X1 \f_reg[13]  ( .D(n2), .CK(clk), .Q(n50), .QN(n227) );
  DFF_X1 \f_reg[14]  ( .D(n80), .CK(clk), .Q(n49), .QN(n228) );
  DFF_X1 \f_reg[15]  ( .D(n8), .CK(clk), .Q(f[15]), .QN(n78) );
  DFF_X1 \data_out_reg[15]  ( .D(n170), .CK(clk), .Q(data_out[15]), .QN(n201)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n171), .CK(clk), .Q(data_out[14]), .QN(n200)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n172), .CK(clk), .Q(data_out[13]), .QN(n199)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n173), .CK(clk), .Q(data_out[12]), .QN(n198)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n174), .CK(clk), .Q(data_out[11]), .QN(n197)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n175), .CK(clk), .Q(data_out[10]), .QN(n196)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n176), .CK(clk), .Q(data_out[9]), .QN(n195) );
  DFF_X1 \data_out_reg[8]  ( .D(n177), .CK(clk), .Q(data_out[8]), .QN(n194) );
  DFF_X1 \data_out_reg[7]  ( .D(n178), .CK(clk), .Q(data_out[7]), .QN(n193) );
  DFF_X1 \data_out_reg[6]  ( .D(n179), .CK(clk), .Q(data_out[6]), .QN(n192) );
  DFF_X1 \data_out_reg[5]  ( .D(n180), .CK(clk), .Q(data_out[5]), .QN(n191) );
  DFF_X1 \data_out_reg[4]  ( .D(n181), .CK(clk), .Q(data_out[4]), .QN(n190) );
  DFF_X1 \data_out_reg[3]  ( .D(n182), .CK(clk), .Q(data_out[3]), .QN(n189) );
  DFF_X1 \data_out_reg[2]  ( .D(n183), .CK(clk), .Q(data_out[2]), .QN(n188) );
  DFF_X1 \data_out_reg[1]  ( .D(n184), .CK(clk), .Q(data_out[1]), .QN(n187) );
  DFF_X1 \data_out_reg[0]  ( .D(n185), .CK(clk), .Q(data_out[0]), .QN(n186) );
  layer1_8_4_8_16_datapath_M8_N4_T16_P8_6_DW_mult_tc_1 mult_183 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer1_8_4_8_16_datapath_M8_N4_T16_P8_6_DW01_add_2 add_184 ( .A({n208, n207, 
        n206, n205, n204, n203, n217, n216, n215, n214, n213, n212, n211, n210, 
        n209, n202}), .B({f[15], n49, n50, n51, n52, n54, f[9:3], n62, n64, 
        n66}), .CI(1'b0), .SUM(adder) );
  DFF_X2 delay_reg ( .D(N27), .CK(clk), .Q(n13), .QN(n245) );
  CLKBUF_X1 U3 ( .A(N40), .Z(n1) );
  NAND3_X1 U4 ( .A1(n5), .A2(n4), .A3(n6), .ZN(n2) );
  NAND2_X1 U5 ( .A1(data_out_b[13]), .A2(n22), .ZN(n4) );
  NAND2_X1 U6 ( .A1(adder[13]), .A2(n21), .ZN(n5) );
  NAND2_X1 U8 ( .A1(n68), .A2(n50), .ZN(n6) );
  MUX2_X2 U9 ( .A(N42), .B(n29), .S(n13), .Z(n206) );
  NAND3_X1 U10 ( .A1(n10), .A2(n9), .A3(n11), .ZN(n7) );
  NAND3_X1 U11 ( .A1(n16), .A2(n15), .A3(n17), .ZN(n8) );
  MUX2_X2 U12 ( .A(n36), .B(N37), .S(n245), .Z(n216) );
  NAND2_X1 U13 ( .A1(data_out_b[12]), .A2(n22), .ZN(n9) );
  NAND2_X1 U14 ( .A1(adder[12]), .A2(n21), .ZN(n10) );
  NAND2_X1 U15 ( .A1(n68), .A2(n51), .ZN(n11) );
  CLKBUF_X1 U16 ( .A(N39), .Z(n12) );
  MUX2_X2 U17 ( .A(N39), .B(n34), .S(n13), .Z(n203) );
  AND2_X1 U18 ( .A1(n20), .A2(n18), .ZN(n14) );
  NAND2_X1 U19 ( .A1(n19), .A2(n14), .ZN(n80) );
  MUX2_X2 U20 ( .A(n32), .B(N41), .S(n245), .Z(n205) );
  NAND2_X1 U21 ( .A1(data_out_b[15]), .A2(n22), .ZN(n15) );
  NAND2_X1 U22 ( .A1(adder[15]), .A2(n21), .ZN(n16) );
  NAND2_X1 U23 ( .A1(n68), .A2(f[15]), .ZN(n17) );
  NAND2_X1 U24 ( .A1(data_out_b[14]), .A2(n22), .ZN(n18) );
  NAND2_X1 U25 ( .A1(adder[14]), .A2(n21), .ZN(n19) );
  NAND2_X1 U26 ( .A1(n68), .A2(n49), .ZN(n20) );
  AND2_X2 U27 ( .A1(n48), .A2(n23), .ZN(n21) );
  INV_X1 U28 ( .A(n23), .ZN(n22) );
  INV_X1 U29 ( .A(n48), .ZN(n68) );
  INV_X1 U30 ( .A(clear_acc), .ZN(n23) );
  NAND2_X1 U31 ( .A1(n169), .A2(N27), .ZN(n247) );
  INV_X1 U32 ( .A(wr_en_y), .ZN(n169) );
  OAI22_X1 U33 ( .A1(n189), .A2(n247), .B1(n70), .B2(n246), .ZN(n182) );
  OAI22_X1 U34 ( .A1(n190), .A2(n247), .B1(n71), .B2(n246), .ZN(n181) );
  OAI22_X1 U35 ( .A1(n191), .A2(n247), .B1(n72), .B2(n246), .ZN(n180) );
  OAI22_X1 U36 ( .A1(n192), .A2(n247), .B1(n73), .B2(n246), .ZN(n179) );
  OAI22_X1 U37 ( .A1(n193), .A2(n247), .B1(n221), .B2(n246), .ZN(n178) );
  OAI22_X1 U38 ( .A1(n194), .A2(n247), .B1(n222), .B2(n246), .ZN(n177) );
  OAI22_X1 U39 ( .A1(n195), .A2(n247), .B1(n223), .B2(n246), .ZN(n176) );
  INV_X1 U40 ( .A(n26), .ZN(n44) );
  MUX2_X1 U41 ( .A(n33), .B(N40), .S(n245), .Z(n204) );
  MUX2_X1 U42 ( .A(n27), .B(N44), .S(n245), .Z(n208) );
  MUX2_X1 U43 ( .A(n28), .B(N43), .S(n245), .Z(n207) );
  AND3_X1 U44 ( .A1(sel[1]), .A2(sel[2]), .A3(sel[0]), .ZN(n25) );
  INV_X1 U45 ( .A(m_ready), .ZN(n24) );
  NAND2_X1 U46 ( .A1(m_valid), .A2(n24), .ZN(n46) );
  OAI21_X1 U47 ( .B1(sel[3]), .B2(n25), .A(n46), .ZN(N27) );
  NAND2_X1 U48 ( .A1(clear_acc_delay), .A2(n245), .ZN(n26) );
  MUX2_X1 U49 ( .A(n27), .B(N44), .S(n44), .Z(n229) );
  MUX2_X1 U50 ( .A(n28), .B(N43), .S(n44), .Z(n230) );
  MUX2_X1 U51 ( .A(n29), .B(N42), .S(n44), .Z(n231) );
  MUX2_X1 U52 ( .A(n32), .B(N41), .S(n44), .Z(n232) );
  MUX2_X1 U53 ( .A(n33), .B(n1), .S(n44), .Z(n233) );
  MUX2_X1 U54 ( .A(n34), .B(n12), .S(n44), .Z(n234) );
  MUX2_X1 U55 ( .A(n35), .B(N38), .S(n44), .Z(n235) );
  MUX2_X1 U56 ( .A(n35), .B(N38), .S(n245), .Z(n217) );
  MUX2_X1 U57 ( .A(n36), .B(N37), .S(n44), .Z(n236) );
  MUX2_X1 U58 ( .A(n37), .B(N36), .S(n44), .Z(n237) );
  MUX2_X1 U59 ( .A(n37), .B(N36), .S(n245), .Z(n215) );
  MUX2_X1 U60 ( .A(n38), .B(N35), .S(n44), .Z(n238) );
  MUX2_X1 U61 ( .A(n38), .B(N35), .S(n245), .Z(n214) );
  MUX2_X1 U62 ( .A(n39), .B(N34), .S(n44), .Z(n239) );
  MUX2_X1 U63 ( .A(n39), .B(N34), .S(n245), .Z(n213) );
  MUX2_X1 U64 ( .A(n40), .B(N33), .S(n44), .Z(n240) );
  MUX2_X1 U65 ( .A(n40), .B(N33), .S(n245), .Z(n212) );
  MUX2_X1 U66 ( .A(n41), .B(N32), .S(n44), .Z(n241) );
  MUX2_X1 U67 ( .A(n41), .B(N32), .S(n245), .Z(n211) );
  MUX2_X1 U68 ( .A(n42), .B(N31), .S(n44), .Z(n242) );
  MUX2_X1 U69 ( .A(n42), .B(N31), .S(n245), .Z(n210) );
  MUX2_X1 U70 ( .A(n43), .B(N30), .S(n44), .Z(n243) );
  MUX2_X1 U71 ( .A(n43), .B(N30), .S(n245), .Z(n209) );
  MUX2_X1 U72 ( .A(n45), .B(N29), .S(n44), .Z(n244) );
  MUX2_X1 U73 ( .A(n45), .B(N29), .S(n245), .Z(n202) );
  INV_X1 U74 ( .A(n46), .ZN(n47) );
  OAI21_X1 U75 ( .B1(n47), .B2(n13), .A(n23), .ZN(n48) );
  AOI222_X1 U76 ( .A1(data_out_b[11]), .A2(n22), .B1(adder[11]), .B2(n21), 
        .C1(n68), .C2(n52), .ZN(n53) );
  INV_X1 U77 ( .A(n53), .ZN(n81) );
  AOI222_X1 U78 ( .A1(data_out_b[10]), .A2(n22), .B1(adder[10]), .B2(n21), 
        .C1(n68), .C2(n54), .ZN(n55) );
  INV_X1 U79 ( .A(n55), .ZN(n82) );
  AOI222_X1 U80 ( .A1(data_out_b[8]), .A2(n22), .B1(adder[8]), .B2(n21), .C1(
        n68), .C2(f[8]), .ZN(n56) );
  INV_X1 U81 ( .A(n56), .ZN(n84) );
  AOI222_X1 U82 ( .A1(data_out_b[7]), .A2(n22), .B1(adder[7]), .B2(n21), .C1(
        n68), .C2(f[7]), .ZN(n57) );
  INV_X1 U83 ( .A(n57), .ZN(n85) );
  AOI222_X1 U84 ( .A1(data_out_b[6]), .A2(n22), .B1(adder[6]), .B2(n21), .C1(
        n68), .C2(f[6]), .ZN(n58) );
  INV_X1 U85 ( .A(n58), .ZN(n87) );
  AOI222_X1 U86 ( .A1(data_out_b[5]), .A2(n22), .B1(adder[5]), .B2(n21), .C1(
        n68), .C2(f[5]), .ZN(n59) );
  INV_X1 U87 ( .A(n59), .ZN(n104) );
  AOI222_X1 U88 ( .A1(data_out_b[4]), .A2(n22), .B1(adder[4]), .B2(n21), .C1(
        n68), .C2(f[4]), .ZN(n60) );
  INV_X1 U89 ( .A(n60), .ZN(n113) );
  AOI222_X1 U90 ( .A1(data_out_b[3]), .A2(n22), .B1(adder[3]), .B2(n21), .C1(
        n68), .C2(f[3]), .ZN(n61) );
  INV_X1 U91 ( .A(n61), .ZN(n114) );
  AOI222_X1 U92 ( .A1(data_out_b[2]), .A2(n22), .B1(adder[2]), .B2(n21), .C1(
        n68), .C2(n62), .ZN(n63) );
  INV_X1 U93 ( .A(n63), .ZN(n115) );
  AOI222_X1 U94 ( .A1(data_out_b[1]), .A2(n22), .B1(adder[1]), .B2(n21), .C1(
        n68), .C2(n64), .ZN(n65) );
  INV_X1 U95 ( .A(n65), .ZN(n116) );
  AOI222_X1 U96 ( .A1(data_out_b[0]), .A2(n22), .B1(adder[0]), .B2(n21), .C1(
        n68), .C2(n66), .ZN(n67) );
  INV_X1 U97 ( .A(n67), .ZN(n168) );
  AOI222_X1 U98 ( .A1(data_out_b[9]), .A2(n22), .B1(adder[9]), .B2(n21), .C1(
        n68), .C2(f[9]), .ZN(n69) );
  INV_X1 U99 ( .A(n69), .ZN(n83) );
  NOR4_X1 U100 ( .A1(n52), .A2(n51), .A3(n50), .A4(n49), .ZN(n77) );
  NOR4_X1 U101 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n54), .ZN(n76) );
  NAND4_X1 U102 ( .A1(n73), .A2(n72), .A3(n71), .A4(n70), .ZN(n74) );
  NOR4_X1 U103 ( .A1(n74), .A2(n66), .A3(n64), .A4(n62), .ZN(n75) );
  NAND3_X1 U104 ( .A1(n77), .A2(n76), .A3(n75), .ZN(n79) );
  NAND3_X1 U105 ( .A1(wr_en_y), .A2(n79), .A3(n78), .ZN(n246) );
  OAI22_X1 U106 ( .A1(n186), .A2(n247), .B1(n218), .B2(n246), .ZN(n185) );
  OAI22_X1 U107 ( .A1(n187), .A2(n247), .B1(n219), .B2(n246), .ZN(n184) );
  OAI22_X1 U108 ( .A1(n188), .A2(n247), .B1(n220), .B2(n246), .ZN(n183) );
  OAI22_X1 U109 ( .A1(n196), .A2(n247), .B1(n224), .B2(n246), .ZN(n175) );
  OAI22_X1 U110 ( .A1(n197), .A2(n247), .B1(n225), .B2(n246), .ZN(n174) );
  OAI22_X1 U111 ( .A1(n198), .A2(n247), .B1(n226), .B2(n246), .ZN(n173) );
  OAI22_X1 U112 ( .A1(n199), .A2(n247), .B1(n227), .B2(n246), .ZN(n172) );
  OAI22_X1 U113 ( .A1(n200), .A2(n247), .B1(n228), .B2(n246), .ZN(n171) );
  OAI22_X1 U114 ( .A1(n201), .A2(n247), .B1(n78), .B2(n246), .ZN(n170) );
endmodule


module layer1_8_4_8_16_datapath_M8_N4_T16_P8_5_DW_mult_tc_1 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n9, n12, n13, n16, n18, n19, n21, n23, n25, n27, n29, n31,
         n32, n34, n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n50,
         n52, n53, n54, n55, n56, n57, n58, n59, n62, n63, n64, n65, n67, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n93, n95, n96, n97, n98, n99,
         n103, n104, n105, n106, n107, n109, n111, n112, n113, n114, n115,
         n117, n119, n120, n122, n125, n127, n131, n133, n135, n139, n141,
         n142, n143, n145, n146, n147, n148, n149, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n237, n247, n249, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n418, n419, n420, n421, n422, n423, n424, n426, n427, n429,
         n430, n431, n490, n491, n492, n493, n494, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U150 ( .A(n271), .B(n146), .Z(n147) );
  XOR2_X1 U152 ( .A(n301), .B(n148), .Z(n149) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U161 ( .A(n177), .B(n168), .CI(n166), .CO(n163), .S(n164) );
  FA_X1 U162 ( .A(n170), .B(n172), .CI(n179), .CO(n165), .S(n166) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n291), .CI(n263), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n317), .B(n252), .CO(n173), .S(n174) );
  FA_X1 U167 ( .A(n180), .B(n187), .CI(n178), .CO(n175), .S(n176) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U169 ( .A(n193), .B(n282), .CI(n191), .CO(n179), .S(n180) );
  FA_X1 U170 ( .A(n268), .B(n292), .CI(n274), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U172 ( .A(n197), .B(n190), .CI(n188), .CO(n185), .S(n186) );
  FA_X1 U173 ( .A(n199), .B(n201), .CI(n192), .CO(n187), .S(n188) );
  FA_X1 U174 ( .A(n275), .B(n293), .CI(n194), .CO(n189), .S(n190) );
  FA_X1 U175 ( .A(n283), .B(n305), .CI(n253), .CO(n191), .S(n192) );
  HA_X1 U176 ( .A(n269), .B(n319), .CO(n193), .S(n194) );
  FA_X1 U177 ( .A(n205), .B(n200), .CI(n198), .CO(n195), .S(n196) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U179 ( .A(n284), .B(n294), .CI(n276), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n320), .B(n270), .CI(n306), .CO(n201), .S(n202) );
  FA_X1 U181 ( .A(n208), .B(n213), .CI(n206), .CO(n203), .S(n204) );
  FA_X1 U182 ( .A(n215), .B(n307), .CI(n210), .CO(n205), .S(n206) );
  FA_X1 U183 ( .A(n295), .B(n285), .CI(n254), .CO(n207), .S(n208) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U185 ( .A(n216), .B(n219), .CI(n214), .CO(n211), .S(n212) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n322), .B(n278), .CI(n308), .CO(n215), .S(n216) );
  FA_X1 U188 ( .A(n225), .B(n222), .CI(n220), .CO(n217), .S(n218) );
  FA_X1 U189 ( .A(n255), .B(n309), .CI(n297), .CO(n219), .S(n220) );
  HA_X1 U190 ( .A(n287), .B(n323), .CO(n221), .S(n222) );
  FA_X1 U191 ( .A(n229), .B(n298), .CI(n226), .CO(n223), .S(n224) );
  FA_X1 U192 ( .A(n288), .B(n310), .CI(n324), .CO(n225), .S(n226) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  HA_X1 U194 ( .A(n311), .B(n325), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n326), .B(n300), .CI(n312), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  BUF_X1 U414 ( .A(n115), .Z(n490) );
  BUF_X2 U415 ( .A(n9), .Z(n547) );
  CLKBUF_X1 U416 ( .A(n104), .Z(n493) );
  OR2_X1 U417 ( .A1(n196), .A2(n203), .ZN(n491) );
  XOR2_X1 U418 ( .A(n553), .B(n249), .Z(n492) );
  BUF_X2 U419 ( .A(n37), .Z(n494) );
  XNOR2_X1 U420 ( .A(n562), .B(a[8]), .ZN(n429) );
  AND2_X1 U421 ( .A1(n224), .A2(n227), .ZN(n497) );
  NAND2_X1 U422 ( .A1(n429), .A2(n27), .ZN(n29) );
  XNOR2_X1 U423 ( .A(n507), .B(n420), .ZN(n338) );
  INV_X1 U424 ( .A(n497), .ZN(n103) );
  AND2_X1 U425 ( .A1(n496), .A2(n122), .ZN(product[1]) );
  OR2_X1 U426 ( .A1(n329), .A2(n258), .ZN(n496) );
  OR2_X2 U427 ( .A1(n227), .A2(n224), .ZN(n542) );
  NOR2_X1 U428 ( .A1(n186), .A2(n195), .ZN(n498) );
  NOR2_X1 U429 ( .A1(n186), .A2(n195), .ZN(n82) );
  AOI21_X1 U430 ( .B1(n80), .B2(n530), .A(n81), .ZN(n45) );
  CLKBUF_X3 U431 ( .A(n19), .Z(n523) );
  XNOR2_X1 U432 ( .A(n533), .B(n499), .ZN(product[12]) );
  AND2_X1 U433 ( .A1(n517), .A2(n79), .ZN(n499) );
  OAI21_X1 U434 ( .B1(n105), .B2(n107), .A(n106), .ZN(n104) );
  OR2_X1 U435 ( .A1(n204), .A2(n211), .ZN(n500) );
  CLKBUF_X1 U436 ( .A(n533), .Z(n501) );
  XOR2_X1 U437 ( .A(n559), .B(a[6]), .Z(n21) );
  XNOR2_X1 U438 ( .A(n88), .B(n502), .ZN(product[10]) );
  NAND2_X1 U439 ( .A1(n491), .A2(n86), .ZN(n502) );
  INV_X2 U440 ( .A(n516), .ZN(n503) );
  INV_X1 U441 ( .A(n516), .ZN(n16) );
  INV_X1 U442 ( .A(n512), .ZN(n504) );
  BUF_X2 U443 ( .A(n9), .Z(n505) );
  OR2_X2 U444 ( .A1(n492), .A2(n249), .ZN(n506) );
  INV_X1 U445 ( .A(n564), .ZN(n507) );
  INV_X1 U446 ( .A(n564), .ZN(n508) );
  INV_X1 U447 ( .A(n564), .ZN(n563) );
  CLKBUF_X1 U448 ( .A(n27), .Z(n509) );
  INV_X1 U449 ( .A(n552), .ZN(n510) );
  INV_X2 U450 ( .A(n553), .ZN(n552) );
  INV_X1 U451 ( .A(n562), .ZN(n511) );
  INV_X1 U452 ( .A(n562), .ZN(n561) );
  INV_X1 U453 ( .A(n559), .ZN(n512) );
  INV_X1 U454 ( .A(n559), .ZN(n557) );
  INV_X1 U455 ( .A(n553), .ZN(n551) );
  OR2_X2 U456 ( .A1(n513), .A2(n529), .ZN(n34) );
  XNOR2_X1 U457 ( .A(n563), .B(a[10]), .ZN(n513) );
  INV_X1 U458 ( .A(n524), .ZN(n534) );
  XOR2_X1 U459 ( .A(n553), .B(a[2]), .Z(n514) );
  CLKBUF_X1 U460 ( .A(n27), .Z(n515) );
  XNOR2_X1 U461 ( .A(n556), .B(a[2]), .ZN(n536) );
  INV_X1 U462 ( .A(n556), .ZN(n554) );
  XNOR2_X1 U463 ( .A(n556), .B(a[4]), .ZN(n516) );
  INV_X1 U464 ( .A(n525), .ZN(n27) );
  OR2_X1 U465 ( .A1(n176), .A2(n185), .ZN(n517) );
  OAI21_X1 U466 ( .B1(n519), .B2(n97), .A(n98), .ZN(n518) );
  AOI21_X1 U467 ( .B1(n104), .B2(n542), .A(n497), .ZN(n519) );
  OAI21_X1 U468 ( .B1(n99), .B2(n97), .A(n98), .ZN(n96) );
  NAND2_X1 U469 ( .A1(n536), .A2(n514), .ZN(n520) );
  NAND2_X1 U470 ( .A1(n536), .A2(n514), .ZN(n521) );
  NAND2_X1 U471 ( .A1(n536), .A2(n514), .ZN(n12) );
  NOR2_X1 U472 ( .A1(n164), .A2(n175), .ZN(n522) );
  XNOR2_X1 U473 ( .A(n560), .B(a[6]), .ZN(n430) );
  NOR2_X1 U474 ( .A1(n164), .A2(n175), .ZN(n75) );
  INV_X1 U475 ( .A(n529), .ZN(n32) );
  XNOR2_X1 U476 ( .A(n559), .B(a[6]), .ZN(n524) );
  XNOR2_X1 U477 ( .A(n560), .B(a[8]), .ZN(n525) );
  OR2_X2 U478 ( .A1(n526), .A2(n249), .ZN(n6) );
  XOR2_X1 U479 ( .A(n553), .B(n249), .Z(n526) );
  INV_X1 U480 ( .A(n249), .ZN(n548) );
  AOI21_X1 U481 ( .B1(n96), .B2(n538), .A(n93), .ZN(n527) );
  AOI21_X1 U482 ( .B1(n518), .B2(n538), .A(n93), .ZN(n528) );
  AOI21_X1 U483 ( .B1(n96), .B2(n538), .A(n93), .ZN(n91) );
  XNOR2_X1 U484 ( .A(n562), .B(a[10]), .ZN(n529) );
  OAI21_X1 U485 ( .B1(n91), .B2(n89), .A(n90), .ZN(n530) );
  XOR2_X1 U486 ( .A(n553), .B(a[2]), .Z(n9) );
  NAND2_X1 U487 ( .A1(n431), .A2(n16), .ZN(n531) );
  NAND2_X1 U488 ( .A1(n431), .A2(n16), .ZN(n532) );
  NAND2_X1 U489 ( .A1(n431), .A2(n16), .ZN(n18) );
  AOI21_X1 U490 ( .B1(n80), .B2(n530), .A(n81), .ZN(n533) );
  XNOR2_X1 U491 ( .A(n557), .B(a[6]), .ZN(n535) );
  OR2_X1 U492 ( .A1(n152), .A2(n163), .ZN(n537) );
  NAND2_X1 U493 ( .A1(n537), .A2(n69), .ZN(n47) );
  INV_X1 U494 ( .A(n73), .ZN(n71) );
  AOI21_X1 U495 ( .B1(n74), .B2(n537), .A(n67), .ZN(n65) );
  INV_X1 U496 ( .A(n69), .ZN(n67) );
  INV_X1 U497 ( .A(n74), .ZN(n72) );
  INV_X1 U498 ( .A(n95), .ZN(n93) );
  NAND2_X1 U499 ( .A1(n500), .A2(n90), .ZN(n52) );
  NAND2_X1 U500 ( .A1(n125), .A2(n76), .ZN(n48) );
  INV_X1 U501 ( .A(n522), .ZN(n125) );
  NAND2_X1 U502 ( .A1(n127), .A2(n83), .ZN(n50) );
  OAI21_X1 U503 ( .B1(n75), .B2(n79), .A(n76), .ZN(n74) );
  NOR2_X1 U504 ( .A1(n522), .A2(n78), .ZN(n73) );
  NAND2_X1 U505 ( .A1(n152), .A2(n163), .ZN(n69) );
  NAND2_X1 U506 ( .A1(n538), .A2(n95), .ZN(n53) );
  INV_X1 U507 ( .A(n119), .ZN(n117) );
  OAI21_X1 U508 ( .B1(n113), .B2(n115), .A(n114), .ZN(n112) );
  NAND2_X1 U509 ( .A1(n133), .A2(n106), .ZN(n56) );
  INV_X1 U510 ( .A(n105), .ZN(n133) );
  NAND2_X1 U511 ( .A1(n131), .A2(n98), .ZN(n54) );
  INV_X1 U512 ( .A(n97), .ZN(n131) );
  NOR2_X1 U513 ( .A1(n176), .A2(n185), .ZN(n78) );
  XOR2_X1 U514 ( .A(n58), .B(n490), .Z(product[3]) );
  NAND2_X1 U515 ( .A1(n135), .A2(n114), .ZN(n58) );
  NOR2_X1 U516 ( .A1(n196), .A2(n203), .ZN(n85) );
  XNOR2_X1 U517 ( .A(n63), .B(n46), .ZN(product[15]) );
  NAND2_X1 U518 ( .A1(n541), .A2(n62), .ZN(n46) );
  NAND2_X1 U519 ( .A1(n73), .A2(n537), .ZN(n64) );
  XNOR2_X1 U520 ( .A(n57), .B(n112), .ZN(product[4]) );
  NAND2_X1 U521 ( .A1(n540), .A2(n111), .ZN(n57) );
  XNOR2_X1 U522 ( .A(n59), .B(n120), .ZN(product[2]) );
  NAND2_X1 U523 ( .A1(n539), .A2(n119), .ZN(n59) );
  NAND2_X1 U524 ( .A1(n176), .A2(n185), .ZN(n79) );
  NAND2_X1 U525 ( .A1(n164), .A2(n175), .ZN(n76) );
  NAND2_X1 U526 ( .A1(n212), .A2(n217), .ZN(n95) );
  INV_X1 U527 ( .A(n122), .ZN(n120) );
  OR2_X1 U528 ( .A1(n212), .A2(n217), .ZN(n538) );
  NAND2_X1 U529 ( .A1(n186), .A2(n195), .ZN(n83) );
  NAND2_X1 U530 ( .A1(n196), .A2(n203), .ZN(n86) );
  NAND2_X1 U531 ( .A1(n329), .A2(n258), .ZN(n122) );
  NAND2_X1 U532 ( .A1(n328), .A2(n314), .ZN(n119) );
  OR2_X1 U533 ( .A1(n328), .A2(n314), .ZN(n539) );
  OR2_X1 U534 ( .A1(n232), .A2(n233), .ZN(n540) );
  NAND2_X1 U535 ( .A1(n228), .A2(n231), .ZN(n106) );
  NAND2_X1 U536 ( .A1(n151), .A2(n139), .ZN(n62) );
  OR2_X1 U537 ( .A1(n151), .A2(n139), .ZN(n541) );
  XNOR2_X1 U538 ( .A(n552), .B(n549), .ZN(n408) );
  XNOR2_X1 U539 ( .A(n155), .B(n543), .ZN(n139) );
  XNOR2_X1 U540 ( .A(n153), .B(n141), .ZN(n543) );
  XNOR2_X1 U541 ( .A(n157), .B(n544), .ZN(n141) );
  XNOR2_X1 U542 ( .A(n145), .B(n143), .ZN(n544) );
  OR2_X1 U543 ( .A1(n549), .A2(n556), .ZN(n392) );
  AND2_X1 U544 ( .A1(n550), .A2(n516), .ZN(n300) );
  AND2_X1 U545 ( .A1(n550), .A2(n524), .ZN(n288) );
  AND2_X1 U546 ( .A1(n550), .A2(n525), .ZN(n278) );
  XNOR2_X1 U547 ( .A(n511), .B(n549), .ZN(n352) );
  OAI22_X1 U548 ( .A1(n42), .A2(n568), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U549 ( .A1(n549), .A2(n568), .ZN(n332) );
  XNOR2_X1 U550 ( .A(n507), .B(n549), .ZN(n343) );
  XNOR2_X1 U551 ( .A(n159), .B(n545), .ZN(n142) );
  XNOR2_X1 U552 ( .A(n315), .B(n261), .ZN(n545) );
  XNOR2_X1 U553 ( .A(n558), .B(n549), .ZN(n376) );
  INV_X1 U554 ( .A(n37), .ZN(n237) );
  XNOR2_X1 U555 ( .A(n565), .B(n549), .ZN(n336) );
  AND2_X1 U556 ( .A1(n550), .A2(n247), .ZN(n314) );
  AND2_X1 U557 ( .A1(n550), .A2(n237), .ZN(n264) );
  OAI22_X1 U558 ( .A1(n39), .A2(n336), .B1(n494), .B2(n335), .ZN(n263) );
  INV_X1 U559 ( .A(n25), .ZN(n562) );
  INV_X1 U560 ( .A(n19), .ZN(n560) );
  INV_X1 U561 ( .A(n1), .ZN(n553) );
  AND2_X1 U562 ( .A1(n550), .A2(n529), .ZN(n270) );
  AND2_X1 U563 ( .A1(n550), .A2(n235), .ZN(n260) );
  OAI22_X1 U564 ( .A1(n39), .A2(n335), .B1(n494), .B2(n334), .ZN(n262) );
  INV_X1 U565 ( .A(n7), .ZN(n556) );
  INV_X1 U566 ( .A(n13), .ZN(n559) );
  INV_X1 U567 ( .A(n41), .ZN(n235) );
  XNOR2_X1 U568 ( .A(n523), .B(n549), .ZN(n363) );
  OAI22_X1 U569 ( .A1(n39), .A2(n566), .B1(n337), .B2(n494), .ZN(n252) );
  OR2_X1 U570 ( .A1(n549), .A2(n566), .ZN(n337) );
  AND2_X1 U571 ( .A1(n550), .A2(n249), .ZN(product[0]) );
  OR2_X1 U572 ( .A1(n549), .A2(n564), .ZN(n344) );
  OR2_X1 U573 ( .A1(n549), .A2(n560), .ZN(n364) );
  OR2_X1 U574 ( .A1(n549), .A2(n562), .ZN(n353) );
  OR2_X1 U575 ( .A1(n549), .A2(n504), .ZN(n377) );
  XNOR2_X1 U576 ( .A(n565), .B(a[14]), .ZN(n41) );
  OAI22_X1 U577 ( .A1(n39), .A2(n334), .B1(n494), .B2(n333), .ZN(n261) );
  XNOR2_X1 U578 ( .A(n565), .B(n422), .ZN(n333) );
  XNOR2_X1 U579 ( .A(n558), .B(b[11]), .ZN(n365) );
  BUF_X2 U580 ( .A(n43), .Z(n549) );
  XNOR2_X1 U581 ( .A(n523), .B(b[9]), .ZN(n354) );
  OAI22_X1 U582 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U583 ( .A(n567), .B(n424), .ZN(n330) );
  XNOR2_X1 U584 ( .A(n567), .B(n549), .ZN(n331) );
  XNOR2_X1 U585 ( .A(n565), .B(n423), .ZN(n334) );
  XNOR2_X1 U586 ( .A(n565), .B(n424), .ZN(n335) );
  XNOR2_X1 U587 ( .A(n511), .B(n418), .ZN(n345) );
  XNOR2_X1 U588 ( .A(n265), .B(n546), .ZN(n145) );
  XNOR2_X1 U589 ( .A(n149), .B(n147), .ZN(n546) );
  XNOR2_X1 U590 ( .A(n555), .B(b[13]), .ZN(n378) );
  NAND2_X1 U591 ( .A1(n427), .A2(n37), .ZN(n39) );
  XNOR2_X1 U592 ( .A(n555), .B(n419), .ZN(n385) );
  XNOR2_X1 U593 ( .A(n508), .B(n422), .ZN(n340) );
  XNOR2_X1 U594 ( .A(n508), .B(n421), .ZN(n339) );
  XNOR2_X1 U595 ( .A(n508), .B(n423), .ZN(n341) );
  XNOR2_X1 U596 ( .A(n507), .B(n424), .ZN(n342) );
  XNOR2_X1 U597 ( .A(n552), .B(n423), .ZN(n406) );
  XNOR2_X1 U598 ( .A(n551), .B(n422), .ZN(n405) );
  XNOR2_X1 U599 ( .A(n511), .B(n422), .ZN(n349) );
  XNOR2_X1 U600 ( .A(n523), .B(n423), .ZN(n361) );
  XNOR2_X1 U601 ( .A(n523), .B(n422), .ZN(n360) );
  XNOR2_X1 U602 ( .A(n561), .B(n423), .ZN(n350) );
  XNOR2_X1 U603 ( .A(n511), .B(n420), .ZN(n347) );
  XNOR2_X1 U604 ( .A(n523), .B(n420), .ZN(n358) );
  XNOR2_X1 U605 ( .A(n561), .B(n421), .ZN(n348) );
  XNOR2_X1 U606 ( .A(n523), .B(n421), .ZN(n359) );
  XNOR2_X1 U607 ( .A(n551), .B(n420), .ZN(n403) );
  XNOR2_X1 U608 ( .A(n551), .B(n421), .ZN(n404) );
  XNOR2_X1 U609 ( .A(n511), .B(n419), .ZN(n346) );
  XNOR2_X1 U610 ( .A(n523), .B(n419), .ZN(n357) );
  XNOR2_X1 U611 ( .A(n551), .B(n419), .ZN(n402) );
  XNOR2_X1 U612 ( .A(n561), .B(n424), .ZN(n351) );
  XNOR2_X1 U613 ( .A(n523), .B(n424), .ZN(n362) );
  XNOR2_X1 U614 ( .A(n552), .B(n424), .ZN(n407) );
  NAND2_X1 U615 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U616 ( .A(n567), .B(a[14]), .Z(n426) );
  CLKBUF_X1 U617 ( .A(n43), .Z(n550) );
  XNOR2_X1 U618 ( .A(n555), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U619 ( .A(n555), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U620 ( .A(n555), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U621 ( .A(n555), .B(n418), .ZN(n384) );
  XNOR2_X1 U622 ( .A(n555), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U623 ( .A(n555), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U624 ( .A(n558), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U625 ( .A(n558), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U626 ( .A(n558), .B(n418), .ZN(n369) );
  XNOR2_X1 U627 ( .A(n558), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U628 ( .A(n552), .B(b[14]), .ZN(n394) );
  XNOR2_X1 U629 ( .A(n552), .B(b[13]), .ZN(n395) );
  XNOR2_X1 U630 ( .A(n552), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U631 ( .A(n552), .B(b[11]), .ZN(n397) );
  XNOR2_X1 U632 ( .A(n523), .B(b[8]), .ZN(n355) );
  XNOR2_X1 U633 ( .A(n523), .B(n418), .ZN(n356) );
  XNOR2_X1 U634 ( .A(n551), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U635 ( .A(n552), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U636 ( .A(n552), .B(n418), .ZN(n401) );
  XNOR2_X1 U637 ( .A(n551), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U638 ( .A(n552), .B(b[15]), .ZN(n393) );
  OAI22_X1 U639 ( .A1(n34), .A2(n339), .B1(n338), .B2(n32), .ZN(n265) );
  OAI22_X1 U640 ( .A1(n34), .A2(n340), .B1(n339), .B2(n32), .ZN(n266) );
  OAI22_X1 U641 ( .A1(n34), .A2(n341), .B1(n340), .B2(n32), .ZN(n267) );
  OAI22_X1 U642 ( .A1(n34), .A2(n342), .B1(n341), .B2(n32), .ZN(n268) );
  OAI22_X1 U643 ( .A1(n34), .A2(n343), .B1(n342), .B2(n32), .ZN(n269) );
  OAI22_X1 U644 ( .A1(n34), .A2(n564), .B1(n344), .B2(n32), .ZN(n253) );
  XOR2_X1 U645 ( .A(n565), .B(a[12]), .Z(n427) );
  XNOR2_X1 U646 ( .A(n563), .B(a[12]), .ZN(n37) );
  NAND2_X1 U647 ( .A1(n218), .A2(n223), .ZN(n98) );
  NOR2_X1 U648 ( .A1(n218), .A2(n223), .ZN(n97) );
  OAI22_X1 U649 ( .A1(n506), .A2(n394), .B1(n393), .B2(n548), .ZN(n315) );
  OAI22_X1 U650 ( .A1(n6), .A2(n395), .B1(n394), .B2(n548), .ZN(n316) );
  OAI22_X1 U651 ( .A1(n506), .A2(n396), .B1(n395), .B2(n548), .ZN(n317) );
  OAI22_X1 U652 ( .A1(n506), .A2(n397), .B1(n396), .B2(n548), .ZN(n318) );
  OAI22_X1 U653 ( .A1(n6), .A2(n398), .B1(n397), .B2(n548), .ZN(n319) );
  OAI22_X1 U654 ( .A1(n506), .A2(n399), .B1(n398), .B2(n548), .ZN(n320) );
  OAI22_X1 U655 ( .A1(n6), .A2(n400), .B1(n399), .B2(n548), .ZN(n321) );
  OAI22_X1 U656 ( .A1(n6), .A2(n408), .B1(n407), .B2(n548), .ZN(n329) );
  OAI22_X1 U657 ( .A1(n6), .A2(n407), .B1(n406), .B2(n548), .ZN(n328) );
  OAI22_X1 U658 ( .A1(n506), .A2(n406), .B1(n405), .B2(n548), .ZN(n327) );
  OAI22_X1 U659 ( .A1(n6), .A2(n405), .B1(n404), .B2(n548), .ZN(n326) );
  OAI22_X1 U660 ( .A1(n506), .A2(n404), .B1(n403), .B2(n548), .ZN(n325) );
  OAI22_X1 U661 ( .A1(n6), .A2(n403), .B1(n402), .B2(n548), .ZN(n324) );
  OAI22_X1 U662 ( .A1(n6), .A2(n402), .B1(n401), .B2(n548), .ZN(n323) );
  OAI22_X1 U663 ( .A1(n506), .A2(n401), .B1(n400), .B2(n548), .ZN(n322) );
  NOR2_X1 U664 ( .A1(n228), .A2(n231), .ZN(n105) );
  INV_X1 U665 ( .A(n113), .ZN(n135) );
  NOR2_X1 U666 ( .A1(n234), .A2(n257), .ZN(n113) );
  NAND2_X1 U667 ( .A1(n232), .A2(n233), .ZN(n111) );
  NAND2_X1 U668 ( .A1(n542), .A2(n103), .ZN(n55) );
  XNOR2_X1 U669 ( .A(n84), .B(n50), .ZN(product[11]) );
  NAND2_X1 U670 ( .A1(n204), .A2(n211), .ZN(n90) );
  NOR2_X1 U671 ( .A1(n204), .A2(n211), .ZN(n89) );
  OAI22_X1 U672 ( .A1(n29), .A2(n346), .B1(n345), .B2(n515), .ZN(n271) );
  OAI22_X1 U673 ( .A1(n29), .A2(n347), .B1(n346), .B2(n515), .ZN(n272) );
  OAI22_X1 U674 ( .A1(n29), .A2(n350), .B1(n349), .B2(n515), .ZN(n275) );
  OAI22_X1 U675 ( .A1(n29), .A2(n351), .B1(n350), .B2(n509), .ZN(n276) );
  OAI22_X1 U676 ( .A1(n29), .A2(n348), .B1(n347), .B2(n509), .ZN(n273) );
  OAI22_X1 U677 ( .A1(n29), .A2(n562), .B1(n353), .B2(n27), .ZN(n254) );
  OAI22_X1 U678 ( .A1(n29), .A2(n349), .B1(n348), .B2(n509), .ZN(n274) );
  OAI22_X1 U679 ( .A1(n29), .A2(n352), .B1(n351), .B2(n509), .ZN(n277) );
  XNOR2_X1 U680 ( .A(n512), .B(n424), .ZN(n375) );
  XNOR2_X1 U681 ( .A(n512), .B(n419), .ZN(n370) );
  XNOR2_X1 U682 ( .A(n557), .B(n420), .ZN(n371) );
  XNOR2_X1 U683 ( .A(n512), .B(n423), .ZN(n374) );
  XNOR2_X1 U684 ( .A(n512), .B(n422), .ZN(n373) );
  XNOR2_X1 U685 ( .A(n512), .B(n421), .ZN(n372) );
  XOR2_X1 U686 ( .A(n557), .B(a[4]), .Z(n431) );
  XNOR2_X1 U687 ( .A(n554), .B(n420), .ZN(n386) );
  XNOR2_X1 U688 ( .A(n554), .B(n549), .ZN(n391) );
  XNOR2_X1 U689 ( .A(n554), .B(n422), .ZN(n388) );
  XNOR2_X1 U690 ( .A(n554), .B(n424), .ZN(n390) );
  XNOR2_X1 U691 ( .A(n554), .B(n423), .ZN(n389) );
  XNOR2_X1 U692 ( .A(n554), .B(n421), .ZN(n387) );
  XNOR2_X1 U693 ( .A(n77), .B(n48), .ZN(product[13]) );
  AOI21_X1 U694 ( .B1(n539), .B2(n120), .A(n117), .ZN(n115) );
  INV_X1 U695 ( .A(n498), .ZN(n127) );
  NOR2_X1 U696 ( .A1(n498), .A2(n85), .ZN(n80) );
  OAI21_X1 U697 ( .B1(n82), .B2(n86), .A(n83), .ZN(n81) );
  OAI21_X1 U698 ( .B1(n87), .B2(n85), .A(n86), .ZN(n84) );
  OAI22_X1 U699 ( .A1(n506), .A2(n510), .B1(n409), .B2(n548), .ZN(n258) );
  OR2_X1 U700 ( .A1(n549), .A2(n510), .ZN(n409) );
  INV_X1 U701 ( .A(n88), .ZN(n87) );
  OAI22_X1 U702 ( .A1(n23), .A2(n358), .B1(n357), .B2(n535), .ZN(n282) );
  OAI22_X1 U703 ( .A1(n23), .A2(n356), .B1(n355), .B2(n534), .ZN(n280) );
  OAI22_X1 U704 ( .A1(n23), .A2(n362), .B1(n361), .B2(n535), .ZN(n286) );
  OAI22_X1 U705 ( .A1(n23), .A2(n560), .B1(n364), .B2(n535), .ZN(n255) );
  OAI22_X1 U706 ( .A1(n23), .A2(n357), .B1(n356), .B2(n534), .ZN(n281) );
  OAI22_X1 U707 ( .A1(n23), .A2(n355), .B1(n354), .B2(n534), .ZN(n279) );
  OAI22_X1 U708 ( .A1(n23), .A2(n361), .B1(n360), .B2(n535), .ZN(n285) );
  OAI22_X1 U709 ( .A1(n23), .A2(n360), .B1(n359), .B2(n534), .ZN(n284) );
  OAI22_X1 U710 ( .A1(n23), .A2(n363), .B1(n362), .B2(n534), .ZN(n287) );
  OAI22_X1 U711 ( .A1(n23), .A2(n359), .B1(n358), .B2(n535), .ZN(n283) );
  NAND2_X2 U712 ( .A1(n430), .A2(n21), .ZN(n23) );
  OAI22_X1 U713 ( .A1(n532), .A2(n375), .B1(n374), .B2(n503), .ZN(n298) );
  OAI22_X1 U714 ( .A1(n532), .A2(n370), .B1(n369), .B2(n503), .ZN(n293) );
  OAI22_X1 U715 ( .A1(n531), .A2(n376), .B1(n375), .B2(n503), .ZN(n299) );
  OAI22_X1 U716 ( .A1(n532), .A2(n504), .B1(n377), .B2(n503), .ZN(n256) );
  OAI22_X1 U717 ( .A1(n531), .A2(n367), .B1(n366), .B2(n503), .ZN(n290) );
  OAI22_X1 U718 ( .A1(n531), .A2(n373), .B1(n372), .B2(n503), .ZN(n296) );
  OAI22_X1 U719 ( .A1(n532), .A2(n372), .B1(n371), .B2(n503), .ZN(n295) );
  OAI22_X1 U720 ( .A1(n531), .A2(n366), .B1(n365), .B2(n503), .ZN(n289) );
  OAI22_X1 U721 ( .A1(n18), .A2(n374), .B1(n373), .B2(n503), .ZN(n297) );
  OAI22_X1 U722 ( .A1(n531), .A2(n368), .B1(n367), .B2(n503), .ZN(n291) );
  OAI22_X1 U723 ( .A1(n18), .A2(n371), .B1(n370), .B2(n503), .ZN(n294) );
  OAI22_X1 U724 ( .A1(n532), .A2(n369), .B1(n368), .B2(n503), .ZN(n292) );
  XOR2_X1 U725 ( .A(n528), .B(n52), .Z(product[9]) );
  OAI21_X1 U726 ( .B1(n527), .B2(n89), .A(n90), .ZN(n88) );
  XNOR2_X1 U727 ( .A(n518), .B(n53), .ZN(product[8]) );
  AOI21_X1 U728 ( .B1(n542), .B2(n104), .A(n497), .ZN(n99) );
  XNOR2_X1 U729 ( .A(n55), .B(n493), .ZN(product[6]) );
  XOR2_X1 U730 ( .A(n54), .B(n519), .Z(product[7]) );
  OAI21_X1 U731 ( .B1(n45), .B2(n78), .A(n79), .ZN(n77) );
  OAI21_X1 U732 ( .B1(n45), .B2(n71), .A(n72), .ZN(n70) );
  XNOR2_X1 U733 ( .A(n70), .B(n47), .ZN(product[14]) );
  OAI21_X1 U734 ( .B1(n64), .B2(n501), .A(n65), .ZN(n63) );
  XOR2_X1 U735 ( .A(n56), .B(n107), .Z(product[5]) );
  AOI21_X1 U736 ( .B1(n540), .B2(n112), .A(n109), .ZN(n107) );
  INV_X1 U737 ( .A(n111), .ZN(n109) );
  OAI22_X1 U738 ( .A1(n520), .A2(n379), .B1(n378), .B2(n505), .ZN(n301) );
  OAI22_X1 U739 ( .A1(n520), .A2(n380), .B1(n379), .B2(n505), .ZN(n302) );
  OAI22_X1 U740 ( .A1(n521), .A2(n385), .B1(n384), .B2(n505), .ZN(n307) );
  OAI22_X1 U741 ( .A1(n521), .A2(n382), .B1(n381), .B2(n505), .ZN(n304) );
  OAI22_X1 U742 ( .A1(n520), .A2(n381), .B1(n380), .B2(n505), .ZN(n303) );
  NAND2_X1 U743 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U744 ( .A1(n520), .A2(n383), .B1(n382), .B2(n547), .ZN(n305) );
  OAI22_X1 U745 ( .A1(n521), .A2(n384), .B1(n383), .B2(n547), .ZN(n306) );
  OAI22_X1 U746 ( .A1(n520), .A2(n386), .B1(n385), .B2(n505), .ZN(n308) );
  OAI22_X1 U747 ( .A1(n521), .A2(n387), .B1(n386), .B2(n505), .ZN(n309) );
  OAI22_X1 U748 ( .A1(n521), .A2(n556), .B1(n392), .B2(n505), .ZN(n257) );
  OAI22_X1 U749 ( .A1(n12), .A2(n389), .B1(n388), .B2(n505), .ZN(n311) );
  OAI22_X1 U750 ( .A1(n12), .A2(n388), .B1(n387), .B2(n547), .ZN(n310) );
  OAI22_X1 U751 ( .A1(n12), .A2(n390), .B1(n389), .B2(n547), .ZN(n312) );
  INV_X1 U752 ( .A(n505), .ZN(n247) );
  OAI22_X1 U753 ( .A1(n520), .A2(n391), .B1(n390), .B2(n505), .ZN(n313) );
  INV_X1 U754 ( .A(n556), .ZN(n555) );
  INV_X1 U755 ( .A(n559), .ZN(n558) );
  INV_X1 U756 ( .A(n31), .ZN(n564) );
  INV_X1 U757 ( .A(n566), .ZN(n565) );
  INV_X1 U758 ( .A(n36), .ZN(n566) );
  INV_X1 U759 ( .A(n568), .ZN(n567) );
  INV_X1 U760 ( .A(n40), .ZN(n568) );
  XOR2_X1 U761 ( .A(n259), .B(n251), .Z(n148) );
  XOR2_X1 U762 ( .A(n289), .B(n279), .Z(n146) );
endmodule


module layer1_8_4_8_16_datapath_M8_N4_T16_P8_5_DW01_add_2 ( A, B, CI, SUM, CO
 );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n18,
         n19, n20, n21, n23, n25, n26, n27, n28, n30, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n48, n49, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n71, n72, n73,
         n74, n75, n77, n79, n80, n81, n82, n83, n85, n87, n88, n90, n93, n98,
         n99, n100, n102, n104, n161, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186;

  OR2_X1 U126 ( .A1(A[11]), .A2(B[11]), .ZN(n161) );
  AND2_X1 U127 ( .A1(n178), .A2(n90), .ZN(SUM[0]) );
  NOR2_X1 U128 ( .A1(A[8]), .A2(B[8]), .ZN(n163) );
  NOR2_X1 U129 ( .A1(A[8]), .A2(B[8]), .ZN(n58) );
  AOI21_X1 U130 ( .B1(n56), .B2(n64), .A(n57), .ZN(n164) );
  AOI21_X1 U131 ( .B1(n56), .B2(n64), .A(n57), .ZN(n55) );
  BUF_X1 U132 ( .A(n169), .Z(n165) );
  AND2_X1 U133 ( .A1(A[9]), .A2(B[9]), .ZN(n166) );
  BUF_X1 U134 ( .A(n40), .Z(n169) );
  NAND2_X1 U135 ( .A1(A[12]), .A2(B[12]), .ZN(n167) );
  XNOR2_X1 U136 ( .A(n172), .B(n5), .ZN(SUM[11]) );
  OR2_X1 U137 ( .A1(A[12]), .A2(B[12]), .ZN(n168) );
  AOI21_X1 U138 ( .B1(n185), .B2(n166), .A(n186), .ZN(n170) );
  NOR2_X1 U139 ( .A1(n36), .A2(n39), .ZN(n171) );
  NOR2_X2 U140 ( .A1(A[11]), .A2(B[11]), .ZN(n39) );
  OAI21_X1 U141 ( .B1(n43), .B2(n55), .A(n170), .ZN(n172) );
  NOR2_X1 U142 ( .A1(A[12]), .A2(B[12]), .ZN(n173) );
  NOR2_X1 U143 ( .A1(A[12]), .A2(B[12]), .ZN(n174) );
  NOR2_X1 U144 ( .A1(A[12]), .A2(B[12]), .ZN(n36) );
  OAI21_X1 U145 ( .B1(n40), .B2(n174), .A(n167), .ZN(n175) );
  OR2_X2 U146 ( .A1(A[10]), .A2(B[10]), .ZN(n185) );
  AOI21_X1 U147 ( .B1(n42), .B2(n34), .A(n35), .ZN(n176) );
  AOI21_X1 U148 ( .B1(n42), .B2(n171), .A(n175), .ZN(n177) );
  OR2_X1 U149 ( .A1(A[0]), .A2(B[0]), .ZN(n178) );
  INV_X1 U150 ( .A(n172), .ZN(n41) );
  INV_X1 U151 ( .A(n71), .ZN(n69) );
  INV_X1 U152 ( .A(n87), .ZN(n85) );
  NOR2_X1 U153 ( .A1(n163), .A2(n61), .ZN(n56) );
  OAI21_X1 U154 ( .B1(n83), .B2(n81), .A(n82), .ZN(n80) );
  AOI21_X1 U155 ( .B1(n182), .B2(n80), .A(n77), .ZN(n75) );
  INV_X1 U156 ( .A(n79), .ZN(n77) );
  AOI21_X1 U157 ( .B1(n172), .B2(n171), .A(n175), .ZN(n33) );
  AOI21_X1 U158 ( .B1(n180), .B2(n54), .A(n166), .ZN(n49) );
  INV_X1 U159 ( .A(n61), .ZN(n99) );
  INV_X1 U160 ( .A(n90), .ZN(n88) );
  NAND2_X1 U161 ( .A1(n98), .A2(n59), .ZN(n8) );
  INV_X1 U162 ( .A(n163), .ZN(n98) );
  NAND2_X1 U163 ( .A1(n180), .A2(n53), .ZN(n7) );
  NAND2_X1 U164 ( .A1(n100), .A2(n66), .ZN(n10) );
  INV_X1 U165 ( .A(n65), .ZN(n100) );
  NAND2_X1 U166 ( .A1(n102), .A2(n74), .ZN(n12) );
  INV_X1 U167 ( .A(n73), .ZN(n102) );
  NAND2_X1 U168 ( .A1(n183), .A2(n87), .ZN(n15) );
  NAND2_X1 U169 ( .A1(n182), .A2(n79), .ZN(n13) );
  NAND2_X1 U170 ( .A1(n179), .A2(n71), .ZN(n11) );
  NAND2_X1 U171 ( .A1(n104), .A2(n82), .ZN(n14) );
  INV_X1 U172 ( .A(n81), .ZN(n104) );
  XNOR2_X1 U173 ( .A(n38), .B(n4), .ZN(SUM[12]) );
  NAND2_X1 U174 ( .A1(n168), .A2(n167), .ZN(n4) );
  XOR2_X1 U175 ( .A(n49), .B(n6), .Z(SUM[10]) );
  XNOR2_X1 U176 ( .A(n54), .B(n7), .ZN(SUM[9]) );
  XNOR2_X1 U177 ( .A(n60), .B(n8), .ZN(SUM[8]) );
  XOR2_X1 U178 ( .A(n63), .B(n9), .Z(SUM[7]) );
  XNOR2_X1 U179 ( .A(n13), .B(n80), .ZN(SUM[3]) );
  XNOR2_X1 U180 ( .A(n15), .B(n88), .ZN(SUM[1]) );
  NAND2_X1 U181 ( .A1(n161), .A2(n169), .ZN(n5) );
  NOR2_X1 U182 ( .A1(A[7]), .A2(B[7]), .ZN(n61) );
  OR2_X1 U183 ( .A1(A[5]), .A2(B[5]), .ZN(n179) );
  OR2_X1 U184 ( .A1(A[9]), .A2(B[9]), .ZN(n180) );
  NAND2_X1 U185 ( .A1(A[11]), .A2(B[11]), .ZN(n40) );
  NAND2_X1 U186 ( .A1(A[3]), .A2(B[3]), .ZN(n79) );
  OR2_X1 U187 ( .A1(A[14]), .A2(B[14]), .ZN(n181) );
  NOR2_X1 U188 ( .A1(A[2]), .A2(B[2]), .ZN(n81) );
  NOR2_X1 U189 ( .A1(A[6]), .A2(B[6]), .ZN(n65) );
  NOR2_X1 U190 ( .A1(A[4]), .A2(B[4]), .ZN(n73) );
  OR2_X1 U191 ( .A1(A[3]), .A2(B[3]), .ZN(n182) );
  NAND2_X1 U192 ( .A1(A[1]), .A2(B[1]), .ZN(n87) );
  NAND2_X1 U193 ( .A1(A[5]), .A2(B[5]), .ZN(n71) );
  NAND2_X1 U194 ( .A1(A[0]), .A2(B[0]), .ZN(n90) );
  NAND2_X1 U195 ( .A1(A[2]), .A2(B[2]), .ZN(n82) );
  NAND2_X1 U196 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  OR2_X1 U197 ( .A1(A[1]), .A2(B[1]), .ZN(n183) );
  NAND2_X1 U198 ( .A1(A[6]), .A2(B[6]), .ZN(n66) );
  NAND2_X1 U199 ( .A1(A[4]), .A2(B[4]), .ZN(n74) );
  OR2_X1 U200 ( .A1(A[15]), .A2(B[15]), .ZN(n184) );
  XOR2_X1 U201 ( .A(n10), .B(n67), .Z(SUM[6]) );
  XOR2_X1 U202 ( .A(n12), .B(n75), .Z(SUM[4]) );
  INV_X1 U203 ( .A(n186), .ZN(n48) );
  OAI21_X1 U204 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  OAI21_X1 U205 ( .B1(n58), .B2(n62), .A(n59), .ZN(n57) );
  NAND2_X1 U206 ( .A1(n99), .A2(n62), .ZN(n9) );
  NAND2_X1 U207 ( .A1(A[7]), .A2(B[7]), .ZN(n62) );
  NAND2_X1 U208 ( .A1(A[8]), .A2(B[8]), .ZN(n59) );
  AND2_X1 U209 ( .A1(A[10]), .A2(B[10]), .ZN(n186) );
  INV_X1 U210 ( .A(n28), .ZN(n30) );
  NAND2_X1 U211 ( .A1(A[12]), .A2(B[12]), .ZN(n37) );
  AOI21_X1 U212 ( .B1(n179), .B2(n72), .A(n69), .ZN(n67) );
  XNOR2_X1 U213 ( .A(n11), .B(n72), .ZN(SUM[5]) );
  OAI21_X1 U214 ( .B1(n75), .B2(n73), .A(n74), .ZN(n72) );
  NAND2_X1 U215 ( .A1(A[9]), .A2(B[9]), .ZN(n53) );
  INV_X1 U216 ( .A(n164), .ZN(n54) );
  AOI21_X1 U217 ( .B1(n181), .B2(n30), .A(n23), .ZN(n21) );
  NAND2_X1 U218 ( .A1(A[15]), .A2(B[15]), .ZN(n18) );
  INV_X1 U219 ( .A(n25), .ZN(n23) );
  NAND2_X1 U220 ( .A1(n181), .A2(n25), .ZN(n2) );
  NAND2_X1 U221 ( .A1(n93), .A2(n181), .ZN(n20) );
  NAND2_X1 U222 ( .A1(n93), .A2(n28), .ZN(n3) );
  INV_X1 U223 ( .A(n27), .ZN(n93) );
  AOI21_X1 U224 ( .B1(n183), .B2(n88), .A(n85), .ZN(n83) );
  INV_X1 U225 ( .A(n64), .ZN(n63) );
  XOR2_X1 U226 ( .A(n14), .B(n83), .Z(SUM[2]) );
  NAND2_X1 U227 ( .A1(A[14]), .A2(B[14]), .ZN(n25) );
  OAI21_X1 U228 ( .B1(n173), .B2(n40), .A(n37), .ZN(n35) );
  NOR2_X1 U229 ( .A1(n36), .A2(n39), .ZN(n34) );
  OAI21_X1 U230 ( .B1(n67), .B2(n65), .A(n66), .ZN(n64) );
  NOR2_X1 U231 ( .A1(A[13]), .A2(B[13]), .ZN(n27) );
  XNOR2_X1 U232 ( .A(n26), .B(n2), .ZN(SUM[14]) );
  XNOR2_X1 U233 ( .A(n19), .B(n1), .ZN(SUM[15]) );
  NAND2_X1 U234 ( .A1(n184), .A2(n18), .ZN(n1) );
  OAI21_X1 U235 ( .B1(n41), .B2(n39), .A(n165), .ZN(n38) );
  NAND2_X1 U236 ( .A1(n185), .A2(n48), .ZN(n6) );
  NAND2_X1 U237 ( .A1(n185), .A2(n180), .ZN(n43) );
  AOI21_X1 U238 ( .B1(n185), .B2(n166), .A(n186), .ZN(n44) );
  XOR2_X1 U239 ( .A(n33), .B(n3), .Z(SUM[13]) );
  OAI21_X1 U240 ( .B1(n176), .B2(n27), .A(n28), .ZN(n26) );
  OAI21_X1 U241 ( .B1(n177), .B2(n20), .A(n21), .ZN(n19) );
  OAI21_X1 U242 ( .B1(n43), .B2(n55), .A(n44), .ZN(n42) );
endmodule


module layer1_8_4_8_16_datapath_M8_N4_T16_P8_5 ( clk, clear_acc, data_out_x, 
        data_out, data_out_w, data_out_b, wr_en_y, m_valid, m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [3:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N27, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, n1, n2, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n87, n104, n113, n114, n115, n116, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n20), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n227), .CK(clk), .Q(n25) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n228), .CK(clk), .Q(n26) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n229), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n230), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n231), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n232), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n233), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n234), .CK(clk), .Q(n34) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n235), .CK(clk), .Q(n35) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n236), .CK(clk), .Q(n36) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n237), .CK(clk), .Q(n37) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n238), .CK(clk), .Q(n38) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n239), .CK(clk), .Q(n39) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n240), .CK(clk), .Q(n40) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n241), .CK(clk), .Q(n41) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n242), .CK(clk), .Q(n43) );
  DFF_X1 \f_reg[0]  ( .D(n115), .CK(clk), .Q(n64), .QN(n216) );
  DFF_X1 \f_reg[1]  ( .D(n114), .CK(clk), .Q(n62), .QN(n217) );
  DFF_X1 \f_reg[2]  ( .D(n113), .CK(clk), .Q(n60), .QN(n218) );
  DFF_X1 \f_reg[3]  ( .D(n104), .CK(clk), .Q(f[3]), .QN(n68) );
  DFF_X1 \f_reg[4]  ( .D(n87), .CK(clk), .Q(f[4]), .QN(n69) );
  DFF_X1 \f_reg[5]  ( .D(n85), .CK(clk), .Q(f[5]), .QN(n70) );
  DFF_X1 \f_reg[6]  ( .D(n84), .CK(clk), .Q(f[6]), .QN(n71) );
  DFF_X1 \f_reg[7]  ( .D(n83), .CK(clk), .Q(f[7]), .QN(n219) );
  DFF_X1 \f_reg[8]  ( .D(n82), .CK(clk), .Q(f[8]), .QN(n220) );
  DFF_X1 \f_reg[9]  ( .D(n81), .CK(clk), .Q(f[9]), .QN(n221) );
  DFF_X1 \f_reg[10]  ( .D(n80), .CK(clk), .Q(n52), .QN(n222) );
  DFF_X1 \f_reg[11]  ( .D(n79), .CK(clk), .Q(n50), .QN(n223) );
  DFF_X1 \f_reg[12]  ( .D(n4), .CK(clk), .Q(n49), .QN(n224) );
  DFF_X1 \f_reg[13]  ( .D(n2), .CK(clk), .Q(n48), .QN(n225) );
  DFF_X1 \f_reg[14]  ( .D(n5), .CK(clk), .Q(n47), .QN(n226) );
  DFF_X1 \f_reg[15]  ( .D(n78), .CK(clk), .Q(f[15]), .QN(n76) );
  DFF_X1 \data_out_reg[15]  ( .D(n168), .CK(clk), .Q(data_out[15]), .QN(n199)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n169), .CK(clk), .Q(data_out[14]), .QN(n198)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n170), .CK(clk), .Q(data_out[13]), .QN(n197)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n171), .CK(clk), .Q(data_out[12]), .QN(n196)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n172), .CK(clk), .Q(data_out[11]), .QN(n195)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n173), .CK(clk), .Q(data_out[10]), .QN(n194)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n174), .CK(clk), .Q(data_out[9]), .QN(n193) );
  DFF_X1 \data_out_reg[8]  ( .D(n175), .CK(clk), .Q(data_out[8]), .QN(n192) );
  DFF_X1 \data_out_reg[7]  ( .D(n176), .CK(clk), .Q(data_out[7]), .QN(n191) );
  DFF_X1 \data_out_reg[6]  ( .D(n177), .CK(clk), .Q(data_out[6]), .QN(n190) );
  DFF_X1 \data_out_reg[5]  ( .D(n178), .CK(clk), .Q(data_out[5]), .QN(n189) );
  DFF_X1 \data_out_reg[4]  ( .D(n179), .CK(clk), .Q(data_out[4]), .QN(n188) );
  DFF_X1 \data_out_reg[3]  ( .D(n180), .CK(clk), .Q(data_out[3]), .QN(n187) );
  DFF_X1 \data_out_reg[2]  ( .D(n181), .CK(clk), .Q(data_out[2]), .QN(n186) );
  DFF_X1 \data_out_reg[1]  ( .D(n182), .CK(clk), .Q(data_out[1]), .QN(n185) );
  DFF_X1 \data_out_reg[0]  ( .D(n183), .CK(clk), .Q(data_out[0]), .QN(n184) );
  layer1_8_4_8_16_datapath_M8_N4_T16_P8_5_DW_mult_tc_1 mult_183 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer1_8_4_8_16_datapath_M8_N4_T16_P8_5_DW01_add_2 add_184 ( .A({n206, n205, 
        n204, n203, n202, n201, n215, n214, n213, n212, n211, n210, n209, n208, 
        n207, n200}), .B({f[15], n47, n48, n49, n50, n52, f[9:3], n60, n62, 
        n64}), .CI(1'b0), .SUM(adder) );
  DFF_X2 delay_reg ( .D(N27), .CK(clk), .Q(n1), .QN(n243) );
  MUX2_X2 U3 ( .A(n33), .B(N38), .S(n243), .Z(n215) );
  NAND3_X1 U4 ( .A1(n14), .A2(n13), .A3(n15), .ZN(n2) );
  NAND3_X1 U5 ( .A1(n8), .A2(n7), .A3(n9), .ZN(n4) );
  MUX2_X2 U6 ( .A(n27), .B(N42), .S(n243), .Z(n204) );
  NAND3_X1 U8 ( .A1(n17), .A2(n16), .A3(n18), .ZN(n5) );
  MUX2_X2 U9 ( .A(n29), .B(N40), .S(n243), .Z(n202) );
  AND2_X1 U10 ( .A1(n12), .A2(n10), .ZN(n6) );
  NAND2_X1 U11 ( .A1(n11), .A2(n6), .ZN(n78) );
  MUX2_X2 U12 ( .A(n34), .B(N37), .S(n243), .Z(n214) );
  MUX2_X2 U13 ( .A(n28), .B(N41), .S(n243), .Z(n203) );
  NAND2_X1 U14 ( .A1(data_out_b[12]), .A2(n20), .ZN(n7) );
  NAND2_X1 U15 ( .A1(adder[12]), .A2(n19), .ZN(n8) );
  NAND2_X1 U16 ( .A1(n66), .A2(n49), .ZN(n9) );
  NAND2_X1 U17 ( .A1(data_out_b[15]), .A2(n20), .ZN(n10) );
  NAND2_X1 U18 ( .A1(adder[15]), .A2(n19), .ZN(n11) );
  NAND2_X1 U19 ( .A1(n66), .A2(f[15]), .ZN(n12) );
  NAND2_X1 U20 ( .A1(data_out_b[13]), .A2(n20), .ZN(n13) );
  NAND2_X1 U21 ( .A1(adder[13]), .A2(n19), .ZN(n14) );
  NAND2_X1 U22 ( .A1(n66), .A2(n48), .ZN(n15) );
  NAND2_X1 U23 ( .A1(data_out_b[14]), .A2(n20), .ZN(n16) );
  NAND2_X1 U24 ( .A1(adder[14]), .A2(n19), .ZN(n17) );
  NAND2_X1 U25 ( .A1(n66), .A2(n47), .ZN(n18) );
  INV_X1 U26 ( .A(n21), .ZN(n20) );
  AND2_X2 U27 ( .A1(n46), .A2(n21), .ZN(n19) );
  INV_X1 U28 ( .A(n46), .ZN(n66) );
  INV_X1 U29 ( .A(clear_acc), .ZN(n21) );
  NAND2_X1 U30 ( .A1(n116), .A2(N27), .ZN(n245) );
  INV_X1 U31 ( .A(wr_en_y), .ZN(n116) );
  OAI22_X1 U32 ( .A1(n187), .A2(n245), .B1(n68), .B2(n244), .ZN(n180) );
  OAI22_X1 U33 ( .A1(n188), .A2(n245), .B1(n69), .B2(n244), .ZN(n179) );
  OAI22_X1 U34 ( .A1(n189), .A2(n245), .B1(n70), .B2(n244), .ZN(n178) );
  OAI22_X1 U35 ( .A1(n190), .A2(n245), .B1(n71), .B2(n244), .ZN(n177) );
  OAI22_X1 U36 ( .A1(n191), .A2(n245), .B1(n219), .B2(n244), .ZN(n176) );
  OAI22_X1 U37 ( .A1(n192), .A2(n245), .B1(n220), .B2(n244), .ZN(n175) );
  OAI22_X1 U38 ( .A1(n193), .A2(n245), .B1(n221), .B2(n244), .ZN(n174) );
  INV_X1 U39 ( .A(n24), .ZN(n42) );
  MUX2_X1 U40 ( .A(n39), .B(N32), .S(n243), .Z(n209) );
  MUX2_X1 U41 ( .A(n26), .B(N43), .S(n243), .Z(n205) );
  AND3_X1 U42 ( .A1(sel[1]), .A2(sel[2]), .A3(sel[0]), .ZN(n23) );
  INV_X1 U43 ( .A(m_ready), .ZN(n22) );
  NAND2_X1 U44 ( .A1(m_valid), .A2(n22), .ZN(n44) );
  OAI21_X1 U45 ( .B1(sel[3]), .B2(n23), .A(n44), .ZN(N27) );
  NAND2_X1 U46 ( .A1(clear_acc_delay), .A2(n243), .ZN(n24) );
  MUX2_X1 U47 ( .A(n25), .B(N44), .S(n42), .Z(n227) );
  MUX2_X1 U48 ( .A(n25), .B(N44), .S(n243), .Z(n206) );
  MUX2_X1 U49 ( .A(n26), .B(N43), .S(n42), .Z(n228) );
  MUX2_X1 U50 ( .A(n27), .B(N42), .S(n42), .Z(n229) );
  MUX2_X1 U51 ( .A(n28), .B(N41), .S(n42), .Z(n230) );
  MUX2_X1 U52 ( .A(n29), .B(N40), .S(n42), .Z(n231) );
  MUX2_X1 U53 ( .A(n32), .B(N39), .S(n42), .Z(n232) );
  MUX2_X1 U54 ( .A(n32), .B(N39), .S(n243), .Z(n201) );
  MUX2_X1 U55 ( .A(n33), .B(N38), .S(n42), .Z(n233) );
  MUX2_X1 U56 ( .A(n34), .B(N37), .S(n42), .Z(n234) );
  MUX2_X1 U57 ( .A(n35), .B(N36), .S(n42), .Z(n235) );
  MUX2_X1 U58 ( .A(n35), .B(N36), .S(n243), .Z(n213) );
  MUX2_X1 U59 ( .A(n36), .B(N35), .S(n42), .Z(n236) );
  MUX2_X1 U60 ( .A(n36), .B(N35), .S(n243), .Z(n212) );
  MUX2_X1 U61 ( .A(n37), .B(N34), .S(n42), .Z(n237) );
  MUX2_X1 U62 ( .A(n37), .B(N34), .S(n243), .Z(n211) );
  MUX2_X1 U63 ( .A(n38), .B(N33), .S(n42), .Z(n238) );
  MUX2_X1 U64 ( .A(n38), .B(N33), .S(n243), .Z(n210) );
  MUX2_X1 U65 ( .A(n39), .B(N32), .S(n42), .Z(n239) );
  MUX2_X1 U66 ( .A(n40), .B(N31), .S(n42), .Z(n240) );
  MUX2_X1 U67 ( .A(n40), .B(N31), .S(n243), .Z(n208) );
  MUX2_X1 U68 ( .A(n41), .B(N30), .S(n42), .Z(n241) );
  MUX2_X1 U69 ( .A(n41), .B(N30), .S(n243), .Z(n207) );
  MUX2_X1 U70 ( .A(n43), .B(N29), .S(n42), .Z(n242) );
  MUX2_X1 U71 ( .A(n43), .B(N29), .S(n243), .Z(n200) );
  INV_X1 U72 ( .A(n44), .ZN(n45) );
  OAI21_X1 U73 ( .B1(n45), .B2(n1), .A(n21), .ZN(n46) );
  AOI222_X1 U74 ( .A1(data_out_b[11]), .A2(n20), .B1(adder[11]), .B2(n19), 
        .C1(n66), .C2(n50), .ZN(n51) );
  INV_X1 U75 ( .A(n51), .ZN(n79) );
  AOI222_X1 U76 ( .A1(data_out_b[10]), .A2(n20), .B1(adder[10]), .B2(n19), 
        .C1(n66), .C2(n52), .ZN(n53) );
  INV_X1 U77 ( .A(n53), .ZN(n80) );
  AOI222_X1 U78 ( .A1(data_out_b[8]), .A2(n20), .B1(adder[8]), .B2(n19), .C1(
        n66), .C2(f[8]), .ZN(n54) );
  INV_X1 U79 ( .A(n54), .ZN(n82) );
  AOI222_X1 U80 ( .A1(data_out_b[7]), .A2(n20), .B1(adder[7]), .B2(n19), .C1(
        n66), .C2(f[7]), .ZN(n55) );
  INV_X1 U81 ( .A(n55), .ZN(n83) );
  AOI222_X1 U82 ( .A1(data_out_b[6]), .A2(n20), .B1(adder[6]), .B2(n19), .C1(
        n66), .C2(f[6]), .ZN(n56) );
  INV_X1 U83 ( .A(n56), .ZN(n84) );
  AOI222_X1 U84 ( .A1(data_out_b[5]), .A2(n20), .B1(adder[5]), .B2(n19), .C1(
        n66), .C2(f[5]), .ZN(n57) );
  INV_X1 U85 ( .A(n57), .ZN(n85) );
  AOI222_X1 U86 ( .A1(data_out_b[4]), .A2(n20), .B1(adder[4]), .B2(n19), .C1(
        n66), .C2(f[4]), .ZN(n58) );
  INV_X1 U87 ( .A(n58), .ZN(n87) );
  AOI222_X1 U88 ( .A1(data_out_b[3]), .A2(n20), .B1(adder[3]), .B2(n19), .C1(
        n66), .C2(f[3]), .ZN(n59) );
  INV_X1 U89 ( .A(n59), .ZN(n104) );
  AOI222_X1 U90 ( .A1(data_out_b[2]), .A2(n20), .B1(adder[2]), .B2(n19), .C1(
        n66), .C2(n60), .ZN(n61) );
  INV_X1 U91 ( .A(n61), .ZN(n113) );
  AOI222_X1 U92 ( .A1(data_out_b[1]), .A2(n20), .B1(adder[1]), .B2(n19), .C1(
        n66), .C2(n62), .ZN(n63) );
  INV_X1 U93 ( .A(n63), .ZN(n114) );
  AOI222_X1 U94 ( .A1(data_out_b[0]), .A2(n20), .B1(adder[0]), .B2(n19), .C1(
        n66), .C2(n64), .ZN(n65) );
  INV_X1 U95 ( .A(n65), .ZN(n115) );
  AOI222_X1 U96 ( .A1(data_out_b[9]), .A2(n20), .B1(adder[9]), .B2(n19), .C1(
        n66), .C2(f[9]), .ZN(n67) );
  INV_X1 U97 ( .A(n67), .ZN(n81) );
  NOR4_X1 U98 ( .A1(n50), .A2(n49), .A3(n48), .A4(n47), .ZN(n75) );
  NOR4_X1 U99 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n52), .ZN(n74) );
  NAND4_X1 U100 ( .A1(n71), .A2(n70), .A3(n69), .A4(n68), .ZN(n72) );
  NOR4_X1 U101 ( .A1(n72), .A2(n64), .A3(n62), .A4(n60), .ZN(n73) );
  NAND3_X1 U102 ( .A1(n75), .A2(n74), .A3(n73), .ZN(n77) );
  NAND3_X1 U103 ( .A1(wr_en_y), .A2(n77), .A3(n76), .ZN(n244) );
  OAI22_X1 U104 ( .A1(n184), .A2(n245), .B1(n216), .B2(n244), .ZN(n183) );
  OAI22_X1 U105 ( .A1(n185), .A2(n245), .B1(n217), .B2(n244), .ZN(n182) );
  OAI22_X1 U106 ( .A1(n186), .A2(n245), .B1(n218), .B2(n244), .ZN(n181) );
  OAI22_X1 U107 ( .A1(n194), .A2(n245), .B1(n222), .B2(n244), .ZN(n173) );
  OAI22_X1 U108 ( .A1(n195), .A2(n245), .B1(n223), .B2(n244), .ZN(n172) );
  OAI22_X1 U109 ( .A1(n196), .A2(n245), .B1(n224), .B2(n244), .ZN(n171) );
  OAI22_X1 U110 ( .A1(n197), .A2(n245), .B1(n225), .B2(n244), .ZN(n170) );
  OAI22_X1 U111 ( .A1(n198), .A2(n245), .B1(n226), .B2(n244), .ZN(n169) );
  OAI22_X1 U112 ( .A1(n199), .A2(n245), .B1(n76), .B2(n244), .ZN(n168) );
endmodule


module layer1_8_4_8_16_datapath_M8_N4_T16_P8_4_DW_mult_tc_1 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n12, n13, n16, n18, n19, n21, n23, n25, n27, n29, n31,
         n32, n34, n36, n37, n39, n40, n41, n42, n43, n46, n47, n48, n50, n51,
         n53, n55, n56, n57, n58, n59, n62, n63, n64, n65, n67, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n93, n95, n96, n97, n98, n99, n101,
         n103, n104, n105, n106, n107, n109, n111, n112, n113, n114, n115,
         n117, n119, n120, n122, n127, n135, n139, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n237, n243, n245, n249, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n418,
         n419, n420, n421, n422, n423, n424, n426, n427, n428, n429, n430,
         n490, n491, n492, n493, n494, n495, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U148 ( .A(n265), .B(n144), .Z(n145) );
  XOR2_X1 U150 ( .A(n271), .B(n146), .Z(n147) );
  XOR2_X1 U152 ( .A(n301), .B(n148), .Z(n149) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U162 ( .A(n170), .B(n172), .CI(n179), .CO(n165), .S(n166) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n263), .CI(n291), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n317), .B(n252), .CO(n173), .S(n174) );
  FA_X1 U167 ( .A(n180), .B(n187), .CI(n178), .CO(n175), .S(n176) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U169 ( .A(n193), .B(n282), .CI(n191), .CO(n179), .S(n180) );
  FA_X1 U170 ( .A(n268), .B(n274), .CI(n292), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U172 ( .A(n197), .B(n190), .CI(n188), .CO(n185), .S(n186) );
  FA_X1 U173 ( .A(n199), .B(n201), .CI(n192), .CO(n187), .S(n188) );
  FA_X1 U174 ( .A(n275), .B(n293), .CI(n194), .CO(n189), .S(n190) );
  FA_X1 U175 ( .A(n253), .B(n305), .CI(n283), .CO(n191), .S(n192) );
  HA_X1 U176 ( .A(n319), .B(n269), .CO(n193), .S(n194) );
  FA_X1 U177 ( .A(n205), .B(n200), .CI(n198), .CO(n195), .S(n196) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U179 ( .A(n276), .B(n284), .CI(n294), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n320), .B(n270), .CI(n306), .CO(n201), .S(n202) );
  FA_X1 U181 ( .A(n208), .B(n213), .CI(n206), .CO(n203), .S(n204) );
  FA_X1 U182 ( .A(n215), .B(n307), .CI(n210), .CO(n205), .S(n206) );
  FA_X1 U183 ( .A(n254), .B(n295), .CI(n285), .CO(n207), .S(n208) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n322), .B(n278), .CI(n308), .CO(n215), .S(n216) );
  FA_X1 U188 ( .A(n225), .B(n222), .CI(n220), .CO(n217), .S(n218) );
  FA_X1 U189 ( .A(n309), .B(n255), .CI(n297), .CO(n219), .S(n220) );
  HA_X1 U190 ( .A(n287), .B(n323), .CO(n221), .S(n222) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  HA_X1 U194 ( .A(n311), .B(n325), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n312), .B(n300), .CI(n326), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  CLKBUF_X1 U414 ( .A(n228), .Z(n490) );
  NAND2_X1 U415 ( .A1(n196), .A2(n203), .ZN(n491) );
  CLKBUF_X1 U416 ( .A(n83), .Z(n492) );
  NOR2_X1 U417 ( .A1(n526), .A2(n85), .ZN(n493) );
  CLKBUF_X2 U418 ( .A(n7), .Z(n494) );
  XNOR2_X1 U419 ( .A(n166), .B(n495), .ZN(n164) );
  XNOR2_X1 U420 ( .A(n177), .B(n168), .ZN(n495) );
  BUF_X1 U421 ( .A(n603), .Z(n581) );
  BUF_X1 U422 ( .A(n32), .Z(n560) );
  OR2_X1 U423 ( .A1(n573), .A2(n249), .ZN(n6) );
  AND2_X1 U424 ( .A1(n498), .A2(n122), .ZN(product[1]) );
  OR2_X1 U425 ( .A1(n164), .A2(n175), .ZN(n497) );
  OR2_X1 U426 ( .A1(n329), .A2(n258), .ZN(n498) );
  XNOR2_X1 U427 ( .A(n583), .B(n499), .ZN(product[7]) );
  AND2_X1 U428 ( .A1(n523), .A2(n98), .ZN(n499) );
  CLKBUF_X1 U429 ( .A(n112), .Z(n500) );
  INV_X1 U430 ( .A(n608), .ZN(n501) );
  FA_X1 U431 ( .A(n205), .B(n200), .CI(n198), .S(n502) );
  NAND2_X1 U432 ( .A1(n429), .A2(n27), .ZN(n503) );
  NAND2_X1 U433 ( .A1(n429), .A2(n27), .ZN(n504) );
  NAND2_X1 U434 ( .A1(n429), .A2(n27), .ZN(n29) );
  CLKBUF_X1 U435 ( .A(n18), .Z(n558) );
  CLKBUF_X1 U436 ( .A(n18), .Z(n557) );
  INV_X1 U437 ( .A(n577), .ZN(n505) );
  BUF_X1 U438 ( .A(n605), .Z(n543) );
  CLKBUF_X1 U439 ( .A(n549), .Z(n506) );
  XNOR2_X1 U440 ( .A(n507), .B(n226), .ZN(n224) );
  XNOR2_X1 U441 ( .A(n229), .B(n298), .ZN(n507) );
  BUF_X1 U442 ( .A(n106), .Z(n508) );
  CLKBUF_X1 U443 ( .A(n559), .Z(n525) );
  XNOR2_X1 U444 ( .A(n582), .B(n509), .ZN(product[9]) );
  AND2_X1 U445 ( .A1(n555), .A2(n90), .ZN(n509) );
  XNOR2_X1 U446 ( .A(n612), .B(a[8]), .ZN(n429) );
  XOR2_X1 U447 ( .A(n581), .B(n418), .Z(n401) );
  CLKBUF_X1 U448 ( .A(n226), .Z(n510) );
  OR2_X2 U449 ( .A1(n573), .A2(n249), .ZN(n511) );
  INV_X1 U450 ( .A(n7), .ZN(n512) );
  BUF_X1 U451 ( .A(n401), .Z(n513) );
  XNOR2_X1 U452 ( .A(n613), .B(a[10]), .ZN(n428) );
  XNOR2_X1 U453 ( .A(n214), .B(n514), .ZN(n212) );
  XNOR2_X1 U454 ( .A(n216), .B(n219), .ZN(n514) );
  BUF_X1 U455 ( .A(n18), .Z(n534) );
  NAND2_X1 U456 ( .A1(n214), .A2(n216), .ZN(n515) );
  NAND2_X1 U457 ( .A1(n214), .A2(n219), .ZN(n516) );
  NAND2_X1 U458 ( .A1(n216), .A2(n219), .ZN(n517) );
  NAND3_X1 U459 ( .A1(n515), .A2(n516), .A3(n517), .ZN(n211) );
  INV_X2 U460 ( .A(n603), .ZN(n602) );
  CLKBUF_X1 U461 ( .A(n491), .Z(n518) );
  CLKBUF_X1 U462 ( .A(n571), .Z(n519) );
  INV_X2 U463 ( .A(n581), .ZN(n598) );
  NAND2_X1 U464 ( .A1(n166), .A2(n177), .ZN(n520) );
  NAND2_X1 U465 ( .A1(n166), .A2(n168), .ZN(n521) );
  NAND2_X1 U466 ( .A1(n177), .A2(n168), .ZN(n522) );
  NAND3_X1 U467 ( .A1(n520), .A2(n521), .A3(n522), .ZN(n163) );
  OR2_X1 U468 ( .A1(n218), .A2(n223), .ZN(n523) );
  CLKBUF_X3 U469 ( .A(n16), .Z(n529) );
  NOR2_X1 U470 ( .A1(n164), .A2(n175), .ZN(n524) );
  NOR2_X1 U471 ( .A1(n164), .A2(n175), .ZN(n75) );
  NOR2_X1 U472 ( .A1(n186), .A2(n195), .ZN(n526) );
  NOR2_X1 U473 ( .A1(n186), .A2(n195), .ZN(n82) );
  INV_X1 U474 ( .A(n580), .ZN(n527) );
  INV_X1 U475 ( .A(n540), .ZN(n528) );
  BUF_X2 U476 ( .A(n609), .Z(n539) );
  CLKBUF_X1 U477 ( .A(n16), .Z(n596) );
  INV_X1 U478 ( .A(n613), .ZN(n530) );
  INV_X1 U479 ( .A(n613), .ZN(n531) );
  INV_X1 U480 ( .A(n541), .ZN(n579) );
  INV_X1 U481 ( .A(n572), .ZN(n532) );
  INV_X1 U482 ( .A(n572), .ZN(n27) );
  BUF_X1 U483 ( .A(n18), .Z(n533) );
  INV_X1 U484 ( .A(n548), .ZN(n535) );
  INV_X1 U485 ( .A(n543), .ZN(n536) );
  BUF_X1 U486 ( .A(n609), .Z(n538) );
  BUF_X1 U487 ( .A(n382), .Z(n537) );
  BUF_X1 U488 ( .A(n609), .Z(n540) );
  INV_X1 U489 ( .A(n610), .ZN(n609) );
  AOI21_X1 U490 ( .B1(n96), .B2(n586), .A(n93), .ZN(n91) );
  XNOR2_X1 U491 ( .A(n603), .B(a[2]), .ZN(n541) );
  XNOR2_X1 U492 ( .A(n603), .B(a[2]), .ZN(n542) );
  XNOR2_X1 U493 ( .A(n531), .B(a[12]), .ZN(n544) );
  XNOR2_X1 U494 ( .A(n530), .B(a[12]), .ZN(n545) );
  INV_X1 U495 ( .A(n612), .ZN(n546) );
  INV_X1 U496 ( .A(n612), .ZN(n611) );
  OR2_X1 U497 ( .A1(n502), .A2(n203), .ZN(n547) );
  INV_X1 U498 ( .A(n608), .ZN(n548) );
  NAND2_X1 U499 ( .A1(n428), .A2(n32), .ZN(n549) );
  OR2_X1 U500 ( .A1(n176), .A2(n185), .ZN(n550) );
  NAND2_X1 U501 ( .A1(n430), .A2(n594), .ZN(n551) );
  NAND2_X1 U502 ( .A1(n430), .A2(n594), .ZN(n552) );
  NAND2_X1 U503 ( .A1(n430), .A2(n594), .ZN(n23) );
  XNOR2_X1 U504 ( .A(n553), .B(n310), .ZN(n226) );
  XNOR2_X1 U505 ( .A(n559), .B(n288), .ZN(n553) );
  AOI21_X1 U506 ( .B1(n568), .B2(n493), .A(n81), .ZN(n554) );
  OR2_X1 U507 ( .A1(n204), .A2(n211), .ZN(n555) );
  AOI21_X1 U508 ( .B1(n589), .B2(n112), .A(n109), .ZN(n556) );
  OAI22_X1 U509 ( .A1(n6), .A2(n403), .B1(n402), .B2(n597), .ZN(n559) );
  INV_X1 U510 ( .A(n577), .ZN(n32) );
  NAND2_X1 U511 ( .A1(n428), .A2(n505), .ZN(n34) );
  NAND2_X1 U512 ( .A1(n525), .A2(n288), .ZN(n561) );
  NAND2_X1 U513 ( .A1(n525), .A2(n310), .ZN(n562) );
  NAND2_X1 U514 ( .A1(n288), .A2(n310), .ZN(n563) );
  NAND3_X1 U515 ( .A1(n561), .A2(n562), .A3(n563), .ZN(n225) );
  NAND2_X1 U516 ( .A1(n229), .A2(n298), .ZN(n564) );
  NAND2_X1 U517 ( .A1(n229), .A2(n510), .ZN(n565) );
  NAND2_X1 U518 ( .A1(n298), .A2(n510), .ZN(n566) );
  NAND3_X1 U519 ( .A1(n564), .A2(n565), .A3(n566), .ZN(n223) );
  XOR2_X1 U520 ( .A(n605), .B(a[2]), .Z(n574) );
  INV_X1 U521 ( .A(n543), .ZN(n604) );
  XOR2_X1 U522 ( .A(n603), .B(n249), .Z(n573) );
  OAI21_X1 U523 ( .B1(n527), .B2(n556), .A(n508), .ZN(n567) );
  OAI21_X1 U524 ( .B1(n91), .B2(n89), .A(n90), .ZN(n568) );
  INV_X1 U525 ( .A(n494), .ZN(n569) );
  OAI21_X1 U526 ( .B1(n89), .B2(n91), .A(n90), .ZN(n88) );
  OR2_X2 U527 ( .A1(n574), .A2(n542), .ZN(n576) );
  XNOR2_X1 U528 ( .A(n610), .B(a[6]), .ZN(n430) );
  OAI21_X1 U529 ( .B1(n105), .B2(n107), .A(n106), .ZN(n104) );
  CLKBUF_X1 U530 ( .A(n96), .Z(n570) );
  AOI21_X1 U531 ( .B1(n80), .B2(n88), .A(n81), .ZN(n571) );
  XNOR2_X1 U532 ( .A(n610), .B(a[8]), .ZN(n572) );
  XOR2_X1 U533 ( .A(n512), .B(a[4]), .Z(n16) );
  XOR2_X1 U534 ( .A(n608), .B(a[6]), .Z(n21) );
  INV_X1 U535 ( .A(n608), .ZN(n606) );
  OR2_X1 U536 ( .A1(n574), .A2(n541), .ZN(n12) );
  OR2_X2 U537 ( .A1(n574), .A2(n542), .ZN(n575) );
  XNOR2_X1 U538 ( .A(n612), .B(a[10]), .ZN(n577) );
  INV_X1 U539 ( .A(n542), .ZN(n578) );
  OR2_X1 U540 ( .A1(n490), .A2(n231), .ZN(n580) );
  CLKBUF_X3 U541 ( .A(n21), .Z(n595) );
  BUF_X1 U542 ( .A(n21), .Z(n594) );
  CLKBUF_X1 U543 ( .A(n91), .Z(n582) );
  AOI21_X1 U544 ( .B1(n590), .B2(n567), .A(n101), .ZN(n583) );
  NAND2_X1 U545 ( .A1(n16), .A2(n584), .ZN(n18) );
  XOR2_X1 U546 ( .A(n606), .B(a[4]), .Z(n584) );
  NAND2_X1 U547 ( .A1(n585), .A2(n69), .ZN(n47) );
  INV_X1 U548 ( .A(n73), .ZN(n71) );
  INV_X1 U549 ( .A(n69), .ZN(n67) );
  NAND2_X1 U550 ( .A1(n73), .A2(n585), .ZN(n64) );
  INV_X1 U551 ( .A(n74), .ZN(n72) );
  NOR2_X1 U552 ( .A1(n526), .A2(n85), .ZN(n80) );
  OAI21_X1 U553 ( .B1(n82), .B2(n86), .A(n83), .ZN(n81) );
  INV_X1 U554 ( .A(n95), .ZN(n93) );
  NAND2_X1 U555 ( .A1(n127), .A2(n492), .ZN(n50) );
  INV_X1 U556 ( .A(n526), .ZN(n127) );
  OR2_X1 U557 ( .A1(n152), .A2(n163), .ZN(n585) );
  NAND2_X1 U558 ( .A1(n497), .A2(n76), .ZN(n48) );
  NAND2_X1 U559 ( .A1(n547), .A2(n491), .ZN(n51) );
  OAI21_X1 U560 ( .B1(n524), .B2(n79), .A(n76), .ZN(n74) );
  NOR2_X1 U561 ( .A1(n75), .A2(n78), .ZN(n73) );
  XNOR2_X1 U562 ( .A(n570), .B(n53), .ZN(product[8]) );
  NAND2_X1 U563 ( .A1(n586), .A2(n95), .ZN(n53) );
  NAND2_X1 U564 ( .A1(n152), .A2(n163), .ZN(n69) );
  INV_X1 U565 ( .A(n103), .ZN(n101) );
  OAI21_X1 U566 ( .B1(n113), .B2(n115), .A(n114), .ZN(n112) );
  OAI21_X1 U567 ( .B1(n99), .B2(n97), .A(n98), .ZN(n96) );
  AOI21_X1 U568 ( .B1(n589), .B2(n112), .A(n109), .ZN(n107) );
  INV_X1 U569 ( .A(n111), .ZN(n109) );
  AOI21_X1 U570 ( .B1(n588), .B2(n120), .A(n117), .ZN(n115) );
  INV_X1 U571 ( .A(n119), .ZN(n117) );
  NOR2_X1 U572 ( .A1(n176), .A2(n185), .ZN(n78) );
  NOR2_X1 U573 ( .A1(n502), .A2(n203), .ZN(n85) );
  XOR2_X1 U574 ( .A(n58), .B(n115), .Z(product[3]) );
  INV_X1 U575 ( .A(n113), .ZN(n135) );
  INV_X1 U576 ( .A(n122), .ZN(n120) );
  XNOR2_X1 U577 ( .A(n59), .B(n120), .ZN(product[2]) );
  NAND2_X1 U578 ( .A1(n588), .A2(n119), .ZN(n59) );
  NAND2_X1 U579 ( .A1(n196), .A2(n203), .ZN(n86) );
  NAND2_X1 U580 ( .A1(n164), .A2(n175), .ZN(n76) );
  NAND2_X1 U581 ( .A1(n186), .A2(n195), .ZN(n83) );
  OR2_X1 U582 ( .A1(n212), .A2(n217), .ZN(n586) );
  NAND2_X1 U583 ( .A1(n176), .A2(n185), .ZN(n79) );
  NAND2_X1 U584 ( .A1(n212), .A2(n217), .ZN(n95) );
  XNOR2_X1 U585 ( .A(n567), .B(n55), .ZN(product[6]) );
  NAND2_X1 U586 ( .A1(n590), .A2(n103), .ZN(n55) );
  XNOR2_X1 U587 ( .A(n57), .B(n500), .ZN(product[4]) );
  NAND2_X1 U588 ( .A1(n589), .A2(n111), .ZN(n57) );
  XNOR2_X1 U589 ( .A(n63), .B(n46), .ZN(product[15]) );
  NAND2_X1 U590 ( .A1(n587), .A2(n62), .ZN(n46) );
  AOI21_X1 U591 ( .B1(n74), .B2(n585), .A(n67), .ZN(n65) );
  NAND2_X1 U592 ( .A1(n580), .A2(n508), .ZN(n56) );
  OR2_X1 U593 ( .A1(n151), .A2(n139), .ZN(n587) );
  NAND2_X1 U594 ( .A1(n329), .A2(n258), .ZN(n122) );
  NAND2_X1 U595 ( .A1(n328), .A2(n314), .ZN(n119) );
  NOR2_X1 U596 ( .A1(n218), .A2(n223), .ZN(n97) );
  OR2_X1 U597 ( .A1(n328), .A2(n314), .ZN(n588) );
  NOR2_X1 U598 ( .A1(n228), .A2(n231), .ZN(n105) );
  NAND2_X1 U599 ( .A1(n218), .A2(n223), .ZN(n98) );
  OR2_X1 U600 ( .A1(n232), .A2(n233), .ZN(n589) );
  NAND2_X1 U601 ( .A1(n228), .A2(n231), .ZN(n106) );
  OR2_X1 U602 ( .A1(n224), .A2(n227), .ZN(n590) );
  OR2_X1 U603 ( .A1(n43), .A2(n599), .ZN(n409) );
  OR2_X1 U604 ( .A1(n43), .A2(n569), .ZN(n392) );
  XNOR2_X1 U605 ( .A(n539), .B(n43), .ZN(n363) );
  OAI22_X1 U606 ( .A1(n39), .A2(n336), .B1(n544), .B2(n335), .ZN(n263) );
  AND2_X1 U607 ( .A1(n601), .A2(n243), .ZN(n288) );
  AND2_X1 U608 ( .A1(n601), .A2(n572), .ZN(n278) );
  AND2_X1 U609 ( .A1(n601), .A2(n577), .ZN(n270) );
  AND2_X1 U610 ( .A1(n601), .A2(n237), .ZN(n264) );
  XNOR2_X1 U611 ( .A(n607), .B(n43), .ZN(n376) );
  XNOR2_X1 U612 ( .A(n155), .B(n591), .ZN(n139) );
  XNOR2_X1 U613 ( .A(n153), .B(n141), .ZN(n591) );
  XNOR2_X1 U614 ( .A(n157), .B(n592), .ZN(n141) );
  XNOR2_X1 U615 ( .A(n145), .B(n143), .ZN(n592) );
  OAI22_X1 U616 ( .A1(n42), .A2(n617), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U617 ( .A1(n43), .A2(n617), .ZN(n332) );
  XNOR2_X1 U618 ( .A(n530), .B(n43), .ZN(n343) );
  AND2_X1 U619 ( .A1(n601), .A2(n245), .ZN(n300) );
  XNOR2_X1 U620 ( .A(n159), .B(n593), .ZN(n142) );
  XNOR2_X1 U621 ( .A(n315), .B(n261), .ZN(n593) );
  INV_X1 U622 ( .A(n545), .ZN(n237) );
  XNOR2_X1 U623 ( .A(n614), .B(n43), .ZN(n336) );
  AND2_X1 U624 ( .A1(n601), .A2(n542), .ZN(n314) );
  INV_X1 U625 ( .A(n19), .ZN(n610) );
  INV_X1 U626 ( .A(n25), .ZN(n612) );
  AND2_X1 U627 ( .A1(n601), .A2(n235), .ZN(n260) );
  OAI22_X1 U628 ( .A1(n39), .A2(n335), .B1(n545), .B2(n334), .ZN(n262) );
  INV_X1 U629 ( .A(n7), .ZN(n605) );
  INV_X1 U630 ( .A(n13), .ZN(n608) );
  INV_X1 U631 ( .A(n41), .ZN(n235) );
  XNOR2_X1 U632 ( .A(n546), .B(n43), .ZN(n352) );
  OAI22_X1 U633 ( .A1(n39), .A2(n615), .B1(n337), .B2(n544), .ZN(n252) );
  OR2_X1 U634 ( .A1(n43), .A2(n615), .ZN(n337) );
  AND2_X1 U635 ( .A1(n601), .A2(n249), .ZN(product[0]) );
  OR2_X1 U636 ( .A1(n43), .A2(n528), .ZN(n364) );
  OR2_X1 U637 ( .A1(n43), .A2(n612), .ZN(n353) );
  OR2_X1 U638 ( .A1(n43), .A2(n613), .ZN(n344) );
  OR2_X1 U639 ( .A1(n43), .A2(n535), .ZN(n377) );
  XNOR2_X1 U640 ( .A(n614), .B(a[14]), .ZN(n41) );
  OAI22_X1 U641 ( .A1(n39), .A2(n334), .B1(n544), .B2(n333), .ZN(n261) );
  XNOR2_X1 U642 ( .A(n614), .B(n422), .ZN(n333) );
  XNOR2_X1 U643 ( .A(n538), .B(b[9]), .ZN(n354) );
  XNOR2_X1 U644 ( .A(n607), .B(b[11]), .ZN(n365) );
  OAI22_X1 U645 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U646 ( .A(n616), .B(n424), .ZN(n330) );
  XNOR2_X1 U647 ( .A(n616), .B(n43), .ZN(n331) );
  XNOR2_X1 U648 ( .A(n614), .B(n424), .ZN(n335) );
  XNOR2_X1 U649 ( .A(n614), .B(n423), .ZN(n334) );
  XNOR2_X1 U650 ( .A(n546), .B(n418), .ZN(n345) );
  XNOR2_X1 U651 ( .A(n530), .B(n420), .ZN(n338) );
  XNOR2_X1 U652 ( .A(n494), .B(b[13]), .ZN(n378) );
  NAND2_X1 U653 ( .A1(n427), .A2(n37), .ZN(n39) );
  XNOR2_X1 U654 ( .A(n540), .B(n424), .ZN(n362) );
  XNOR2_X1 U655 ( .A(n611), .B(n424), .ZN(n351) );
  XNOR2_X1 U656 ( .A(n531), .B(n424), .ZN(n342) );
  XNOR2_X1 U657 ( .A(n536), .B(n418), .ZN(n384) );
  XNOR2_X1 U658 ( .A(n604), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U659 ( .A(n536), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U660 ( .A(n494), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U661 ( .A(n494), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U662 ( .A(n494), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U663 ( .A(n494), .B(n419), .ZN(n385) );
  XNOR2_X1 U664 ( .A(n531), .B(n423), .ZN(n341) );
  XNOR2_X1 U665 ( .A(n530), .B(n422), .ZN(n340) );
  XNOR2_X1 U666 ( .A(n531), .B(n421), .ZN(n339) );
  XNOR2_X1 U667 ( .A(n607), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U668 ( .A(n607), .B(n418), .ZN(n369) );
  XNOR2_X1 U669 ( .A(n607), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U670 ( .A(n607), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U671 ( .A(n538), .B(n423), .ZN(n361) );
  XNOR2_X1 U672 ( .A(n539), .B(n422), .ZN(n360) );
  XNOR2_X1 U673 ( .A(n611), .B(n423), .ZN(n350) );
  XNOR2_X1 U674 ( .A(n546), .B(n422), .ZN(n349) );
  XNOR2_X1 U675 ( .A(n539), .B(n421), .ZN(n359) );
  XNOR2_X1 U676 ( .A(n538), .B(n420), .ZN(n358) );
  XNOR2_X1 U677 ( .A(n546), .B(n421), .ZN(n348) );
  XNOR2_X1 U678 ( .A(n611), .B(n420), .ZN(n347) );
  XNOR2_X1 U679 ( .A(n538), .B(n418), .ZN(n356) );
  XNOR2_X1 U680 ( .A(n539), .B(n419), .ZN(n357) );
  XNOR2_X1 U681 ( .A(n546), .B(n419), .ZN(n346) );
  XNOR2_X1 U682 ( .A(n602), .B(b[13]), .ZN(n395) );
  XNOR2_X1 U683 ( .A(n598), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U684 ( .A(n598), .B(b[14]), .ZN(n394) );
  XNOR2_X1 U685 ( .A(n539), .B(b[8]), .ZN(n355) );
  XNOR2_X1 U686 ( .A(n602), .B(b[11]), .ZN(n397) );
  NAND2_X1 U687 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U688 ( .A(n616), .B(a[14]), .Z(n426) );
  CLKBUF_X1 U689 ( .A(n43), .Z(n601) );
  XNOR2_X1 U690 ( .A(n598), .B(b[15]), .ZN(n393) );
  XOR2_X1 U691 ( .A(n614), .B(a[12]), .Z(n427) );
  XNOR2_X1 U692 ( .A(n530), .B(a[12]), .ZN(n37) );
  OAI22_X1 U693 ( .A1(n506), .A2(n339), .B1(n338), .B2(n560), .ZN(n265) );
  OAI22_X1 U694 ( .A1(n506), .A2(n340), .B1(n339), .B2(n560), .ZN(n266) );
  OAI22_X1 U695 ( .A1(n549), .A2(n342), .B1(n341), .B2(n560), .ZN(n268) );
  OAI22_X1 U696 ( .A1(n549), .A2(n341), .B1(n340), .B2(n560), .ZN(n267) );
  OAI22_X1 U697 ( .A1(n549), .A2(n343), .B1(n342), .B2(n505), .ZN(n269) );
  OAI22_X1 U698 ( .A1(n34), .A2(n613), .B1(n344), .B2(n505), .ZN(n253) );
  INV_X1 U699 ( .A(n249), .ZN(n597) );
  INV_X1 U700 ( .A(n602), .ZN(n599) );
  INV_X1 U701 ( .A(n1), .ZN(n603) );
  XNOR2_X1 U702 ( .A(n571), .B(n600), .ZN(product[12]) );
  AND2_X1 U703 ( .A1(n550), .A2(n79), .ZN(n600) );
  NAND2_X1 U704 ( .A1(n204), .A2(n211), .ZN(n90) );
  NOR2_X1 U705 ( .A1(n204), .A2(n211), .ZN(n89) );
  OAI22_X1 U706 ( .A1(n503), .A2(n350), .B1(n349), .B2(n532), .ZN(n275) );
  OAI22_X1 U707 ( .A1(n503), .A2(n346), .B1(n345), .B2(n532), .ZN(n271) );
  OAI22_X1 U708 ( .A1(n504), .A2(n347), .B1(n346), .B2(n532), .ZN(n272) );
  OAI22_X1 U709 ( .A1(n504), .A2(n348), .B1(n347), .B2(n532), .ZN(n273) );
  OAI22_X1 U710 ( .A1(n504), .A2(n349), .B1(n348), .B2(n532), .ZN(n274) );
  OAI22_X1 U711 ( .A1(n29), .A2(n612), .B1(n353), .B2(n532), .ZN(n254) );
  OAI22_X1 U712 ( .A1(n29), .A2(n351), .B1(n350), .B2(n532), .ZN(n276) );
  OAI22_X1 U713 ( .A1(n503), .A2(n352), .B1(n351), .B2(n532), .ZN(n277) );
  XOR2_X1 U714 ( .A(n56), .B(n556), .Z(product[5]) );
  XNOR2_X1 U715 ( .A(n88), .B(n51), .ZN(product[10]) );
  NOR2_X1 U716 ( .A1(n234), .A2(n257), .ZN(n113) );
  XNOR2_X1 U717 ( .A(n77), .B(n48), .ZN(product[13]) );
  NAND2_X1 U718 ( .A1(n224), .A2(n227), .ZN(n103) );
  OAI22_X1 U719 ( .A1(n552), .A2(n358), .B1(n357), .B2(n595), .ZN(n282) );
  OAI22_X1 U720 ( .A1(n551), .A2(n356), .B1(n355), .B2(n595), .ZN(n280) );
  OAI22_X1 U721 ( .A1(n552), .A2(n355), .B1(n354), .B2(n595), .ZN(n279) );
  OAI22_X1 U722 ( .A1(n551), .A2(n357), .B1(n356), .B2(n595), .ZN(n281) );
  OAI22_X1 U723 ( .A1(n551), .A2(n362), .B1(n361), .B2(n595), .ZN(n286) );
  OAI22_X1 U724 ( .A1(n551), .A2(n528), .B1(n364), .B2(n595), .ZN(n255) );
  OAI22_X1 U725 ( .A1(n552), .A2(n361), .B1(n360), .B2(n595), .ZN(n285) );
  OAI22_X1 U726 ( .A1(n552), .A2(n360), .B1(n359), .B2(n595), .ZN(n284) );
  OAI22_X1 U727 ( .A1(n23), .A2(n363), .B1(n362), .B2(n595), .ZN(n287) );
  XNOR2_X1 U728 ( .A(n548), .B(n424), .ZN(n375) );
  XNOR2_X1 U729 ( .A(n606), .B(n421), .ZN(n372) );
  XNOR2_X1 U730 ( .A(n548), .B(n423), .ZN(n374) );
  XNOR2_X1 U731 ( .A(n548), .B(n422), .ZN(n373) );
  OAI22_X1 U732 ( .A1(n359), .A2(n23), .B1(n358), .B2(n595), .ZN(n283) );
  XNOR2_X1 U733 ( .A(n501), .B(n419), .ZN(n370) );
  XNOR2_X1 U734 ( .A(n501), .B(n420), .ZN(n371) );
  INV_X1 U735 ( .A(n595), .ZN(n243) );
  OAI21_X1 U736 ( .B1(n87), .B2(n85), .A(n518), .ZN(n84) );
  OAI22_X1 U737 ( .A1(n511), .A2(n394), .B1(n393), .B2(n597), .ZN(n315) );
  OAI22_X1 U738 ( .A1(n511), .A2(n395), .B1(n394), .B2(n597), .ZN(n316) );
  OAI22_X1 U739 ( .A1(n511), .A2(n396), .B1(n395), .B2(n597), .ZN(n317) );
  OAI22_X1 U740 ( .A1(n511), .A2(n400), .B1(n399), .B2(n597), .ZN(n321) );
  OAI22_X1 U741 ( .A1(n401), .A2(n6), .B1(n400), .B2(n597), .ZN(n322) );
  OAI22_X1 U742 ( .A1(n511), .A2(n397), .B1(n396), .B2(n597), .ZN(n318) );
  OAI22_X1 U743 ( .A1(n511), .A2(n398), .B1(n397), .B2(n597), .ZN(n319) );
  OAI22_X1 U744 ( .A1(n6), .A2(n399), .B1(n398), .B2(n597), .ZN(n320) );
  OAI22_X1 U745 ( .A1(n402), .A2(n511), .B1(n513), .B2(n597), .ZN(n323) );
  OAI22_X1 U746 ( .A1(n6), .A2(n404), .B1(n403), .B2(n597), .ZN(n325) );
  OAI22_X1 U747 ( .A1(n511), .A2(n405), .B1(n404), .B2(n597), .ZN(n326) );
  OAI22_X1 U748 ( .A1(n511), .A2(n406), .B1(n405), .B2(n597), .ZN(n327) );
  OAI22_X1 U749 ( .A1(n511), .A2(n407), .B1(n406), .B2(n597), .ZN(n328) );
  OAI22_X1 U750 ( .A1(n511), .A2(n408), .B1(n407), .B2(n597), .ZN(n329) );
  OAI22_X1 U751 ( .A1(n511), .A2(n599), .B1(n409), .B2(n597), .ZN(n258) );
  AOI21_X1 U752 ( .B1(n104), .B2(n590), .A(n101), .ZN(n99) );
  XNOR2_X1 U753 ( .A(n84), .B(n50), .ZN(product[11]) );
  NAND2_X1 U754 ( .A1(n232), .A2(n233), .ZN(n111) );
  NAND2_X1 U755 ( .A1(n151), .A2(n139), .ZN(n62) );
  OAI22_X1 U756 ( .A1(n558), .A2(n370), .B1(n369), .B2(n529), .ZN(n293) );
  OAI22_X1 U757 ( .A1(n533), .A2(n367), .B1(n366), .B2(n529), .ZN(n290) );
  OAI22_X1 U758 ( .A1(n557), .A2(n368), .B1(n367), .B2(n529), .ZN(n291) );
  OAI22_X1 U759 ( .A1(n533), .A2(n375), .B1(n374), .B2(n529), .ZN(n298) );
  OAI22_X1 U760 ( .A1(n534), .A2(n372), .B1(n371), .B2(n529), .ZN(n295) );
  OAI22_X1 U761 ( .A1(n558), .A2(n373), .B1(n372), .B2(n529), .ZN(n296) );
  OAI22_X1 U762 ( .A1(n557), .A2(n371), .B1(n370), .B2(n529), .ZN(n294) );
  OAI22_X1 U763 ( .A1(n534), .A2(n374), .B1(n373), .B2(n596), .ZN(n297) );
  OAI22_X1 U764 ( .A1(n533), .A2(n369), .B1(n368), .B2(n529), .ZN(n292) );
  OAI22_X1 U765 ( .A1(n533), .A2(n376), .B1(n375), .B2(n529), .ZN(n299) );
  OAI22_X1 U766 ( .A1(n557), .A2(n535), .B1(n377), .B2(n529), .ZN(n256) );
  XNOR2_X1 U767 ( .A(n494), .B(n420), .ZN(n386) );
  OAI22_X1 U768 ( .A1(n558), .A2(n366), .B1(n365), .B2(n529), .ZN(n289) );
  INV_X1 U769 ( .A(n596), .ZN(n245) );
  XNOR2_X1 U770 ( .A(n494), .B(n421), .ZN(n387) );
  XNOR2_X1 U771 ( .A(n494), .B(n43), .ZN(n391) );
  XNOR2_X1 U772 ( .A(n494), .B(n422), .ZN(n388) );
  XNOR2_X1 U773 ( .A(n494), .B(n424), .ZN(n390) );
  XNOR2_X1 U774 ( .A(n604), .B(n423), .ZN(n389) );
  INV_X1 U775 ( .A(n568), .ZN(n87) );
  NAND2_X1 U776 ( .A1(n135), .A2(n114), .ZN(n58) );
  XNOR2_X1 U777 ( .A(n602), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U778 ( .A(n602), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U779 ( .A(n602), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U780 ( .A(n602), .B(n420), .ZN(n403) );
  XNOR2_X1 U781 ( .A(n598), .B(n419), .ZN(n402) );
  XNOR2_X1 U782 ( .A(n602), .B(n421), .ZN(n404) );
  XNOR2_X1 U783 ( .A(n598), .B(n422), .ZN(n405) );
  XNOR2_X1 U784 ( .A(n598), .B(n43), .ZN(n408) );
  XNOR2_X1 U785 ( .A(n602), .B(n423), .ZN(n406) );
  XNOR2_X1 U786 ( .A(n602), .B(n424), .ZN(n407) );
  OAI21_X1 U787 ( .B1(n64), .B2(n519), .A(n65), .ZN(n63) );
  XNOR2_X1 U788 ( .A(n70), .B(n47), .ZN(product[14]) );
  OAI21_X1 U789 ( .B1(n554), .B2(n78), .A(n79), .ZN(n77) );
  OAI21_X1 U790 ( .B1(n554), .B2(n71), .A(n72), .ZN(n70) );
  OAI22_X1 U791 ( .A1(n575), .A2(n379), .B1(n378), .B2(n578), .ZN(n301) );
  OAI22_X1 U792 ( .A1(n575), .A2(n380), .B1(n379), .B2(n578), .ZN(n302) );
  OAI22_X1 U793 ( .A1(n575), .A2(n385), .B1(n384), .B2(n579), .ZN(n307) );
  OAI22_X1 U794 ( .A1(n575), .A2(n537), .B1(n381), .B2(n579), .ZN(n304) );
  OAI22_X1 U795 ( .A1(n575), .A2(n381), .B1(n380), .B2(n579), .ZN(n303) );
  NAND2_X1 U796 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U797 ( .A1(n383), .A2(n576), .B1(n382), .B2(n579), .ZN(n305) );
  OAI22_X1 U798 ( .A1(n576), .A2(n384), .B1(n578), .B2(n383), .ZN(n306) );
  OAI22_X1 U799 ( .A1(n575), .A2(n386), .B1(n385), .B2(n578), .ZN(n308) );
  OAI22_X1 U800 ( .A1(n575), .A2(n387), .B1(n386), .B2(n578), .ZN(n309) );
  OAI22_X1 U801 ( .A1(n575), .A2(n569), .B1(n392), .B2(n579), .ZN(n257) );
  OAI22_X1 U802 ( .A1(n576), .A2(n389), .B1(n388), .B2(n579), .ZN(n311) );
  OAI22_X1 U803 ( .A1(n12), .A2(n388), .B1(n387), .B2(n578), .ZN(n310) );
  OAI22_X1 U804 ( .A1(n12), .A2(n390), .B1(n389), .B2(n579), .ZN(n312) );
  OAI22_X1 U805 ( .A1(n575), .A2(n391), .B1(n390), .B2(n579), .ZN(n313) );
  INV_X1 U806 ( .A(n608), .ZN(n607) );
  INV_X1 U807 ( .A(n31), .ZN(n613) );
  INV_X1 U808 ( .A(n615), .ZN(n614) );
  INV_X1 U809 ( .A(n36), .ZN(n615) );
  INV_X1 U810 ( .A(n617), .ZN(n616) );
  INV_X1 U811 ( .A(n40), .ZN(n617) );
  XOR2_X1 U812 ( .A(n259), .B(n251), .Z(n148) );
  XOR2_X1 U813 ( .A(n289), .B(n279), .Z(n146) );
  XOR2_X1 U814 ( .A(n149), .B(n147), .Z(n144) );
endmodule


module layer1_8_4_8_16_datapath_M8_N4_T16_P8_4_DW01_add_2 ( A, B, CI, SUM, CO
 );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n18,
         n19, n20, n21, n23, n25, n26, n28, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n48, n49, n51, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n71, n72, n73, n74,
         n75, n77, n79, n80, n81, n82, n83, n85, n87, n88, n90, n94, n95, n98,
         n99, n100, n102, n104, n161, n162, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177;

  INV_X1 U126 ( .A(n95), .ZN(n161) );
  NOR2_X2 U127 ( .A1(A[8]), .A2(B[8]), .ZN(n58) );
  NOR2_X1 U128 ( .A1(A[11]), .A2(B[11]), .ZN(n39) );
  AND2_X1 U129 ( .A1(A[13]), .A2(B[13]), .ZN(n162) );
  AND2_X1 U130 ( .A1(n169), .A2(n90), .ZN(SUM[0]) );
  OR2_X1 U131 ( .A1(A[15]), .A2(B[15]), .ZN(n164) );
  AOI21_X2 U132 ( .B1(n176), .B2(n72), .A(n69), .ZN(n67) );
  INV_X1 U133 ( .A(n166), .ZN(n48) );
  OR2_X2 U134 ( .A1(A[10]), .A2(B[10]), .ZN(n175) );
  XNOR2_X1 U135 ( .A(n41), .B(n165), .ZN(SUM[11]) );
  AND2_X1 U136 ( .A1(n95), .A2(n40), .ZN(n165) );
  AND2_X1 U137 ( .A1(A[10]), .A2(B[10]), .ZN(n166) );
  NOR2_X1 U138 ( .A1(A[13]), .A2(B[13]), .ZN(n167) );
  AOI21_X1 U139 ( .B1(n42), .B2(n34), .A(n35), .ZN(n168) );
  AOI21_X1 U140 ( .B1(n42), .B2(n34), .A(n35), .ZN(n33) );
  OR2_X1 U141 ( .A1(A[0]), .A2(B[0]), .ZN(n169) );
  INV_X1 U142 ( .A(n64), .ZN(n63) );
  INV_X1 U143 ( .A(n55), .ZN(n54) );
  AOI21_X1 U144 ( .B1(n175), .B2(n51), .A(n166), .ZN(n44) );
  AOI21_X1 U145 ( .B1(n171), .B2(n80), .A(n77), .ZN(n75) );
  INV_X1 U146 ( .A(n79), .ZN(n77) );
  AOI21_X1 U147 ( .B1(n172), .B2(n88), .A(n85), .ZN(n83) );
  INV_X1 U148 ( .A(n87), .ZN(n85) );
  OAI21_X1 U149 ( .B1(n83), .B2(n81), .A(n82), .ZN(n80) );
  INV_X1 U150 ( .A(n71), .ZN(n69) );
  OAI21_X1 U151 ( .B1(n75), .B2(n73), .A(n74), .ZN(n72) );
  AOI21_X1 U152 ( .B1(n56), .B2(n64), .A(n57), .ZN(n55) );
  AOI21_X1 U153 ( .B1(n54), .B2(n170), .A(n51), .ZN(n49) );
  INV_X1 U154 ( .A(n90), .ZN(n88) );
  OAI21_X1 U155 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  INV_X1 U156 ( .A(n53), .ZN(n51) );
  NAND2_X1 U157 ( .A1(n102), .A2(n74), .ZN(n12) );
  INV_X1 U158 ( .A(n73), .ZN(n102) );
  INV_X1 U159 ( .A(n39), .ZN(n95) );
  NAND2_X1 U160 ( .A1(n170), .A2(n53), .ZN(n7) );
  NAND2_X1 U161 ( .A1(n99), .A2(n62), .ZN(n9) );
  INV_X1 U162 ( .A(n61), .ZN(n99) );
  NAND2_X1 U163 ( .A1(n104), .A2(n82), .ZN(n14) );
  INV_X1 U164 ( .A(n81), .ZN(n104) );
  NAND2_X1 U165 ( .A1(n98), .A2(n59), .ZN(n8) );
  NAND2_X1 U166 ( .A1(n176), .A2(n71), .ZN(n11) );
  NAND2_X1 U167 ( .A1(n171), .A2(n79), .ZN(n13) );
  NAND2_X1 U168 ( .A1(n172), .A2(n87), .ZN(n15) );
  NAND2_X1 U169 ( .A1(n100), .A2(n66), .ZN(n10) );
  INV_X1 U170 ( .A(n65), .ZN(n100) );
  XNOR2_X1 U171 ( .A(n38), .B(n4), .ZN(SUM[12]) );
  XNOR2_X1 U172 ( .A(n54), .B(n7), .ZN(SUM[9]) );
  XOR2_X1 U173 ( .A(n63), .B(n9), .Z(SUM[7]) );
  XNOR2_X1 U174 ( .A(n11), .B(n72), .ZN(SUM[5]) );
  XOR2_X1 U175 ( .A(n12), .B(n75), .Z(SUM[4]) );
  XNOR2_X1 U176 ( .A(n13), .B(n80), .ZN(SUM[3]) );
  NOR2_X1 U177 ( .A1(A[7]), .A2(B[7]), .ZN(n61) );
  OR2_X1 U178 ( .A1(A[9]), .A2(B[9]), .ZN(n170) );
  NOR2_X1 U179 ( .A1(A[4]), .A2(B[4]), .ZN(n73) );
  NOR2_X1 U180 ( .A1(A[2]), .A2(B[2]), .ZN(n81) );
  XOR2_X1 U181 ( .A(n49), .B(n6), .Z(SUM[10]) );
  OR2_X1 U182 ( .A1(A[3]), .A2(B[3]), .ZN(n171) );
  OR2_X1 U183 ( .A1(A[1]), .A2(B[1]), .ZN(n172) );
  OR2_X1 U184 ( .A1(A[13]), .A2(B[13]), .ZN(n173) );
  OR2_X1 U185 ( .A1(A[14]), .A2(B[14]), .ZN(n174) );
  XNOR2_X1 U186 ( .A(n60), .B(n8), .ZN(SUM[8]) );
  NOR2_X1 U187 ( .A1(A[6]), .A2(B[6]), .ZN(n65) );
  NAND2_X1 U188 ( .A1(A[7]), .A2(B[7]), .ZN(n62) );
  OR2_X1 U189 ( .A1(A[5]), .A2(B[5]), .ZN(n176) );
  NAND2_X1 U190 ( .A1(A[4]), .A2(B[4]), .ZN(n74) );
  NAND2_X1 U191 ( .A1(A[2]), .A2(B[2]), .ZN(n82) );
  NAND2_X1 U192 ( .A1(A[5]), .A2(B[5]), .ZN(n71) );
  NAND2_X1 U193 ( .A1(A[1]), .A2(B[1]), .ZN(n87) );
  NAND2_X1 U194 ( .A1(A[3]), .A2(B[3]), .ZN(n79) );
  NAND2_X1 U195 ( .A1(A[0]), .A2(B[0]), .ZN(n90) );
  NAND2_X1 U196 ( .A1(A[6]), .A2(B[6]), .ZN(n66) );
  NAND2_X1 U197 ( .A1(A[8]), .A2(B[8]), .ZN(n59) );
  XOR2_X1 U198 ( .A(n14), .B(n83), .Z(SUM[2]) );
  XNOR2_X1 U199 ( .A(n15), .B(n88), .ZN(SUM[1]) );
  NAND2_X1 U200 ( .A1(n164), .A2(n18), .ZN(n1) );
  NOR2_X1 U201 ( .A1(A[12]), .A2(B[12]), .ZN(n177) );
  NOR2_X1 U202 ( .A1(A[12]), .A2(B[12]), .ZN(n36) );
  NAND2_X1 U203 ( .A1(A[12]), .A2(B[12]), .ZN(n37) );
  NAND2_X1 U204 ( .A1(n37), .A2(n94), .ZN(n4) );
  INV_X1 U205 ( .A(n25), .ZN(n23) );
  INV_X1 U206 ( .A(n58), .ZN(n98) );
  NOR2_X1 U207 ( .A1(n58), .A2(n61), .ZN(n56) );
  OAI21_X1 U208 ( .B1(n58), .B2(n62), .A(n59), .ZN(n57) );
  NAND2_X1 U209 ( .A1(A[9]), .A2(B[9]), .ZN(n53) );
  NAND2_X1 U210 ( .A1(n173), .A2(n28), .ZN(n3) );
  NAND2_X1 U211 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  NAND2_X1 U212 ( .A1(A[11]), .A2(B[11]), .ZN(n40) );
  NAND2_X1 U213 ( .A1(A[14]), .A2(B[14]), .ZN(n25) );
  XOR2_X1 U214 ( .A(n10), .B(n67), .Z(SUM[6]) );
  OAI21_X1 U215 ( .B1(n67), .B2(n65), .A(n66), .ZN(n64) );
  INV_X1 U216 ( .A(n177), .ZN(n94) );
  NOR2_X1 U217 ( .A1(n177), .A2(n39), .ZN(n34) );
  OAI21_X1 U218 ( .B1(n36), .B2(n40), .A(n37), .ZN(n35) );
  NAND2_X1 U219 ( .A1(A[15]), .A2(B[15]), .ZN(n18) );
  OAI21_X1 U220 ( .B1(n41), .B2(n161), .A(n40), .ZN(n38) );
  INV_X1 U221 ( .A(n42), .ZN(n41) );
  OAI21_X1 U222 ( .B1(n43), .B2(n55), .A(n44), .ZN(n42) );
  NAND2_X1 U223 ( .A1(n174), .A2(n25), .ZN(n2) );
  NAND2_X1 U224 ( .A1(n174), .A2(n173), .ZN(n20) );
  AOI21_X1 U225 ( .B1(n174), .B2(n162), .A(n23), .ZN(n21) );
  XNOR2_X1 U226 ( .A(n19), .B(n1), .ZN(SUM[15]) );
  NAND2_X1 U227 ( .A1(n175), .A2(n48), .ZN(n6) );
  NAND2_X1 U228 ( .A1(n175), .A2(n170), .ZN(n43) );
  XNOR2_X1 U229 ( .A(n26), .B(n2), .ZN(SUM[14]) );
  XOR2_X1 U230 ( .A(n168), .B(n3), .Z(SUM[13]) );
  OAI21_X1 U231 ( .B1(n33), .B2(n167), .A(n28), .ZN(n26) );
  OAI21_X1 U232 ( .B1(n168), .B2(n20), .A(n21), .ZN(n19) );
endmodule


module layer1_8_4_8_16_datapath_M8_N4_T16_P8_4 ( clk, clear_acc, data_out_x, 
        data_out, data_out_w, data_out_b, wr_en_y, m_valid, m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [3:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N27, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, n1, n2, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n87, n104, n113, n114, n115, n116, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n8), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n217), .CK(clk), .Q(n13) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n218), .CK(clk), .Q(n14) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n219), .CK(clk), .Q(n15) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n220), .CK(clk), .Q(n16) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n221), .CK(clk), .Q(n17) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n222), .CK(clk), .Q(n18) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n223), .CK(clk), .Q(n19) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n224), .CK(clk), .Q(n20) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n225), .CK(clk), .Q(n21) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n226), .CK(clk), .Q(n22) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n227), .CK(clk), .Q(n23) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n228), .CK(clk), .Q(n24) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n229), .CK(clk), .Q(n25) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n230), .CK(clk), .Q(n26) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n231), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n232), .CK(clk), .Q(n29) );
  DFF_X1 \f_reg[0]  ( .D(n85), .CK(clk), .Q(n56), .QN(n206) );
  DFF_X1 \f_reg[1]  ( .D(n84), .CK(clk), .Q(n54), .QN(n207) );
  DFF_X1 \f_reg[2]  ( .D(n83), .CK(clk), .Q(n52), .QN(n208) );
  DFF_X1 \f_reg[3]  ( .D(n82), .CK(clk), .Q(f[3]), .QN(n60) );
  DFF_X1 \f_reg[4]  ( .D(n81), .CK(clk), .Q(f[4]), .QN(n61) );
  DFF_X1 \f_reg[5]  ( .D(n80), .CK(clk), .Q(f[5]), .QN(n62) );
  DFF_X1 \f_reg[6]  ( .D(n79), .CK(clk), .Q(f[6]), .QN(n63) );
  DFF_X1 \f_reg[7]  ( .D(n78), .CK(clk), .Q(f[7]), .QN(n209) );
  DFF_X1 \f_reg[8]  ( .D(n77), .CK(clk), .Q(f[8]), .QN(n210) );
  DFF_X1 \f_reg[9]  ( .D(n76), .CK(clk), .Q(f[9]), .QN(n211) );
  DFF_X1 \f_reg[10]  ( .D(n75), .CK(clk), .Q(n44), .QN(n212) );
  DFF_X1 \f_reg[11]  ( .D(n74), .CK(clk), .Q(n42), .QN(n213) );
  DFF_X1 \f_reg[12]  ( .D(n73), .CK(clk), .Q(n40), .QN(n214) );
  DFF_X1 \f_reg[13]  ( .D(n72), .CK(clk), .Q(n38), .QN(n215) );
  DFF_X1 \f_reg[14]  ( .D(n71), .CK(clk), .Q(n36), .QN(n216) );
  DFF_X1 \f_reg[15]  ( .D(n70), .CK(clk), .Q(f[15]), .QN(n68) );
  DFF_X1 \data_out_reg[15]  ( .D(n104), .CK(clk), .Q(data_out[15]), .QN(n189)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n113), .CK(clk), .Q(data_out[14]), .QN(n188)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n114), .CK(clk), .Q(data_out[13]), .QN(n187)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n115), .CK(clk), .Q(data_out[12]), .QN(n186)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n116), .CK(clk), .Q(data_out[11]), .QN(n185)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n163), .CK(clk), .Q(data_out[10]), .QN(n184)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n164), .CK(clk), .Q(data_out[9]), .QN(n183) );
  DFF_X1 \data_out_reg[8]  ( .D(n165), .CK(clk), .Q(data_out[8]), .QN(n182) );
  DFF_X1 \data_out_reg[7]  ( .D(n166), .CK(clk), .Q(data_out[7]), .QN(n181) );
  DFF_X1 \data_out_reg[6]  ( .D(n167), .CK(clk), .Q(data_out[6]), .QN(n180) );
  DFF_X1 \data_out_reg[5]  ( .D(n168), .CK(clk), .Q(data_out[5]), .QN(n179) );
  DFF_X1 \data_out_reg[4]  ( .D(n169), .CK(clk), .Q(data_out[4]), .QN(n178) );
  DFF_X1 \data_out_reg[3]  ( .D(n170), .CK(clk), .Q(data_out[3]), .QN(n177) );
  DFF_X1 \data_out_reg[2]  ( .D(n171), .CK(clk), .Q(data_out[2]), .QN(n176) );
  DFF_X1 \data_out_reg[1]  ( .D(n172), .CK(clk), .Q(data_out[1]), .QN(n175) );
  DFF_X1 \data_out_reg[0]  ( .D(n173), .CK(clk), .Q(data_out[0]), .QN(n174) );
  layer1_8_4_8_16_datapath_M8_N4_T16_P8_4_DW_mult_tc_1 mult_183 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer1_8_4_8_16_datapath_M8_N4_T16_P8_4_DW01_add_2 add_184 ( .A({n196, n195, 
        n194, n193, n192, n191, n205, n204, n203, n202, n201, n200, n199, n198, 
        n197, n190}), .B({f[15], n36, n38, n40, n42, n44, f[9:3], n52, n54, 
        n56}), .CI(1'b0), .SUM(adder) );
  DFF_X2 delay_reg ( .D(N27), .CK(clk), .Q(n6), .QN(n233) );
  CLKBUF_X1 U3 ( .A(N39), .Z(n1) );
  MUX2_X2 U4 ( .A(n20), .B(N37), .S(n233), .Z(n204) );
  AND2_X1 U5 ( .A1(n58), .A2(f[15]), .ZN(n2) );
  AND2_X1 U6 ( .A1(data_out_b[15]), .A2(n8), .ZN(n4) );
  MUX2_X1 U8 ( .A(N43), .B(n14), .S(n6), .Z(n195) );
  MUX2_X2 U9 ( .A(N39), .B(n18), .S(n6), .Z(n191) );
  MUX2_X2 U10 ( .A(n15), .B(N42), .S(n233), .Z(n194) );
  CLKBUF_X1 U11 ( .A(N41), .Z(n5) );
  AOI211_X1 U12 ( .C1(adder[15]), .C2(n7), .A(n2), .B(n4), .ZN(n35) );
  MUX2_X2 U13 ( .A(n17), .B(N40), .S(n233), .Z(n192) );
  AND2_X2 U14 ( .A1(n34), .A2(n9), .ZN(n7) );
  MUX2_X2 U15 ( .A(n16), .B(N41), .S(n233), .Z(n193) );
  INV_X1 U16 ( .A(n9), .ZN(n8) );
  INV_X1 U17 ( .A(n34), .ZN(n58) );
  INV_X1 U18 ( .A(clear_acc), .ZN(n9) );
  NAND2_X1 U19 ( .A1(n87), .A2(N27), .ZN(n235) );
  INV_X1 U20 ( .A(wr_en_y), .ZN(n87) );
  OAI22_X1 U21 ( .A1(n177), .A2(n235), .B1(n60), .B2(n234), .ZN(n170) );
  OAI22_X1 U22 ( .A1(n178), .A2(n235), .B1(n61), .B2(n234), .ZN(n169) );
  OAI22_X1 U23 ( .A1(n179), .A2(n235), .B1(n62), .B2(n234), .ZN(n168) );
  OAI22_X1 U24 ( .A1(n180), .A2(n235), .B1(n63), .B2(n234), .ZN(n167) );
  OAI22_X1 U25 ( .A1(n181), .A2(n235), .B1(n209), .B2(n234), .ZN(n166) );
  OAI22_X1 U26 ( .A1(n182), .A2(n235), .B1(n210), .B2(n234), .ZN(n165) );
  OAI22_X1 U27 ( .A1(n183), .A2(n235), .B1(n211), .B2(n234), .ZN(n164) );
  INV_X1 U28 ( .A(n12), .ZN(n28) );
  AND3_X1 U29 ( .A1(sel[1]), .A2(sel[2]), .A3(sel[0]), .ZN(n11) );
  INV_X1 U30 ( .A(m_ready), .ZN(n10) );
  NAND2_X1 U31 ( .A1(m_valid), .A2(n10), .ZN(n32) );
  OAI21_X1 U32 ( .B1(sel[3]), .B2(n11), .A(n32), .ZN(N27) );
  NAND2_X1 U33 ( .A1(clear_acc_delay), .A2(n233), .ZN(n12) );
  MUX2_X1 U34 ( .A(n13), .B(N44), .S(n28), .Z(n217) );
  MUX2_X1 U35 ( .A(n13), .B(N44), .S(n233), .Z(n196) );
  MUX2_X1 U36 ( .A(n14), .B(N43), .S(n28), .Z(n218) );
  MUX2_X1 U37 ( .A(n15), .B(N42), .S(n28), .Z(n219) );
  MUX2_X1 U38 ( .A(n16), .B(n5), .S(n28), .Z(n220) );
  MUX2_X1 U39 ( .A(n17), .B(N40), .S(n28), .Z(n221) );
  MUX2_X1 U40 ( .A(n18), .B(n1), .S(n28), .Z(n222) );
  MUX2_X1 U41 ( .A(n19), .B(N38), .S(n28), .Z(n223) );
  MUX2_X1 U42 ( .A(n19), .B(N38), .S(n233), .Z(n205) );
  MUX2_X1 U43 ( .A(n20), .B(N37), .S(n28), .Z(n224) );
  MUX2_X1 U44 ( .A(n21), .B(N36), .S(n28), .Z(n225) );
  MUX2_X1 U45 ( .A(n21), .B(N36), .S(n233), .Z(n203) );
  MUX2_X1 U46 ( .A(n22), .B(N35), .S(n28), .Z(n226) );
  MUX2_X1 U47 ( .A(n22), .B(N35), .S(n233), .Z(n202) );
  MUX2_X1 U48 ( .A(n23), .B(N34), .S(n28), .Z(n227) );
  MUX2_X1 U49 ( .A(n23), .B(N34), .S(n233), .Z(n201) );
  MUX2_X1 U50 ( .A(n24), .B(N33), .S(n28), .Z(n228) );
  MUX2_X1 U51 ( .A(n24), .B(N33), .S(n233), .Z(n200) );
  MUX2_X1 U52 ( .A(n25), .B(N32), .S(n28), .Z(n229) );
  MUX2_X1 U53 ( .A(n25), .B(N32), .S(n233), .Z(n199) );
  MUX2_X1 U54 ( .A(n26), .B(N31), .S(n28), .Z(n230) );
  MUX2_X1 U55 ( .A(n26), .B(N31), .S(n233), .Z(n198) );
  MUX2_X1 U56 ( .A(n27), .B(N30), .S(n28), .Z(n231) );
  MUX2_X1 U57 ( .A(n27), .B(N30), .S(n233), .Z(n197) );
  MUX2_X1 U58 ( .A(n29), .B(N29), .S(n28), .Z(n232) );
  MUX2_X1 U59 ( .A(n29), .B(N29), .S(n233), .Z(n190) );
  INV_X1 U60 ( .A(n32), .ZN(n33) );
  OAI21_X1 U61 ( .B1(n33), .B2(n6), .A(n9), .ZN(n34) );
  INV_X1 U62 ( .A(n35), .ZN(n70) );
  AOI222_X1 U63 ( .A1(data_out_b[14]), .A2(n8), .B1(adder[14]), .B2(n7), .C1(
        n58), .C2(n36), .ZN(n37) );
  INV_X1 U64 ( .A(n37), .ZN(n71) );
  AOI222_X1 U65 ( .A1(data_out_b[13]), .A2(n8), .B1(adder[13]), .B2(n7), .C1(
        n58), .C2(n38), .ZN(n39) );
  INV_X1 U66 ( .A(n39), .ZN(n72) );
  AOI222_X1 U67 ( .A1(data_out_b[12]), .A2(n8), .B1(adder[12]), .B2(n7), .C1(
        n58), .C2(n40), .ZN(n41) );
  INV_X1 U68 ( .A(n41), .ZN(n73) );
  AOI222_X1 U69 ( .A1(data_out_b[11]), .A2(n8), .B1(adder[11]), .B2(n7), .C1(
        n58), .C2(n42), .ZN(n43) );
  INV_X1 U70 ( .A(n43), .ZN(n74) );
  AOI222_X1 U71 ( .A1(data_out_b[10]), .A2(n8), .B1(adder[10]), .B2(n7), .C1(
        n58), .C2(n44), .ZN(n45) );
  INV_X1 U72 ( .A(n45), .ZN(n75) );
  AOI222_X1 U73 ( .A1(data_out_b[8]), .A2(n8), .B1(adder[8]), .B2(n7), .C1(n58), .C2(f[8]), .ZN(n46) );
  INV_X1 U74 ( .A(n46), .ZN(n77) );
  AOI222_X1 U75 ( .A1(data_out_b[7]), .A2(n8), .B1(adder[7]), .B2(n7), .C1(n58), .C2(f[7]), .ZN(n47) );
  INV_X1 U76 ( .A(n47), .ZN(n78) );
  AOI222_X1 U77 ( .A1(data_out_b[6]), .A2(n8), .B1(adder[6]), .B2(n7), .C1(n58), .C2(f[6]), .ZN(n48) );
  INV_X1 U78 ( .A(n48), .ZN(n79) );
  AOI222_X1 U79 ( .A1(data_out_b[5]), .A2(n8), .B1(adder[5]), .B2(n7), .C1(n58), .C2(f[5]), .ZN(n49) );
  INV_X1 U80 ( .A(n49), .ZN(n80) );
  AOI222_X1 U81 ( .A1(data_out_b[4]), .A2(n8), .B1(adder[4]), .B2(n7), .C1(n58), .C2(f[4]), .ZN(n50) );
  INV_X1 U82 ( .A(n50), .ZN(n81) );
  AOI222_X1 U83 ( .A1(data_out_b[3]), .A2(n8), .B1(adder[3]), .B2(n7), .C1(n58), .C2(f[3]), .ZN(n51) );
  INV_X1 U84 ( .A(n51), .ZN(n82) );
  AOI222_X1 U85 ( .A1(data_out_b[2]), .A2(n8), .B1(adder[2]), .B2(n7), .C1(n58), .C2(n52), .ZN(n53) );
  INV_X1 U86 ( .A(n53), .ZN(n83) );
  AOI222_X1 U87 ( .A1(data_out_b[1]), .A2(n8), .B1(adder[1]), .B2(n7), .C1(n58), .C2(n54), .ZN(n55) );
  INV_X1 U88 ( .A(n55), .ZN(n84) );
  AOI222_X1 U89 ( .A1(data_out_b[0]), .A2(n8), .B1(adder[0]), .B2(n7), .C1(n58), .C2(n56), .ZN(n57) );
  INV_X1 U90 ( .A(n57), .ZN(n85) );
  AOI222_X1 U91 ( .A1(data_out_b[9]), .A2(n8), .B1(adder[9]), .B2(n7), .C1(n58), .C2(f[9]), .ZN(n59) );
  INV_X1 U92 ( .A(n59), .ZN(n76) );
  NOR4_X1 U93 ( .A1(n42), .A2(n40), .A3(n38), .A4(n36), .ZN(n67) );
  NOR4_X1 U94 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n44), .ZN(n66) );
  NAND4_X1 U95 ( .A1(n63), .A2(n62), .A3(n61), .A4(n60), .ZN(n64) );
  NOR4_X1 U96 ( .A1(n64), .A2(n56), .A3(n54), .A4(n52), .ZN(n65) );
  NAND3_X1 U97 ( .A1(n67), .A2(n66), .A3(n65), .ZN(n69) );
  NAND3_X1 U98 ( .A1(wr_en_y), .A2(n69), .A3(n68), .ZN(n234) );
  OAI22_X1 U99 ( .A1(n174), .A2(n235), .B1(n206), .B2(n234), .ZN(n173) );
  OAI22_X1 U100 ( .A1(n175), .A2(n235), .B1(n207), .B2(n234), .ZN(n172) );
  OAI22_X1 U101 ( .A1(n176), .A2(n235), .B1(n208), .B2(n234), .ZN(n171) );
  OAI22_X1 U102 ( .A1(n184), .A2(n235), .B1(n212), .B2(n234), .ZN(n163) );
  OAI22_X1 U103 ( .A1(n185), .A2(n235), .B1(n213), .B2(n234), .ZN(n116) );
  OAI22_X1 U104 ( .A1(n186), .A2(n235), .B1(n214), .B2(n234), .ZN(n115) );
  OAI22_X1 U105 ( .A1(n187), .A2(n235), .B1(n215), .B2(n234), .ZN(n114) );
  OAI22_X1 U106 ( .A1(n188), .A2(n235), .B1(n216), .B2(n234), .ZN(n113) );
  OAI22_X1 U107 ( .A1(n189), .A2(n235), .B1(n68), .B2(n234), .ZN(n104) );
endmodule


module layer1_8_4_8_16_datapath_M8_N4_T16_P8_3_DW_mult_tc_1 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n9, n12, n13, n16, n18, n19, n21, n23, n25, n27, n29, n31,
         n32, n34, n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n50,
         n53, n54, n55, n56, n57, n58, n59, n62, n63, n64, n65, n67, n69, n70,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n89, n90, n91, n93, n95, n96, n97, n98, n99, n101, n103,
         n104, n105, n106, n107, n109, n111, n112, n113, n114, n115, n117,
         n119, n120, n122, n125, n127, n128, n135, n139, n141, n142, n143,
         n144, n145, n146, n148, n149, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n237, n245, n247, n249, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n418, n419, n420, n421, n422, n423, n424, n426, n427, n429, n430,
         n433, n490, n491, n492, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U148 ( .A(n265), .B(n144), .Z(n145) );
  XOR2_X1 U152 ( .A(n301), .B(n148), .Z(n149) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U162 ( .A(n170), .B(n172), .CI(n179), .CO(n165), .S(n166) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n263), .CI(n291), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n252), .B(n317), .CO(n173), .S(n174) );
  FA_X1 U167 ( .A(n180), .B(n187), .CI(n178), .CO(n175), .S(n176) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U169 ( .A(n193), .B(n282), .CI(n191), .CO(n179), .S(n180) );
  FA_X1 U170 ( .A(n268), .B(n274), .CI(n292), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U172 ( .A(n197), .B(n190), .CI(n188), .CO(n185), .S(n186) );
  FA_X1 U173 ( .A(n199), .B(n201), .CI(n192), .CO(n187), .S(n188) );
  FA_X1 U174 ( .A(n275), .B(n293), .CI(n194), .CO(n189), .S(n190) );
  FA_X1 U175 ( .A(n305), .B(n253), .CI(n283), .CO(n191), .S(n192) );
  HA_X1 U176 ( .A(n269), .B(n319), .CO(n193), .S(n194) );
  FA_X1 U177 ( .A(n205), .B(n200), .CI(n198), .CO(n195), .S(n196) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U180 ( .A(n320), .B(n270), .CI(n306), .CO(n201), .S(n202) );
  FA_X1 U181 ( .A(n208), .B(n213), .CI(n206), .CO(n203), .S(n204) );
  FA_X1 U182 ( .A(n215), .B(n307), .CI(n210), .CO(n205), .S(n206) );
  FA_X1 U183 ( .A(n285), .B(n254), .CI(n295), .CO(n207), .S(n208) );
  HA_X1 U184 ( .A(n321), .B(n277), .CO(n209), .S(n210) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n308), .B(n278), .CI(n322), .CO(n215), .S(n216) );
  FA_X1 U188 ( .A(n225), .B(n222), .CI(n220), .CO(n217), .S(n218) );
  FA_X1 U189 ( .A(n255), .B(n309), .CI(n297), .CO(n219), .S(n220) );
  HA_X1 U190 ( .A(n323), .B(n287), .CO(n221), .S(n222) );
  FA_X1 U192 ( .A(n324), .B(n288), .CI(n310), .CO(n225), .S(n226) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  HA_X1 U194 ( .A(n325), .B(n311), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n326), .B(n300), .CI(n312), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  BUF_X1 U414 ( .A(n107), .Z(n490) );
  BUF_X2 U415 ( .A(n12), .Z(n537) );
  XOR2_X1 U416 ( .A(n590), .B(a[6]), .Z(n491) );
  NAND2_X1 U417 ( .A1(n429), .A2(n27), .ZN(n29) );
  BUF_X2 U418 ( .A(n16), .Z(n580) );
  INV_X2 U419 ( .A(n249), .ZN(n582) );
  OR2_X1 U420 ( .A1(n212), .A2(n217), .ZN(n492) );
  BUF_X1 U421 ( .A(n27), .Z(n544) );
  BUF_X1 U422 ( .A(n587), .Z(n518) );
  AND2_X1 U423 ( .A1(n569), .A2(n122), .ZN(product[1]) );
  CLKBUF_X1 U424 ( .A(n85), .Z(n494) );
  XNOR2_X1 U425 ( .A(n592), .B(a[4]), .ZN(n571) );
  XNOR2_X1 U426 ( .A(n214), .B(n495), .ZN(n212) );
  XNOR2_X1 U427 ( .A(n216), .B(n219), .ZN(n495) );
  CLKBUF_X3 U428 ( .A(n498), .Z(n496) );
  CLKBUF_X1 U429 ( .A(n498), .Z(n581) );
  BUF_X1 U430 ( .A(n533), .Z(n497) );
  XNOR2_X1 U431 ( .A(n585), .B(a[2]), .ZN(n498) );
  CLKBUF_X1 U432 ( .A(n23), .Z(n499) );
  OAI21_X1 U433 ( .B1(n75), .B2(n79), .A(n76), .ZN(n500) );
  INV_X1 U434 ( .A(n542), .ZN(n501) );
  OAI21_X1 U435 ( .B1(n545), .B2(n501), .A(n90), .ZN(n502) );
  OR2_X1 U436 ( .A1(n541), .A2(n78), .ZN(n503) );
  XNOR2_X1 U437 ( .A(n166), .B(n504), .ZN(n164) );
  XNOR2_X1 U438 ( .A(n177), .B(n168), .ZN(n504) );
  CLKBUF_X1 U439 ( .A(n79), .Z(n505) );
  XNOR2_X1 U440 ( .A(n545), .B(n506), .ZN(product[9]) );
  AND2_X1 U441 ( .A1(n542), .A2(n90), .ZN(n506) );
  OR2_X1 U442 ( .A1(n218), .A2(n223), .ZN(n507) );
  XNOR2_X1 U443 ( .A(n45), .B(n508), .ZN(product[12]) );
  AND2_X1 U444 ( .A1(n540), .A2(n79), .ZN(n508) );
  BUF_X2 U445 ( .A(n12), .Z(n538) );
  XNOR2_X1 U446 ( .A(n226), .B(n509), .ZN(n224) );
  XNOR2_X1 U447 ( .A(n229), .B(n298), .ZN(n509) );
  CLKBUF_X1 U448 ( .A(n104), .Z(n510) );
  OAI21_X1 U449 ( .B1(n91), .B2(n89), .A(n90), .ZN(n511) );
  NOR2_X1 U450 ( .A1(n186), .A2(n195), .ZN(n512) );
  NOR2_X1 U451 ( .A1(n186), .A2(n195), .ZN(n82) );
  BUF_X1 U452 ( .A(n37), .Z(n513) );
  CLKBUF_X1 U453 ( .A(n568), .Z(n514) );
  CLKBUF_X1 U454 ( .A(n568), .Z(n515) );
  NOR2_X1 U455 ( .A1(n196), .A2(n203), .ZN(n85) );
  INV_X1 U456 ( .A(n85), .ZN(n128) );
  CLKBUF_X1 U457 ( .A(n45), .Z(n548) );
  OAI21_X1 U458 ( .B1(n512), .B2(n86), .A(n83), .ZN(n516) );
  OR2_X1 U459 ( .A1(n228), .A2(n231), .ZN(n517) );
  XNOR2_X2 U460 ( .A(n590), .B(a[6]), .ZN(n568) );
  XOR2_X1 U461 ( .A(n294), .B(n276), .Z(n519) );
  XOR2_X1 U462 ( .A(n519), .B(n284), .Z(n200) );
  NAND2_X1 U463 ( .A1(n284), .A2(n294), .ZN(n520) );
  NAND2_X1 U464 ( .A1(n284), .A2(n276), .ZN(n521) );
  NAND2_X1 U465 ( .A1(n294), .A2(n276), .ZN(n522) );
  NAND3_X1 U466 ( .A1(n520), .A2(n521), .A3(n522), .ZN(n199) );
  NAND2_X1 U467 ( .A1(n166), .A2(n177), .ZN(n523) );
  NAND2_X1 U468 ( .A1(n166), .A2(n168), .ZN(n524) );
  NAND2_X1 U469 ( .A1(n177), .A2(n168), .ZN(n525) );
  NAND3_X1 U470 ( .A1(n523), .A2(n524), .A3(n525), .ZN(n163) );
  OR2_X2 U471 ( .A1(n152), .A2(n163), .ZN(n572) );
  CLKBUF_X3 U472 ( .A(n19), .Z(n557) );
  XNOR2_X1 U473 ( .A(n593), .B(a[6]), .ZN(n430) );
  INV_X1 U474 ( .A(n497), .ZN(n526) );
  XNOR2_X1 U475 ( .A(n589), .B(a[2]), .ZN(n570) );
  CLKBUF_X1 U476 ( .A(n568), .Z(n527) );
  INV_X2 U477 ( .A(n589), .ZN(n554) );
  XNOR2_X1 U478 ( .A(n595), .B(a[8]), .ZN(n429) );
  BUF_X1 U479 ( .A(n587), .Z(n528) );
  INV_X1 U480 ( .A(n27), .ZN(n529) );
  INV_X1 U481 ( .A(n529), .ZN(n530) );
  INV_X1 U482 ( .A(n597), .ZN(n531) );
  INV_X1 U483 ( .A(n597), .ZN(n532) );
  INV_X1 U484 ( .A(n597), .ZN(n596) );
  BUF_X1 U485 ( .A(n12), .Z(n536) );
  INV_X1 U486 ( .A(n592), .ZN(n533) );
  NAND2_X1 U487 ( .A1(n571), .A2(n555), .ZN(n534) );
  NAND2_X1 U488 ( .A1(n571), .A2(n555), .ZN(n18) );
  XNOR2_X1 U489 ( .A(n528), .B(n249), .ZN(n433) );
  CLKBUF_X1 U490 ( .A(n16), .Z(n555) );
  INV_X1 U491 ( .A(n595), .ZN(n535) );
  INV_X1 U492 ( .A(n595), .ZN(n594) );
  NAND2_X1 U493 ( .A1(n9), .A2(n570), .ZN(n12) );
  XNOR2_X1 U494 ( .A(n149), .B(n539), .ZN(n144) );
  XNOR2_X1 U495 ( .A(n146), .B(n271), .ZN(n539) );
  OR2_X1 U496 ( .A1(n185), .A2(n176), .ZN(n540) );
  NOR2_X1 U497 ( .A1(n164), .A2(n175), .ZN(n541) );
  NOR2_X1 U498 ( .A1(n164), .A2(n175), .ZN(n75) );
  OR2_X1 U499 ( .A1(n204), .A2(n211), .ZN(n542) );
  OR2_X2 U500 ( .A1(n563), .A2(n543), .ZN(n34) );
  XNOR2_X1 U501 ( .A(n596), .B(a[10]), .ZN(n543) );
  INV_X1 U502 ( .A(n563), .ZN(n32) );
  AOI21_X1 U503 ( .B1(n96), .B2(n492), .A(n93), .ZN(n545) );
  AOI21_X1 U504 ( .B1(n96), .B2(n492), .A(n93), .ZN(n91) );
  CLKBUF_X1 U505 ( .A(n99), .Z(n546) );
  OAI21_X1 U506 ( .B1(n91), .B2(n89), .A(n90), .ZN(n547) );
  XNOR2_X1 U507 ( .A(n502), .B(n549), .ZN(product[10]) );
  NAND2_X1 U508 ( .A1(n128), .A2(n86), .ZN(n549) );
  NAND2_X1 U509 ( .A1(n214), .A2(n216), .ZN(n550) );
  NAND2_X1 U510 ( .A1(n214), .A2(n219), .ZN(n551) );
  NAND2_X1 U511 ( .A1(n216), .A2(n219), .ZN(n552) );
  NAND3_X1 U512 ( .A1(n550), .A2(n551), .A3(n552), .ZN(n211) );
  NAND2_X1 U513 ( .A1(n21), .A2(n430), .ZN(n553) );
  NAND2_X1 U514 ( .A1(n21), .A2(n430), .ZN(n23) );
  INV_X1 U515 ( .A(n564), .ZN(n27) );
  AOI21_X1 U516 ( .B1(n80), .B2(n511), .A(n81), .ZN(n567) );
  INV_X1 U517 ( .A(n589), .ZN(n588) );
  INV_X1 U518 ( .A(n592), .ZN(n590) );
  INV_X2 U519 ( .A(n592), .ZN(n591) );
  INV_X1 U520 ( .A(n554), .ZN(n556) );
  NAND2_X1 U521 ( .A1(n433), .A2(n582), .ZN(n558) );
  NAND2_X1 U522 ( .A1(n433), .A2(n582), .ZN(n559) );
  NAND2_X1 U523 ( .A1(n433), .A2(n582), .ZN(n6) );
  XOR2_X1 U524 ( .A(n589), .B(a[4]), .Z(n16) );
  NAND2_X1 U525 ( .A1(n226), .A2(n229), .ZN(n560) );
  NAND2_X1 U526 ( .A1(n226), .A2(n298), .ZN(n561) );
  NAND2_X1 U527 ( .A1(n229), .A2(n298), .ZN(n562) );
  NAND3_X1 U528 ( .A1(n560), .A2(n561), .A3(n562), .ZN(n223) );
  XNOR2_X1 U529 ( .A(n595), .B(a[10]), .ZN(n563) );
  XNOR2_X1 U530 ( .A(n593), .B(a[8]), .ZN(n564) );
  INV_X1 U531 ( .A(n518), .ZN(n565) );
  INV_X1 U532 ( .A(n528), .ZN(n566) );
  INV_X1 U533 ( .A(n587), .ZN(n585) );
  XNOR2_X1 U534 ( .A(n533), .B(a[6]), .ZN(n21) );
  NAND2_X1 U535 ( .A1(n176), .A2(n185), .ZN(n79) );
  OR2_X1 U536 ( .A1(n224), .A2(n227), .ZN(n574) );
  OR2_X1 U537 ( .A1(n329), .A2(n258), .ZN(n569) );
  NAND2_X1 U538 ( .A1(n572), .A2(n69), .ZN(n47) );
  AOI21_X1 U539 ( .B1(n500), .B2(n572), .A(n67), .ZN(n65) );
  INV_X1 U540 ( .A(n69), .ZN(n67) );
  INV_X1 U541 ( .A(n74), .ZN(n72) );
  INV_X1 U542 ( .A(n95), .ZN(n93) );
  NAND2_X1 U543 ( .A1(n125), .A2(n76), .ZN(n48) );
  INV_X1 U544 ( .A(n541), .ZN(n125) );
  NAND2_X1 U545 ( .A1(n492), .A2(n95), .ZN(n53) );
  OAI21_X1 U546 ( .B1(n75), .B2(n79), .A(n76), .ZN(n74) );
  NOR2_X1 U547 ( .A1(n541), .A2(n78), .ZN(n73) );
  XNOR2_X1 U548 ( .A(n84), .B(n50), .ZN(product[11]) );
  NAND2_X1 U549 ( .A1(n127), .A2(n83), .ZN(n50) );
  NAND2_X1 U550 ( .A1(n152), .A2(n163), .ZN(n69) );
  INV_X1 U551 ( .A(n113), .ZN(n135) );
  NAND2_X1 U552 ( .A1(n507), .A2(n98), .ZN(n54) );
  NOR2_X1 U553 ( .A1(n176), .A2(n185), .ZN(n78) );
  NAND2_X1 U554 ( .A1(n574), .A2(n103), .ZN(n55) );
  OAI21_X1 U555 ( .B1(n113), .B2(n115), .A(n114), .ZN(n112) );
  AOI21_X1 U556 ( .B1(n573), .B2(n120), .A(n117), .ZN(n115) );
  INV_X1 U557 ( .A(n119), .ZN(n117) );
  INV_X1 U558 ( .A(n122), .ZN(n120) );
  NAND2_X1 U559 ( .A1(n186), .A2(n195), .ZN(n83) );
  NOR2_X1 U560 ( .A1(n211), .A2(n204), .ZN(n89) );
  NAND2_X1 U561 ( .A1(n164), .A2(n175), .ZN(n76) );
  NAND2_X1 U562 ( .A1(n196), .A2(n203), .ZN(n86) );
  NAND2_X1 U563 ( .A1(n204), .A2(n211), .ZN(n90) );
  NAND2_X1 U564 ( .A1(n212), .A2(n217), .ZN(n95) );
  XNOR2_X1 U565 ( .A(n59), .B(n120), .ZN(product[2]) );
  NAND2_X1 U566 ( .A1(n573), .A2(n119), .ZN(n59) );
  XNOR2_X1 U567 ( .A(n63), .B(n46), .ZN(product[15]) );
  NAND2_X1 U568 ( .A1(n575), .A2(n62), .ZN(n46) );
  NAND2_X1 U569 ( .A1(n73), .A2(n572), .ZN(n64) );
  NAND2_X1 U570 ( .A1(n517), .A2(n106), .ZN(n56) );
  NAND2_X1 U571 ( .A1(n329), .A2(n258), .ZN(n122) );
  NAND2_X1 U572 ( .A1(n328), .A2(n314), .ZN(n119) );
  OR2_X1 U573 ( .A1(n328), .A2(n314), .ZN(n573) );
  NOR2_X1 U574 ( .A1(n218), .A2(n223), .ZN(n97) );
  NAND2_X1 U575 ( .A1(n218), .A2(n223), .ZN(n98) );
  NAND2_X1 U576 ( .A1(n224), .A2(n227), .ZN(n103) );
  NAND2_X1 U577 ( .A1(n228), .A2(n231), .ZN(n106) );
  OR2_X1 U578 ( .A1(n139), .A2(n151), .ZN(n575) );
  NAND2_X1 U579 ( .A1(n232), .A2(n233), .ZN(n111) );
  OR2_X1 U580 ( .A1(n232), .A2(n233), .ZN(n576) );
  OR2_X1 U581 ( .A1(n583), .A2(n556), .ZN(n392) );
  AND2_X1 U582 ( .A1(n584), .A2(n564), .ZN(n278) );
  XNOR2_X1 U583 ( .A(n535), .B(n583), .ZN(n352) );
  XNOR2_X1 U584 ( .A(n155), .B(n577), .ZN(n139) );
  XNOR2_X1 U585 ( .A(n153), .B(n141), .ZN(n577) );
  XNOR2_X1 U586 ( .A(n157), .B(n578), .ZN(n141) );
  XNOR2_X1 U587 ( .A(n145), .B(n143), .ZN(n578) );
  OAI22_X1 U588 ( .A1(n42), .A2(n601), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U589 ( .A1(n583), .A2(n601), .ZN(n332) );
  XNOR2_X1 U590 ( .A(n531), .B(n583), .ZN(n343) );
  XNOR2_X1 U591 ( .A(n159), .B(n579), .ZN(n142) );
  XNOR2_X1 U592 ( .A(n315), .B(n261), .ZN(n579) );
  XNOR2_X1 U593 ( .A(n591), .B(n583), .ZN(n376) );
  AND2_X1 U594 ( .A1(n584), .A2(n245), .ZN(n300) );
  XNOR2_X1 U595 ( .A(n598), .B(n583), .ZN(n336) );
  OAI22_X1 U596 ( .A1(n39), .A2(n336), .B1(n513), .B2(n335), .ZN(n263) );
  AND2_X1 U597 ( .A1(n584), .A2(n237), .ZN(n264) );
  INV_X1 U598 ( .A(n19), .ZN(n593) );
  INV_X1 U599 ( .A(n25), .ZN(n595) );
  AND2_X1 U600 ( .A1(n584), .A2(n491), .ZN(n288) );
  AND2_X1 U601 ( .A1(n584), .A2(n563), .ZN(n270) );
  AND2_X1 U602 ( .A1(n584), .A2(n235), .ZN(n260) );
  OAI22_X1 U603 ( .A1(n39), .A2(n335), .B1(n513), .B2(n334), .ZN(n262) );
  INV_X1 U604 ( .A(n7), .ZN(n589) );
  INV_X1 U605 ( .A(n13), .ZN(n592) );
  INV_X1 U606 ( .A(n41), .ZN(n235) );
  INV_X1 U607 ( .A(n37), .ZN(n237) );
  XNOR2_X1 U608 ( .A(n557), .B(n583), .ZN(n363) );
  OAI22_X1 U609 ( .A1(n39), .A2(n599), .B1(n337), .B2(n513), .ZN(n252) );
  OR2_X1 U610 ( .A1(n583), .A2(n599), .ZN(n337) );
  AND2_X1 U611 ( .A1(n584), .A2(n247), .ZN(n314) );
  AND2_X1 U612 ( .A1(n584), .A2(n249), .ZN(product[0]) );
  OR2_X1 U613 ( .A1(n583), .A2(n526), .ZN(n377) );
  OR2_X1 U614 ( .A1(n583), .A2(n593), .ZN(n364) );
  OR2_X1 U615 ( .A1(n583), .A2(n595), .ZN(n353) );
  OR2_X1 U616 ( .A1(n583), .A2(n597), .ZN(n344) );
  XNOR2_X1 U617 ( .A(n596), .B(a[12]), .ZN(n37) );
  XNOR2_X1 U618 ( .A(n598), .B(a[14]), .ZN(n41) );
  OAI22_X1 U619 ( .A1(n39), .A2(n334), .B1(n513), .B2(n333), .ZN(n261) );
  XNOR2_X1 U620 ( .A(n598), .B(n422), .ZN(n333) );
  XNOR2_X1 U621 ( .A(n557), .B(b[9]), .ZN(n354) );
  XNOR2_X1 U622 ( .A(n591), .B(b[11]), .ZN(n365) );
  OAI22_X1 U623 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U624 ( .A(n600), .B(n424), .ZN(n330) );
  XNOR2_X1 U625 ( .A(n600), .B(n583), .ZN(n331) );
  XNOR2_X1 U626 ( .A(n598), .B(n424), .ZN(n335) );
  XNOR2_X1 U627 ( .A(n535), .B(n418), .ZN(n345) );
  XNOR2_X1 U628 ( .A(n531), .B(n420), .ZN(n338) );
  XNOR2_X1 U629 ( .A(n554), .B(b[13]), .ZN(n378) );
  XNOR2_X1 U630 ( .A(n557), .B(n424), .ZN(n362) );
  XNOR2_X1 U631 ( .A(n594), .B(n424), .ZN(n351) );
  XNOR2_X1 U632 ( .A(n532), .B(n424), .ZN(n342) );
  XNOR2_X1 U633 ( .A(n531), .B(n422), .ZN(n340) );
  XNOR2_X1 U634 ( .A(n532), .B(n421), .ZN(n339) );
  XNOR2_X1 U635 ( .A(n554), .B(n418), .ZN(n384) );
  XNOR2_X1 U636 ( .A(n554), .B(n419), .ZN(n385) );
  XNOR2_X1 U637 ( .A(n554), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U638 ( .A(n554), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U639 ( .A(n554), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U640 ( .A(n554), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U641 ( .A(n554), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U642 ( .A(n591), .B(n418), .ZN(n369) );
  XNOR2_X1 U643 ( .A(n591), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U644 ( .A(n591), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U645 ( .A(n591), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U646 ( .A(n566), .B(b[11]), .ZN(n397) );
  XNOR2_X1 U647 ( .A(n566), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U648 ( .A(n565), .B(b[13]), .ZN(n395) );
  XNOR2_X1 U649 ( .A(n586), .B(b[14]), .ZN(n394) );
  XNOR2_X1 U650 ( .A(n557), .B(n420), .ZN(n358) );
  XNOR2_X1 U651 ( .A(n557), .B(n421), .ZN(n359) );
  XNOR2_X1 U652 ( .A(n594), .B(n421), .ZN(n348) );
  XNOR2_X1 U653 ( .A(n535), .B(n420), .ZN(n347) );
  XNOR2_X1 U654 ( .A(n557), .B(n418), .ZN(n356) );
  XNOR2_X1 U655 ( .A(n557), .B(n419), .ZN(n357) );
  XNOR2_X1 U656 ( .A(n535), .B(n419), .ZN(n346) );
  NAND2_X1 U657 ( .A1(n427), .A2(n37), .ZN(n39) );
  XNOR2_X1 U658 ( .A(n557), .B(b[8]), .ZN(n355) );
  XNOR2_X1 U659 ( .A(n535), .B(n422), .ZN(n349) );
  XNOR2_X1 U660 ( .A(n557), .B(n422), .ZN(n360) );
  NAND2_X1 U661 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U662 ( .A(n600), .B(a[14]), .Z(n426) );
  XNOR2_X1 U663 ( .A(n598), .B(n423), .ZN(n334) );
  XNOR2_X1 U664 ( .A(n586), .B(b[15]), .ZN(n393) );
  BUF_X1 U665 ( .A(n43), .Z(n584) );
  XNOR2_X1 U666 ( .A(n532), .B(n423), .ZN(n341) );
  XNOR2_X1 U667 ( .A(n594), .B(n423), .ZN(n350) );
  XNOR2_X1 U668 ( .A(n557), .B(n423), .ZN(n361) );
  XOR2_X1 U669 ( .A(n598), .B(a[12]), .Z(n427) );
  XNOR2_X1 U670 ( .A(n585), .B(a[2]), .ZN(n9) );
  NOR2_X1 U671 ( .A1(n228), .A2(n231), .ZN(n105) );
  XNOR2_X1 U672 ( .A(n77), .B(n48), .ZN(product[13]) );
  XNOR2_X1 U673 ( .A(n70), .B(n47), .ZN(product[14]) );
  INV_X1 U674 ( .A(n512), .ZN(n127) );
  NOR2_X1 U675 ( .A1(n85), .A2(n82), .ZN(n80) );
  OAI21_X1 U676 ( .B1(n82), .B2(n86), .A(n83), .ZN(n81) );
  OAI22_X1 U677 ( .A1(n34), .A2(n339), .B1(n338), .B2(n32), .ZN(n265) );
  OAI22_X1 U678 ( .A1(n34), .A2(n340), .B1(n339), .B2(n32), .ZN(n266) );
  OAI22_X1 U679 ( .A1(n34), .A2(n341), .B1(n340), .B2(n32), .ZN(n267) );
  OAI22_X1 U680 ( .A1(n34), .A2(n342), .B1(n341), .B2(n32), .ZN(n268) );
  OAI22_X1 U681 ( .A1(n34), .A2(n343), .B1(n342), .B2(n32), .ZN(n269) );
  OAI22_X1 U682 ( .A1(n34), .A2(n597), .B1(n344), .B2(n32), .ZN(n253) );
  OAI22_X1 U683 ( .A1(n29), .A2(n346), .B1(n345), .B2(n544), .ZN(n271) );
  OAI22_X1 U684 ( .A1(n29), .A2(n350), .B1(n349), .B2(n544), .ZN(n275) );
  OAI22_X1 U685 ( .A1(n29), .A2(n347), .B1(n346), .B2(n544), .ZN(n272) );
  OAI22_X1 U686 ( .A1(n29), .A2(n348), .B1(n347), .B2(n544), .ZN(n273) );
  OAI22_X1 U687 ( .A1(n29), .A2(n349), .B1(n348), .B2(n530), .ZN(n274) );
  OAI22_X1 U688 ( .A1(n29), .A2(n595), .B1(n353), .B2(n530), .ZN(n254) );
  OAI22_X1 U689 ( .A1(n29), .A2(n351), .B1(n350), .B2(n530), .ZN(n276) );
  OAI22_X1 U690 ( .A1(n29), .A2(n352), .B1(n351), .B2(n544), .ZN(n277) );
  XOR2_X1 U691 ( .A(n546), .B(n54), .Z(product[7]) );
  XNOR2_X1 U692 ( .A(n55), .B(n510), .ZN(product[6]) );
  NAND2_X1 U693 ( .A1(n576), .A2(n111), .ZN(n57) );
  INV_X1 U694 ( .A(n518), .ZN(n586) );
  OR2_X1 U695 ( .A1(n583), .A2(n528), .ZN(n409) );
  INV_X1 U696 ( .A(n1), .ZN(n587) );
  AOI21_X1 U697 ( .B1(n104), .B2(n574), .A(n101), .ZN(n99) );
  OAI21_X1 U698 ( .B1(n105), .B2(n107), .A(n106), .ZN(n104) );
  INV_X1 U699 ( .A(n103), .ZN(n101) );
  NAND2_X1 U700 ( .A1(n151), .A2(n139), .ZN(n62) );
  XNOR2_X1 U701 ( .A(n591), .B(n424), .ZN(n375) );
  XNOR2_X1 U702 ( .A(n591), .B(n423), .ZN(n374) );
  XNOR2_X1 U703 ( .A(n591), .B(n421), .ZN(n372) );
  XNOR2_X1 U704 ( .A(n591), .B(n422), .ZN(n373) );
  XNOR2_X1 U705 ( .A(n591), .B(n419), .ZN(n370) );
  XNOR2_X1 U706 ( .A(n591), .B(n420), .ZN(n371) );
  NOR2_X1 U707 ( .A1(n234), .A2(n257), .ZN(n113) );
  XOR2_X1 U708 ( .A(n58), .B(n115), .Z(product[3]) );
  NAND2_X1 U709 ( .A1(n135), .A2(n114), .ZN(n58) );
  XNOR2_X1 U710 ( .A(n96), .B(n53), .ZN(product[8]) );
  OAI21_X1 U711 ( .B1(n99), .B2(n97), .A(n98), .ZN(n96) );
  XNOR2_X1 U712 ( .A(n57), .B(n112), .ZN(product[4]) );
  OAI22_X1 U713 ( .A1(n559), .A2(n395), .B1(n394), .B2(n582), .ZN(n316) );
  OAI22_X1 U714 ( .A1(n559), .A2(n394), .B1(n393), .B2(n582), .ZN(n315) );
  OAI22_X1 U715 ( .A1(n558), .A2(n396), .B1(n395), .B2(n582), .ZN(n317) );
  OAI22_X1 U716 ( .A1(n559), .A2(n397), .B1(n396), .B2(n582), .ZN(n318) );
  OAI22_X1 U717 ( .A1(n558), .A2(n402), .B1(n401), .B2(n582), .ZN(n323) );
  OAI22_X1 U718 ( .A1(n558), .A2(n401), .B1(n400), .B2(n582), .ZN(n322) );
  OAI22_X1 U719 ( .A1(n559), .A2(n398), .B1(n397), .B2(n582), .ZN(n319) );
  OAI22_X1 U720 ( .A1(n558), .A2(n400), .B1(n399), .B2(n582), .ZN(n321) );
  OAI22_X1 U721 ( .A1(n558), .A2(n399), .B1(n398), .B2(n582), .ZN(n320) );
  OAI22_X1 U722 ( .A1(n6), .A2(n404), .B1(n403), .B2(n582), .ZN(n325) );
  OAI22_X1 U723 ( .A1(n6), .A2(n405), .B1(n404), .B2(n582), .ZN(n326) );
  OAI22_X1 U724 ( .A1(n559), .A2(n403), .B1(n402), .B2(n582), .ZN(n324) );
  OAI22_X1 U725 ( .A1(n6), .A2(n406), .B1(n405), .B2(n582), .ZN(n327) );
  OAI22_X1 U726 ( .A1(n559), .A2(n407), .B1(n406), .B2(n582), .ZN(n328) );
  OAI22_X1 U727 ( .A1(n6), .A2(n408), .B1(n407), .B2(n582), .ZN(n329) );
  OAI22_X1 U728 ( .A1(n6), .A2(n518), .B1(n409), .B2(n582), .ZN(n258) );
  OAI22_X1 U729 ( .A1(n499), .A2(n362), .B1(n361), .B2(n514), .ZN(n286) );
  OAI22_X1 U730 ( .A1(n553), .A2(n358), .B1(n357), .B2(n515), .ZN(n282) );
  OAI22_X1 U731 ( .A1(n553), .A2(n356), .B1(n355), .B2(n527), .ZN(n280) );
  OAI22_X1 U732 ( .A1(n23), .A2(n593), .B1(n364), .B2(n568), .ZN(n255) );
  OAI22_X1 U733 ( .A1(n553), .A2(n363), .B1(n362), .B2(n568), .ZN(n287) );
  OAI22_X1 U734 ( .A1(n499), .A2(n357), .B1(n356), .B2(n527), .ZN(n281) );
  OAI22_X1 U735 ( .A1(n553), .A2(n361), .B1(n360), .B2(n568), .ZN(n285) );
  OAI22_X1 U736 ( .A1(n553), .A2(n360), .B1(n359), .B2(n568), .ZN(n284) );
  OAI22_X1 U737 ( .A1(n553), .A2(n355), .B1(n354), .B2(n568), .ZN(n279) );
  OAI22_X1 U738 ( .A1(n23), .A2(n359), .B1(n358), .B2(n568), .ZN(n283) );
  OAI21_X1 U739 ( .B1(n87), .B2(n494), .A(n86), .ZN(n84) );
  OAI22_X1 U740 ( .A1(n534), .A2(n370), .B1(n369), .B2(n580), .ZN(n293) );
  OAI22_X1 U741 ( .A1(n534), .A2(n367), .B1(n366), .B2(n580), .ZN(n290) );
  OAI22_X1 U742 ( .A1(n534), .A2(n375), .B1(n374), .B2(n580), .ZN(n298) );
  OAI22_X1 U743 ( .A1(n18), .A2(n372), .B1(n371), .B2(n580), .ZN(n295) );
  OAI22_X1 U744 ( .A1(n534), .A2(n368), .B1(n367), .B2(n580), .ZN(n291) );
  OAI22_X1 U745 ( .A1(n18), .A2(n369), .B1(n368), .B2(n580), .ZN(n292) );
  OAI22_X1 U746 ( .A1(n18), .A2(n371), .B1(n370), .B2(n580), .ZN(n294) );
  OAI22_X1 U747 ( .A1(n534), .A2(n526), .B1(n377), .B2(n580), .ZN(n256) );
  OAI22_X1 U748 ( .A1(n534), .A2(n373), .B1(n372), .B2(n580), .ZN(n296) );
  OAI22_X1 U749 ( .A1(n534), .A2(n376), .B1(n375), .B2(n580), .ZN(n299) );
  OAI22_X1 U750 ( .A1(n18), .A2(n374), .B1(n373), .B2(n580), .ZN(n297) );
  OAI22_X1 U751 ( .A1(n534), .A2(n366), .B1(n365), .B2(n580), .ZN(n289) );
  XNOR2_X1 U752 ( .A(n554), .B(n420), .ZN(n386) );
  INV_X1 U753 ( .A(n580), .ZN(n245) );
  XNOR2_X1 U754 ( .A(n588), .B(n422), .ZN(n388) );
  XNOR2_X1 U755 ( .A(n554), .B(n583), .ZN(n391) );
  XNOR2_X1 U756 ( .A(n554), .B(n421), .ZN(n387) );
  XNOR2_X1 U757 ( .A(n554), .B(n424), .ZN(n390) );
  XNOR2_X1 U758 ( .A(n588), .B(n423), .ZN(n389) );
  INV_X1 U759 ( .A(n547), .ZN(n87) );
  XNOR2_X1 U760 ( .A(n565), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U761 ( .A(n586), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U762 ( .A(n586), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U763 ( .A(n566), .B(n418), .ZN(n401) );
  XNOR2_X1 U764 ( .A(n566), .B(n421), .ZN(n404) );
  XNOR2_X1 U765 ( .A(n565), .B(n422), .ZN(n405) );
  XNOR2_X1 U766 ( .A(n586), .B(n420), .ZN(n403) );
  XNOR2_X1 U767 ( .A(n565), .B(n419), .ZN(n402) );
  AOI21_X1 U768 ( .B1(n576), .B2(n112), .A(n109), .ZN(n107) );
  OAI21_X1 U769 ( .B1(n567), .B2(n78), .A(n505), .ZN(n77) );
  OAI21_X1 U770 ( .B1(n64), .B2(n548), .A(n65), .ZN(n63) );
  AOI21_X1 U771 ( .B1(n80), .B2(n511), .A(n516), .ZN(n45) );
  XNOR2_X1 U772 ( .A(n566), .B(n424), .ZN(n407) );
  XNOR2_X1 U773 ( .A(n565), .B(n583), .ZN(n408) );
  XNOR2_X1 U774 ( .A(n565), .B(n423), .ZN(n406) );
  XOR2_X1 U775 ( .A(n56), .B(n490), .Z(product[5]) );
  OAI21_X1 U776 ( .B1(n567), .B2(n503), .A(n72), .ZN(n70) );
  INV_X1 U777 ( .A(n111), .ZN(n109) );
  OAI22_X1 U778 ( .A1(n538), .A2(n379), .B1(n378), .B2(n496), .ZN(n301) );
  OAI22_X1 U779 ( .A1(n538), .A2(n380), .B1(n379), .B2(n496), .ZN(n302) );
  OAI22_X1 U780 ( .A1(n537), .A2(n385), .B1(n384), .B2(n496), .ZN(n307) );
  OAI22_X1 U781 ( .A1(n537), .A2(n382), .B1(n381), .B2(n496), .ZN(n304) );
  OAI22_X1 U782 ( .A1(n538), .A2(n381), .B1(n380), .B2(n496), .ZN(n303) );
  NAND2_X1 U783 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U784 ( .A1(n536), .A2(n383), .B1(n382), .B2(n581), .ZN(n305) );
  OAI22_X1 U785 ( .A1(n538), .A2(n384), .B1(n383), .B2(n496), .ZN(n306) );
  OAI22_X1 U786 ( .A1(n537), .A2(n386), .B1(n385), .B2(n581), .ZN(n308) );
  OAI22_X1 U787 ( .A1(n538), .A2(n387), .B1(n386), .B2(n496), .ZN(n309) );
  OAI22_X1 U788 ( .A1(n537), .A2(n556), .B1(n392), .B2(n496), .ZN(n257) );
  OAI22_X1 U789 ( .A1(n536), .A2(n389), .B1(n388), .B2(n581), .ZN(n311) );
  OAI22_X1 U790 ( .A1(n537), .A2(n388), .B1(n387), .B2(n496), .ZN(n310) );
  OAI22_X1 U791 ( .A1(n537), .A2(n390), .B1(n389), .B2(n496), .ZN(n312) );
  INV_X1 U792 ( .A(n496), .ZN(n247) );
  OAI22_X1 U793 ( .A1(n538), .A2(n391), .B1(n390), .B2(n496), .ZN(n313) );
  BUF_X4 U794 ( .A(n43), .Z(n583) );
  INV_X1 U795 ( .A(n31), .ZN(n597) );
  INV_X1 U796 ( .A(n599), .ZN(n598) );
  INV_X1 U797 ( .A(n36), .ZN(n599) );
  INV_X1 U798 ( .A(n601), .ZN(n600) );
  INV_X1 U799 ( .A(n40), .ZN(n601) );
  XOR2_X1 U800 ( .A(n259), .B(n251), .Z(n148) );
  XOR2_X1 U801 ( .A(n289), .B(n279), .Z(n146) );
endmodule


module layer1_8_4_8_16_datapath_M8_N4_T16_P8_3_DW01_add_2 ( A, B, CI, SUM, CO
 );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n19, n20, n21, n25, n26, n27, n28, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n48, n49, n51, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n71, n72, n73, n74,
         n75, n77, n79, n80, n81, n82, n83, n85, n87, n88, n90, n94, n95, n98,
         n99, n100, n102, n104, n161, n162, n163, n164, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190;

  OR2_X2 U126 ( .A1(A[10]), .A2(B[10]), .ZN(n189) );
  OR2_X1 U127 ( .A1(A[10]), .A2(B[10]), .ZN(n169) );
  OR2_X1 U128 ( .A1(A[14]), .A2(B[14]), .ZN(n161) );
  OR2_X1 U129 ( .A1(A[14]), .A2(B[14]), .ZN(n188) );
  NAND2_X1 U130 ( .A1(A[11]), .A2(B[11]), .ZN(n162) );
  INV_X1 U131 ( .A(n173), .ZN(n163) );
  OR2_X1 U132 ( .A1(A[9]), .A2(B[9]), .ZN(n164) );
  AND2_X1 U133 ( .A1(n183), .A2(n90), .ZN(SUM[0]) );
  NOR2_X1 U134 ( .A1(A[8]), .A2(B[8]), .ZN(n166) );
  NOR2_X1 U135 ( .A1(A[8]), .A2(B[8]), .ZN(n58) );
  XNOR2_X1 U136 ( .A(n49), .B(n167), .ZN(SUM[10]) );
  AND2_X1 U137 ( .A1(n189), .A2(n48), .ZN(n167) );
  AOI21_X1 U138 ( .B1(n56), .B2(n64), .A(n57), .ZN(n168) );
  AOI21_X1 U139 ( .B1(n56), .B2(n64), .A(n57), .ZN(n55) );
  XNOR2_X1 U140 ( .A(n178), .B(n5), .ZN(SUM[11]) );
  CLKBUF_X1 U141 ( .A(n37), .Z(n170) );
  INV_X1 U142 ( .A(n174), .ZN(n25) );
  OR2_X1 U143 ( .A1(A[13]), .A2(B[13]), .ZN(n171) );
  NOR2_X1 U144 ( .A1(n36), .A2(n39), .ZN(n172) );
  NOR2_X2 U145 ( .A1(A[11]), .A2(B[11]), .ZN(n39) );
  AND2_X1 U146 ( .A1(A[13]), .A2(B[13]), .ZN(n173) );
  OR2_X1 U147 ( .A1(n185), .A2(n17), .ZN(n1) );
  AND2_X1 U148 ( .A1(A[14]), .A2(B[14]), .ZN(n174) );
  AOI21_X1 U149 ( .B1(n189), .B2(n51), .A(n190), .ZN(n175) );
  NOR2_X1 U150 ( .A1(A[12]), .A2(B[12]), .ZN(n176) );
  NOR2_X1 U151 ( .A1(A[12]), .A2(B[12]), .ZN(n177) );
  NOR2_X1 U152 ( .A1(A[12]), .A2(B[12]), .ZN(n36) );
  OAI21_X1 U153 ( .B1(n43), .B2(n55), .A(n175), .ZN(n178) );
  OAI21_X1 U154 ( .B1(n177), .B2(n40), .A(n37), .ZN(n179) );
  OAI21_X1 U155 ( .B1(n177), .B2(n40), .A(n37), .ZN(n180) );
  AOI21_X1 U156 ( .B1(n178), .B2(n34), .A(n179), .ZN(n181) );
  AOI21_X1 U157 ( .B1(n42), .B2(n34), .A(n35), .ZN(n182) );
  NOR2_X1 U158 ( .A1(A[7]), .A2(B[7]), .ZN(n61) );
  OR2_X1 U159 ( .A1(A[0]), .A2(B[0]), .ZN(n183) );
  INV_X1 U160 ( .A(n64), .ZN(n63) );
  INV_X1 U161 ( .A(n168), .ZN(n54) );
  AOI21_X1 U162 ( .B1(n42), .B2(n172), .A(n180), .ZN(n33) );
  AOI21_X1 U163 ( .B1(n184), .B2(n88), .A(n85), .ZN(n83) );
  INV_X1 U164 ( .A(n87), .ZN(n85) );
  AOI21_X1 U165 ( .B1(n187), .B2(n72), .A(n69), .ZN(n67) );
  INV_X1 U166 ( .A(n71), .ZN(n69) );
  AOI21_X1 U167 ( .B1(n186), .B2(n80), .A(n77), .ZN(n75) );
  INV_X1 U168 ( .A(n79), .ZN(n77) );
  OAI21_X1 U169 ( .B1(n83), .B2(n81), .A(n82), .ZN(n80) );
  INV_X1 U170 ( .A(n90), .ZN(n88) );
  OAI21_X1 U171 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  INV_X1 U172 ( .A(n39), .ZN(n95) );
  NAND2_X1 U173 ( .A1(n164), .A2(n53), .ZN(n7) );
  NAND2_X1 U174 ( .A1(n99), .A2(n62), .ZN(n9) );
  INV_X1 U175 ( .A(n61), .ZN(n99) );
  NAND2_X1 U176 ( .A1(n187), .A2(n71), .ZN(n11) );
  NAND2_X1 U177 ( .A1(n104), .A2(n82), .ZN(n14) );
  INV_X1 U178 ( .A(n81), .ZN(n104) );
  NAND2_X1 U179 ( .A1(n98), .A2(n59), .ZN(n8) );
  NAND2_X1 U180 ( .A1(n186), .A2(n79), .ZN(n13) );
  NAND2_X1 U181 ( .A1(n184), .A2(n87), .ZN(n15) );
  NAND2_X1 U182 ( .A1(n100), .A2(n66), .ZN(n10) );
  INV_X1 U183 ( .A(n65), .ZN(n100) );
  NAND2_X1 U184 ( .A1(n102), .A2(n74), .ZN(n12) );
  INV_X1 U185 ( .A(n73), .ZN(n102) );
  NAND2_X1 U186 ( .A1(n94), .A2(n170), .ZN(n4) );
  NAND2_X1 U187 ( .A1(n95), .A2(n162), .ZN(n5) );
  XOR2_X1 U188 ( .A(n63), .B(n9), .Z(SUM[7]) );
  XNOR2_X1 U189 ( .A(n15), .B(n88), .ZN(SUM[1]) );
  NAND2_X1 U190 ( .A1(n171), .A2(n28), .ZN(n3) );
  NOR2_X1 U191 ( .A1(A[2]), .A2(B[2]), .ZN(n81) );
  NAND2_X1 U192 ( .A1(A[11]), .A2(B[11]), .ZN(n40) );
  OR2_X1 U193 ( .A1(A[1]), .A2(B[1]), .ZN(n184) );
  AND2_X1 U194 ( .A1(A[15]), .A2(B[15]), .ZN(n185) );
  XNOR2_X1 U195 ( .A(n60), .B(n8), .ZN(SUM[8]) );
  XNOR2_X1 U196 ( .A(n54), .B(n7), .ZN(SUM[9]) );
  NOR2_X1 U197 ( .A1(A[6]), .A2(B[6]), .ZN(n65) );
  NOR2_X1 U198 ( .A1(A[4]), .A2(B[4]), .ZN(n73) );
  NAND2_X1 U199 ( .A1(A[7]), .A2(B[7]), .ZN(n62) );
  OR2_X1 U200 ( .A1(A[3]), .A2(B[3]), .ZN(n186) );
  NAND2_X1 U201 ( .A1(A[2]), .A2(B[2]), .ZN(n82) );
  OR2_X1 U202 ( .A1(A[5]), .A2(B[5]), .ZN(n187) );
  NAND2_X1 U203 ( .A1(A[3]), .A2(B[3]), .ZN(n79) );
  NAND2_X1 U204 ( .A1(A[1]), .A2(B[1]), .ZN(n87) );
  NAND2_X1 U205 ( .A1(A[0]), .A2(B[0]), .ZN(n90) );
  NAND2_X1 U206 ( .A1(A[6]), .A2(B[6]), .ZN(n66) );
  NAND2_X1 U207 ( .A1(A[4]), .A2(B[4]), .ZN(n74) );
  NAND2_X1 U208 ( .A1(A[8]), .A2(B[8]), .ZN(n59) );
  XNOR2_X1 U209 ( .A(n13), .B(n80), .ZN(SUM[3]) );
  XOR2_X1 U210 ( .A(n14), .B(n83), .Z(SUM[2]) );
  INV_X1 U211 ( .A(n190), .ZN(n48) );
  XOR2_X1 U212 ( .A(n10), .B(n67), .Z(SUM[6]) );
  OAI21_X1 U213 ( .B1(n67), .B2(n65), .A(n66), .ZN(n64) );
  NAND2_X1 U214 ( .A1(A[5]), .A2(B[5]), .ZN(n71) );
  AND2_X1 U215 ( .A1(A[10]), .A2(B[10]), .ZN(n190) );
  XNOR2_X1 U216 ( .A(n19), .B(n1), .ZN(SUM[15]) );
  NAND2_X1 U217 ( .A1(n161), .A2(n25), .ZN(n2) );
  XNOR2_X1 U218 ( .A(n38), .B(n4), .ZN(SUM[12]) );
  OAI21_X1 U219 ( .B1(n41), .B2(n39), .A(n162), .ZN(n38) );
  INV_X1 U220 ( .A(n178), .ZN(n41) );
  NAND2_X1 U221 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  NOR2_X1 U222 ( .A1(A[13]), .A2(B[13]), .ZN(n27) );
  AOI21_X1 U223 ( .B1(n54), .B2(n164), .A(n51), .ZN(n49) );
  NAND2_X1 U224 ( .A1(A[9]), .A2(B[9]), .ZN(n53) );
  INV_X1 U225 ( .A(n53), .ZN(n51) );
  NOR2_X1 U226 ( .A1(n36), .A2(n39), .ZN(n34) );
  OAI21_X1 U227 ( .B1(n176), .B2(n40), .A(n37), .ZN(n35) );
  INV_X1 U228 ( .A(n176), .ZN(n94) );
  AOI21_X1 U229 ( .B1(n188), .B2(n173), .A(n174), .ZN(n21) );
  NAND2_X1 U230 ( .A1(A[12]), .A2(B[12]), .ZN(n37) );
  OAI21_X1 U231 ( .B1(n43), .B2(n55), .A(n44), .ZN(n42) );
  AOI21_X1 U232 ( .B1(n189), .B2(n51), .A(n190), .ZN(n44) );
  XNOR2_X1 U233 ( .A(n11), .B(n72), .ZN(SUM[5]) );
  OAI21_X1 U234 ( .B1(n75), .B2(n73), .A(n74), .ZN(n72) );
  XOR2_X1 U235 ( .A(n12), .B(n75), .Z(SUM[4]) );
  INV_X1 U236 ( .A(n166), .ZN(n98) );
  NOR2_X1 U237 ( .A1(n166), .A2(n61), .ZN(n56) );
  OAI21_X1 U238 ( .B1(n58), .B2(n62), .A(n59), .ZN(n57) );
  NOR2_X1 U239 ( .A1(A[15]), .A2(B[15]), .ZN(n17) );
  NAND2_X1 U240 ( .A1(n169), .A2(n164), .ZN(n43) );
  NAND2_X1 U241 ( .A1(n161), .A2(n171), .ZN(n20) );
  XNOR2_X1 U242 ( .A(n26), .B(n2), .ZN(SUM[14]) );
  XOR2_X1 U243 ( .A(n33), .B(n3), .Z(SUM[13]) );
  OAI21_X1 U244 ( .B1(n182), .B2(n27), .A(n163), .ZN(n26) );
  OAI21_X1 U245 ( .B1(n181), .B2(n20), .A(n21), .ZN(n19) );
endmodule


module layer1_8_4_8_16_datapath_M8_N4_T16_P8_3 ( clk, clear_acc, data_out_x, 
        data_out, data_out_w, data_out_b, wr_en_y, m_valid, m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [3:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N27, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, n1, n2, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n87, n104, n113, n114, n115, n116, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n16), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n221), .CK(clk), .Q(n21) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n222), .CK(clk), .Q(n22) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n223), .CK(clk), .Q(n23) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n224), .CK(clk), .Q(n24) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n225), .CK(clk), .Q(n25) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n226), .CK(clk), .Q(n26) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n227), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n228), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n229), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n230), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n231), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n232), .CK(clk), .Q(n34) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n233), .CK(clk), .Q(n35) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n234), .CK(clk), .Q(n36) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n235), .CK(clk), .Q(n37) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n236), .CK(clk), .Q(n39) );
  DFF_X1 \f_reg[0]  ( .D(n104), .CK(clk), .Q(n61), .QN(n210) );
  DFF_X1 \f_reg[1]  ( .D(n87), .CK(clk), .Q(n59), .QN(n211) );
  DFF_X1 \f_reg[2]  ( .D(n85), .CK(clk), .Q(n57), .QN(n212) );
  DFF_X1 \f_reg[3]  ( .D(n84), .CK(clk), .Q(f[3]), .QN(n65) );
  DFF_X1 \f_reg[4]  ( .D(n83), .CK(clk), .Q(f[4]), .QN(n66) );
  DFF_X1 \f_reg[5]  ( .D(n82), .CK(clk), .Q(f[5]), .QN(n67) );
  DFF_X1 \f_reg[6]  ( .D(n81), .CK(clk), .Q(f[6]), .QN(n68) );
  DFF_X1 \f_reg[7]  ( .D(n80), .CK(clk), .Q(f[7]), .QN(n213) );
  DFF_X1 \f_reg[8]  ( .D(n79), .CK(clk), .Q(f[8]), .QN(n214) );
  DFF_X1 \f_reg[9]  ( .D(n78), .CK(clk), .Q(f[9]), .QN(n215) );
  DFF_X1 \f_reg[10]  ( .D(n77), .CK(clk), .Q(n49), .QN(n216) );
  DFF_X1 \f_reg[11]  ( .D(n76), .CK(clk), .Q(n47), .QN(n217) );
  DFF_X1 \f_reg[12]  ( .D(n2), .CK(clk), .Q(n46), .QN(n218) );
  DFF_X1 \f_reg[13]  ( .D(n75), .CK(clk), .Q(n44), .QN(n219) );
  DFF_X1 \f_reg[14]  ( .D(n1), .CK(clk), .Q(n43), .QN(n220) );
  DFF_X1 \f_reg[15]  ( .D(n4), .CK(clk), .Q(f[15]), .QN(n73) );
  DFF_X1 \data_out_reg[1]  ( .D(n176), .CK(clk), .Q(data_out[1]), .QN(n179) );
  DFF_X1 \data_out_reg[0]  ( .D(n177), .CK(clk), .Q(data_out[0]), .QN(n178) );
  layer1_8_4_8_16_datapath_M8_N4_T16_P8_3_DW_mult_tc_1 mult_183 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer1_8_4_8_16_datapath_M8_N4_T16_P8_3_DW01_add_2 add_184 ( .A({n200, n199, 
        n198, n197, n196, n195, n209, n208, n207, n206, n205, n204, n203, n202, 
        n201, n194}), .B({f[15], n43, n44, n46, n47, n49, f[9:3], n57, n59, 
        n61}), .CI(1'b0), .SUM(adder) );
  DFF_X2 delay_reg ( .D(N27), .CK(clk), .Q(n5), .QN(n237) );
  DFF_X1 \data_out_reg[15]  ( .D(n114), .CK(clk), .Q(data_out[15]), .QN(n193)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n115), .CK(clk), .Q(data_out[14]), .QN(n192)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n116), .CK(clk), .Q(data_out[13]), .QN(n191)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n165), .CK(clk), .Q(data_out[12]), .QN(n190)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n166), .CK(clk), .Q(data_out[11]), .QN(n189)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n167), .CK(clk), .Q(data_out[10]), .QN(n188)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n168), .CK(clk), .Q(data_out[9]), .QN(n187) );
  DFF_X1 \data_out_reg[8]  ( .D(n169), .CK(clk), .Q(data_out[8]), .QN(n186) );
  DFF_X1 \data_out_reg[7]  ( .D(n170), .CK(clk), .Q(data_out[7]), .QN(n185) );
  DFF_X1 \data_out_reg[6]  ( .D(n171), .CK(clk), .Q(data_out[6]), .QN(n184) );
  DFF_X1 \data_out_reg[5]  ( .D(n172), .CK(clk), .Q(data_out[5]), .QN(n183) );
  DFF_X1 \data_out_reg[4]  ( .D(n173), .CK(clk), .Q(data_out[4]), .QN(n182) );
  DFF_X1 \data_out_reg[3]  ( .D(n174), .CK(clk), .Q(data_out[3]), .QN(n181) );
  DFF_X1 \data_out_reg[2]  ( .D(n175), .CK(clk), .Q(data_out[2]), .QN(n180) );
  NAND3_X1 U3 ( .A1(n10), .A2(n9), .A3(n11), .ZN(n1) );
  NAND3_X1 U4 ( .A1(n7), .A2(n6), .A3(n8), .ZN(n2) );
  MUX2_X2 U5 ( .A(n26), .B(N39), .S(n237), .Z(n195) );
  NAND3_X1 U6 ( .A1(n13), .A2(n12), .A3(n14), .ZN(n4) );
  MUX2_X2 U8 ( .A(n23), .B(N42), .S(n237), .Z(n198) );
  MUX2_X2 U9 ( .A(n28), .B(N37), .S(n237), .Z(n208) );
  MUX2_X2 U10 ( .A(N44), .B(n21), .S(n5), .Z(n200) );
  MUX2_X2 U11 ( .A(n24), .B(N41), .S(n237), .Z(n197) );
  NAND2_X1 U12 ( .A1(data_out_b[12]), .A2(n16), .ZN(n6) );
  NAND2_X1 U13 ( .A1(adder[12]), .A2(n15), .ZN(n7) );
  NAND2_X1 U14 ( .A1(n63), .A2(n46), .ZN(n8) );
  NAND2_X1 U15 ( .A1(data_out_b[14]), .A2(n16), .ZN(n9) );
  NAND2_X1 U16 ( .A1(adder[14]), .A2(n15), .ZN(n10) );
  NAND2_X1 U17 ( .A1(n63), .A2(n43), .ZN(n11) );
  NAND2_X1 U18 ( .A1(data_out_b[15]), .A2(n16), .ZN(n12) );
  NAND2_X1 U19 ( .A1(adder[15]), .A2(n15), .ZN(n13) );
  NAND2_X1 U20 ( .A1(n63), .A2(f[15]), .ZN(n14) );
  MUX2_X2 U21 ( .A(n25), .B(N40), .S(n237), .Z(n196) );
  INV_X1 U22 ( .A(n17), .ZN(n16) );
  AND2_X2 U23 ( .A1(n42), .A2(n17), .ZN(n15) );
  INV_X1 U24 ( .A(n42), .ZN(n63) );
  INV_X1 U25 ( .A(clear_acc), .ZN(n17) );
  NAND2_X1 U26 ( .A1(n113), .A2(N27), .ZN(n239) );
  INV_X1 U27 ( .A(wr_en_y), .ZN(n113) );
  OAI22_X1 U28 ( .A1(n181), .A2(n239), .B1(n65), .B2(n238), .ZN(n174) );
  OAI22_X1 U29 ( .A1(n182), .A2(n239), .B1(n66), .B2(n238), .ZN(n173) );
  OAI22_X1 U30 ( .A1(n183), .A2(n239), .B1(n67), .B2(n238), .ZN(n172) );
  OAI22_X1 U31 ( .A1(n184), .A2(n239), .B1(n68), .B2(n238), .ZN(n171) );
  OAI22_X1 U32 ( .A1(n185), .A2(n239), .B1(n213), .B2(n238), .ZN(n170) );
  OAI22_X1 U33 ( .A1(n186), .A2(n239), .B1(n214), .B2(n238), .ZN(n169) );
  OAI22_X1 U34 ( .A1(n187), .A2(n239), .B1(n215), .B2(n238), .ZN(n168) );
  INV_X1 U35 ( .A(n20), .ZN(n38) );
  AND3_X1 U36 ( .A1(sel[1]), .A2(sel[2]), .A3(sel[0]), .ZN(n19) );
  INV_X1 U37 ( .A(m_ready), .ZN(n18) );
  NAND2_X1 U38 ( .A1(m_valid), .A2(n18), .ZN(n40) );
  OAI21_X1 U39 ( .B1(sel[3]), .B2(n19), .A(n40), .ZN(N27) );
  NAND2_X1 U40 ( .A1(clear_acc_delay), .A2(n237), .ZN(n20) );
  MUX2_X1 U41 ( .A(n21), .B(N44), .S(n38), .Z(n221) );
  MUX2_X1 U42 ( .A(n22), .B(N43), .S(n38), .Z(n222) );
  MUX2_X1 U43 ( .A(n22), .B(N43), .S(n237), .Z(n199) );
  MUX2_X1 U44 ( .A(n23), .B(N42), .S(n38), .Z(n223) );
  MUX2_X1 U45 ( .A(n24), .B(N41), .S(n38), .Z(n224) );
  MUX2_X1 U46 ( .A(n25), .B(N40), .S(n38), .Z(n225) );
  MUX2_X1 U47 ( .A(n26), .B(N39), .S(n38), .Z(n226) );
  MUX2_X1 U48 ( .A(n27), .B(N38), .S(n38), .Z(n227) );
  MUX2_X1 U49 ( .A(n27), .B(N38), .S(n237), .Z(n209) );
  MUX2_X1 U50 ( .A(n28), .B(N37), .S(n38), .Z(n228) );
  MUX2_X1 U51 ( .A(n29), .B(N36), .S(n38), .Z(n229) );
  MUX2_X1 U52 ( .A(n29), .B(N36), .S(n237), .Z(n207) );
  MUX2_X1 U53 ( .A(n32), .B(N35), .S(n38), .Z(n230) );
  MUX2_X1 U54 ( .A(n32), .B(N35), .S(n237), .Z(n206) );
  MUX2_X1 U55 ( .A(n33), .B(N34), .S(n38), .Z(n231) );
  MUX2_X1 U56 ( .A(n33), .B(N34), .S(n237), .Z(n205) );
  MUX2_X1 U57 ( .A(n34), .B(N33), .S(n38), .Z(n232) );
  MUX2_X1 U58 ( .A(n34), .B(N33), .S(n237), .Z(n204) );
  MUX2_X1 U59 ( .A(n35), .B(N32), .S(n38), .Z(n233) );
  MUX2_X1 U60 ( .A(n35), .B(N32), .S(n237), .Z(n203) );
  MUX2_X1 U61 ( .A(n36), .B(N31), .S(n38), .Z(n234) );
  MUX2_X1 U62 ( .A(n36), .B(N31), .S(n237), .Z(n202) );
  MUX2_X1 U63 ( .A(n37), .B(N30), .S(n38), .Z(n235) );
  MUX2_X1 U64 ( .A(n37), .B(N30), .S(n237), .Z(n201) );
  MUX2_X1 U65 ( .A(n39), .B(N29), .S(n38), .Z(n236) );
  MUX2_X1 U66 ( .A(n39), .B(N29), .S(n237), .Z(n194) );
  INV_X1 U67 ( .A(n40), .ZN(n41) );
  OAI21_X1 U68 ( .B1(n41), .B2(n5), .A(n17), .ZN(n42) );
  AOI222_X1 U69 ( .A1(data_out_b[13]), .A2(n16), .B1(adder[13]), .B2(n15), 
        .C1(n63), .C2(n44), .ZN(n45) );
  INV_X1 U70 ( .A(n45), .ZN(n75) );
  AOI222_X1 U71 ( .A1(data_out_b[11]), .A2(n16), .B1(adder[11]), .B2(n15), 
        .C1(n63), .C2(n47), .ZN(n48) );
  INV_X1 U72 ( .A(n48), .ZN(n76) );
  AOI222_X1 U73 ( .A1(data_out_b[10]), .A2(n16), .B1(adder[10]), .B2(n15), 
        .C1(n63), .C2(n49), .ZN(n50) );
  INV_X1 U74 ( .A(n50), .ZN(n77) );
  AOI222_X1 U75 ( .A1(data_out_b[8]), .A2(n16), .B1(adder[8]), .B2(n15), .C1(
        n63), .C2(f[8]), .ZN(n51) );
  INV_X1 U76 ( .A(n51), .ZN(n79) );
  AOI222_X1 U77 ( .A1(data_out_b[7]), .A2(n16), .B1(adder[7]), .B2(n15), .C1(
        n63), .C2(f[7]), .ZN(n52) );
  INV_X1 U78 ( .A(n52), .ZN(n80) );
  AOI222_X1 U79 ( .A1(data_out_b[6]), .A2(n16), .B1(adder[6]), .B2(n15), .C1(
        n63), .C2(f[6]), .ZN(n53) );
  INV_X1 U80 ( .A(n53), .ZN(n81) );
  AOI222_X1 U81 ( .A1(data_out_b[5]), .A2(n16), .B1(adder[5]), .B2(n15), .C1(
        n63), .C2(f[5]), .ZN(n54) );
  INV_X1 U82 ( .A(n54), .ZN(n82) );
  AOI222_X1 U83 ( .A1(data_out_b[4]), .A2(n16), .B1(adder[4]), .B2(n15), .C1(
        n63), .C2(f[4]), .ZN(n55) );
  INV_X1 U84 ( .A(n55), .ZN(n83) );
  AOI222_X1 U85 ( .A1(data_out_b[3]), .A2(n16), .B1(adder[3]), .B2(n15), .C1(
        n63), .C2(f[3]), .ZN(n56) );
  INV_X1 U86 ( .A(n56), .ZN(n84) );
  AOI222_X1 U87 ( .A1(data_out_b[2]), .A2(n16), .B1(adder[2]), .B2(n15), .C1(
        n63), .C2(n57), .ZN(n58) );
  INV_X1 U88 ( .A(n58), .ZN(n85) );
  AOI222_X1 U89 ( .A1(data_out_b[1]), .A2(n16), .B1(adder[1]), .B2(n15), .C1(
        n63), .C2(n59), .ZN(n60) );
  INV_X1 U90 ( .A(n60), .ZN(n87) );
  AOI222_X1 U91 ( .A1(data_out_b[0]), .A2(n16), .B1(adder[0]), .B2(n15), .C1(
        n63), .C2(n61), .ZN(n62) );
  INV_X1 U92 ( .A(n62), .ZN(n104) );
  AOI222_X1 U93 ( .A1(data_out_b[9]), .A2(n16), .B1(adder[9]), .B2(n15), .C1(
        n63), .C2(f[9]), .ZN(n64) );
  INV_X1 U94 ( .A(n64), .ZN(n78) );
  NOR4_X1 U95 ( .A1(n47), .A2(n46), .A3(n44), .A4(n43), .ZN(n72) );
  NOR4_X1 U96 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n49), .ZN(n71) );
  NAND4_X1 U97 ( .A1(n68), .A2(n67), .A3(n66), .A4(n65), .ZN(n69) );
  NOR4_X1 U98 ( .A1(n69), .A2(n61), .A3(n59), .A4(n57), .ZN(n70) );
  NAND3_X1 U99 ( .A1(n72), .A2(n71), .A3(n70), .ZN(n74) );
  NAND3_X1 U100 ( .A1(wr_en_y), .A2(n74), .A3(n73), .ZN(n238) );
  OAI22_X1 U101 ( .A1(n178), .A2(n239), .B1(n210), .B2(n238), .ZN(n177) );
  OAI22_X1 U102 ( .A1(n179), .A2(n239), .B1(n211), .B2(n238), .ZN(n176) );
  OAI22_X1 U103 ( .A1(n180), .A2(n239), .B1(n212), .B2(n238), .ZN(n175) );
  OAI22_X1 U104 ( .A1(n188), .A2(n239), .B1(n216), .B2(n238), .ZN(n167) );
  OAI22_X1 U105 ( .A1(n189), .A2(n239), .B1(n217), .B2(n238), .ZN(n166) );
  OAI22_X1 U106 ( .A1(n190), .A2(n239), .B1(n218), .B2(n238), .ZN(n165) );
  OAI22_X1 U107 ( .A1(n191), .A2(n239), .B1(n219), .B2(n238), .ZN(n116) );
  OAI22_X1 U108 ( .A1(n192), .A2(n239), .B1(n220), .B2(n238), .ZN(n115) );
  OAI22_X1 U109 ( .A1(n193), .A2(n239), .B1(n73), .B2(n238), .ZN(n114) );
endmodule


module layer1_8_4_8_16_datapath_M8_N4_T16_P8_2_DW_mult_tc_1 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n9, n12, n13, n16, n18, n19, n21, n23, n25, n27, n29, n31,
         n32, n34, n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n50,
         n53, n54, n55, n56, n57, n58, n59, n62, n63, n64, n65, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n86, n87, n88, n89, n90, n91, n93, n95, n96, n97, n98, n99, n101,
         n103, n104, n105, n106, n107, n111, n112, n113, n114, n115, n117,
         n119, n120, n122, n125, n127, n133, n135, n139, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n237, n245, n247, n249, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n418, n419, n420, n421, n422, n423, n424, n426, n427,
         n429, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U148 ( .A(n265), .B(n144), .Z(n145) );
  XOR2_X1 U150 ( .A(n271), .B(n146), .Z(n147) );
  XOR2_X1 U152 ( .A(n301), .B(n148), .Z(n149) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U161 ( .A(n177), .B(n168), .CI(n166), .CO(n163), .S(n164) );
  FA_X1 U162 ( .A(n170), .B(n172), .CI(n179), .CO(n165), .S(n166) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n263), .CI(n291), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n317), .B(n252), .CO(n173), .S(n174) );
  FA_X1 U167 ( .A(n180), .B(n187), .CI(n178), .CO(n175), .S(n176) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U169 ( .A(n193), .B(n282), .CI(n191), .CO(n179), .S(n180) );
  FA_X1 U170 ( .A(n268), .B(n292), .CI(n274), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U172 ( .A(n197), .B(n190), .CI(n188), .CO(n185), .S(n186) );
  FA_X1 U173 ( .A(n199), .B(n201), .CI(n192), .CO(n187), .S(n188) );
  FA_X1 U174 ( .A(n275), .B(n293), .CI(n194), .CO(n189), .S(n190) );
  FA_X1 U175 ( .A(n305), .B(n283), .CI(n253), .CO(n191), .S(n192) );
  HA_X1 U176 ( .A(n319), .B(n269), .CO(n193), .S(n194) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U180 ( .A(n306), .B(n270), .CI(n320), .CO(n201), .S(n202) );
  FA_X1 U181 ( .A(n208), .B(n213), .CI(n206), .CO(n203), .S(n204) );
  FA_X1 U182 ( .A(n210), .B(n307), .CI(n215), .CO(n205), .S(n206) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n308), .B(n278), .CI(n322), .CO(n215), .S(n216) );
  FA_X1 U188 ( .A(n225), .B(n222), .CI(n220), .CO(n217), .S(n218) );
  FA_X1 U189 ( .A(n309), .B(n255), .CI(n297), .CO(n219), .S(n220) );
  HA_X1 U190 ( .A(n287), .B(n323), .CO(n221), .S(n222) );
  FA_X1 U192 ( .A(n324), .B(n288), .CI(n310), .CO(n225), .S(n226) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  HA_X1 U194 ( .A(n325), .B(n311), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n312), .B(n300), .CI(n326), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  CLKBUF_X1 U414 ( .A(n16), .Z(n531) );
  BUF_X1 U415 ( .A(n105), .Z(n498) );
  XNOR2_X1 U416 ( .A(n214), .B(n490), .ZN(n212) );
  XNOR2_X1 U417 ( .A(n219), .B(n216), .ZN(n490) );
  INV_X1 U418 ( .A(n595), .ZN(n491) );
  XOR2_X1 U419 ( .A(n536), .B(n492), .Z(product[9]) );
  NAND2_X1 U420 ( .A1(n511), .A2(n90), .ZN(n492) );
  BUF_X1 U421 ( .A(n533), .Z(n493) );
  AOI21_X1 U422 ( .B1(n537), .B2(n80), .A(n517), .ZN(n533) );
  OR2_X1 U423 ( .A1(n196), .A2(n203), .ZN(n494) );
  OR2_X1 U424 ( .A1(n329), .A2(n258), .ZN(n495) );
  OR2_X1 U425 ( .A1(n218), .A2(n223), .ZN(n496) );
  INV_X1 U426 ( .A(n585), .ZN(n497) );
  INV_X2 U427 ( .A(n598), .ZN(n597) );
  AOI21_X1 U428 ( .B1(n569), .B2(n104), .A(n101), .ZN(n499) );
  CLKBUF_X1 U429 ( .A(n21), .Z(n500) );
  INV_X1 U430 ( .A(n510), .ZN(n501) );
  BUF_X1 U431 ( .A(n584), .Z(n510) );
  CLKBUF_X1 U432 ( .A(n575), .Z(n502) );
  XNOR2_X1 U433 ( .A(n503), .B(n45), .ZN(product[12]) );
  AND2_X1 U434 ( .A1(n504), .A2(n79), .ZN(n503) );
  OR2_X1 U435 ( .A1(n176), .A2(n185), .ZN(n504) );
  NOR2_X1 U436 ( .A1(n186), .A2(n195), .ZN(n505) );
  NOR2_X1 U437 ( .A1(n186), .A2(n195), .ZN(n82) );
  INV_X1 U438 ( .A(n587), .ZN(n586) );
  INV_X2 U439 ( .A(n587), .ZN(n585) );
  CLKBUF_X1 U440 ( .A(n21), .Z(n506) );
  XNOR2_X1 U441 ( .A(n276), .B(n507), .ZN(n200) );
  XNOR2_X1 U442 ( .A(n294), .B(n284), .ZN(n507) );
  CLKBUF_X1 U443 ( .A(n575), .Z(n508) );
  NOR2_X1 U444 ( .A1(n176), .A2(n185), .ZN(n78) );
  XNOR2_X1 U445 ( .A(n587), .B(a[2]), .ZN(n563) );
  INV_X1 U446 ( .A(n591), .ZN(n509) );
  OR2_X1 U447 ( .A1(n204), .A2(n211), .ZN(n511) );
  BUF_X2 U448 ( .A(n9), .Z(n575) );
  INV_X1 U449 ( .A(n19), .ZN(n592) );
  XNOR2_X1 U450 ( .A(n226), .B(n512), .ZN(n224) );
  XNOR2_X1 U451 ( .A(n229), .B(n298), .ZN(n512) );
  XOR2_X1 U452 ( .A(n205), .B(n200), .Z(n513) );
  XOR2_X1 U453 ( .A(n198), .B(n513), .Z(n196) );
  NAND2_X1 U454 ( .A1(n198), .A2(n205), .ZN(n514) );
  NAND2_X1 U455 ( .A1(n198), .A2(n200), .ZN(n515) );
  NAND2_X1 U456 ( .A1(n205), .A2(n200), .ZN(n516) );
  NAND3_X1 U457 ( .A1(n514), .A2(n515), .A3(n516), .ZN(n195) );
  OAI21_X1 U458 ( .B1(n505), .B2(n86), .A(n83), .ZN(n517) );
  XNOR2_X1 U459 ( .A(n88), .B(n518), .ZN(product[10]) );
  NAND2_X1 U460 ( .A1(n494), .A2(n86), .ZN(n518) );
  CLKBUF_X1 U461 ( .A(n104), .Z(n519) );
  NAND2_X1 U462 ( .A1(n429), .A2(n27), .ZN(n520) );
  NAND2_X1 U463 ( .A1(n429), .A2(n27), .ZN(n29) );
  NOR2_X1 U464 ( .A1(n164), .A2(n175), .ZN(n521) );
  NOR2_X1 U465 ( .A1(n164), .A2(n175), .ZN(n75) );
  XNOR2_X1 U466 ( .A(n501), .B(n249), .ZN(n522) );
  NOR2_X1 U467 ( .A1(n196), .A2(n203), .ZN(n523) );
  OAI21_X1 U468 ( .B1(n499), .B2(n97), .A(n98), .ZN(n524) );
  INV_X1 U469 ( .A(n589), .ZN(n525) );
  INV_X1 U470 ( .A(n596), .ZN(n526) );
  INV_X1 U471 ( .A(n596), .ZN(n527) );
  INV_X1 U472 ( .A(n596), .ZN(n595) );
  XNOR2_X1 U473 ( .A(n582), .B(a[2]), .ZN(n9) );
  INV_X1 U474 ( .A(n594), .ZN(n528) );
  NAND2_X1 U475 ( .A1(n9), .A2(n563), .ZN(n529) );
  NAND2_X1 U476 ( .A1(n9), .A2(n563), .ZN(n12) );
  OAI21_X1 U477 ( .B1(n113), .B2(n115), .A(n114), .ZN(n530) );
  INV_X1 U478 ( .A(n553), .ZN(n532) );
  INV_X1 U479 ( .A(n553), .ZN(n27) );
  AOI21_X1 U480 ( .B1(n537), .B2(n80), .A(n81), .ZN(n45) );
  BUF_X2 U481 ( .A(n576), .Z(n534) );
  INV_X1 U482 ( .A(n594), .ZN(n535) );
  INV_X1 U483 ( .A(n594), .ZN(n593) );
  NAND2_X2 U484 ( .A1(n564), .A2(n531), .ZN(n18) );
  AOI21_X1 U485 ( .B1(n96), .B2(n566), .A(n93), .ZN(n536) );
  OAI21_X1 U486 ( .B1(n536), .B2(n89), .A(n90), .ZN(n537) );
  NAND2_X1 U487 ( .A1(n276), .A2(n294), .ZN(n538) );
  NAND2_X1 U488 ( .A1(n276), .A2(n284), .ZN(n539) );
  NAND2_X1 U489 ( .A1(n294), .A2(n284), .ZN(n540) );
  NAND3_X1 U490 ( .A1(n538), .A2(n539), .A3(n540), .ZN(n199) );
  OR2_X2 U491 ( .A1(n557), .A2(n541), .ZN(n34) );
  XNOR2_X1 U492 ( .A(n595), .B(a[10]), .ZN(n541) );
  INV_X1 U493 ( .A(n557), .ZN(n32) );
  XOR2_X1 U494 ( .A(n592), .B(a[6]), .Z(n551) );
  XOR2_X1 U495 ( .A(n254), .B(n295), .Z(n542) );
  XOR2_X1 U496 ( .A(n542), .B(n285), .Z(n208) );
  NAND2_X1 U497 ( .A1(n285), .A2(n254), .ZN(n543) );
  NAND2_X1 U498 ( .A1(n285), .A2(n295), .ZN(n544) );
  NAND2_X1 U499 ( .A1(n254), .A2(n295), .ZN(n545) );
  NAND3_X1 U500 ( .A1(n543), .A2(n544), .A3(n545), .ZN(n207) );
  INV_X1 U501 ( .A(n247), .ZN(n546) );
  XOR2_X1 U502 ( .A(n587), .B(a[4]), .Z(n16) );
  NAND2_X1 U503 ( .A1(n226), .A2(n229), .ZN(n547) );
  NAND2_X1 U504 ( .A1(n226), .A2(n298), .ZN(n548) );
  NAND2_X1 U505 ( .A1(n229), .A2(n298), .ZN(n549) );
  NAND3_X1 U506 ( .A1(n547), .A2(n548), .A3(n549), .ZN(n223) );
  CLKBUF_X1 U507 ( .A(n499), .Z(n550) );
  OR2_X2 U508 ( .A1(n556), .A2(n551), .ZN(n23) );
  INV_X1 U509 ( .A(n556), .ZN(n21) );
  INV_X1 U510 ( .A(n574), .ZN(n552) );
  CLKBUF_X3 U511 ( .A(n582), .Z(n574) );
  XNOR2_X1 U512 ( .A(n592), .B(a[8]), .ZN(n553) );
  OR2_X1 U513 ( .A1(n522), .A2(n558), .ZN(n6) );
  OR2_X2 U514 ( .A1(n522), .A2(n558), .ZN(n554) );
  OR2_X2 U515 ( .A1(n522), .A2(n558), .ZN(n555) );
  XNOR2_X1 U516 ( .A(n590), .B(a[6]), .ZN(n556) );
  XNOR2_X1 U517 ( .A(n594), .B(a[10]), .ZN(n557) );
  INV_X1 U518 ( .A(n249), .ZN(n576) );
  OAI21_X1 U519 ( .B1(n89), .B2(n91), .A(n90), .ZN(n88) );
  INV_X1 U520 ( .A(n576), .ZN(n558) );
  INV_X1 U521 ( .A(n590), .ZN(n588) );
  INV_X2 U522 ( .A(n590), .ZN(n589) );
  CLKBUF_X1 U523 ( .A(n12), .Z(n559) );
  NAND2_X1 U524 ( .A1(n214), .A2(n219), .ZN(n560) );
  NAND2_X1 U525 ( .A1(n214), .A2(n216), .ZN(n561) );
  NAND2_X1 U526 ( .A1(n219), .A2(n216), .ZN(n562) );
  NAND3_X1 U527 ( .A1(n560), .A2(n561), .A3(n562), .ZN(n211) );
  CLKBUF_X3 U528 ( .A(n16), .Z(n573) );
  INV_X2 U529 ( .A(n592), .ZN(n591) );
  XOR2_X1 U530 ( .A(n588), .B(a[4]), .Z(n564) );
  BUF_X1 U531 ( .A(n43), .Z(n580) );
  NAND2_X1 U532 ( .A1(n73), .A2(n565), .ZN(n64) );
  INV_X1 U533 ( .A(n69), .ZN(n67) );
  NAND2_X1 U534 ( .A1(n565), .A2(n69), .ZN(n47) );
  INV_X1 U535 ( .A(n74), .ZN(n72) );
  OAI21_X1 U536 ( .B1(n521), .B2(n79), .A(n76), .ZN(n74) );
  OR2_X1 U537 ( .A1(n152), .A2(n163), .ZN(n565) );
  AOI21_X1 U538 ( .B1(n524), .B2(n566), .A(n93), .ZN(n91) );
  INV_X1 U539 ( .A(n95), .ZN(n93) );
  NAND2_X1 U540 ( .A1(n125), .A2(n76), .ZN(n48) );
  XNOR2_X1 U541 ( .A(n84), .B(n50), .ZN(product[11]) );
  NAND2_X1 U542 ( .A1(n127), .A2(n83), .ZN(n50) );
  XNOR2_X1 U543 ( .A(n96), .B(n53), .ZN(product[8]) );
  NAND2_X1 U544 ( .A1(n566), .A2(n95), .ZN(n53) );
  NAND2_X1 U545 ( .A1(n152), .A2(n163), .ZN(n69) );
  OAI21_X1 U546 ( .B1(n113), .B2(n115), .A(n114), .ZN(n112) );
  OAI21_X1 U547 ( .B1(n99), .B2(n97), .A(n98), .ZN(n96) );
  NAND2_X1 U548 ( .A1(n133), .A2(n106), .ZN(n56) );
  NAND2_X1 U549 ( .A1(n496), .A2(n98), .ZN(n54) );
  AOI21_X1 U550 ( .B1(n567), .B2(n120), .A(n117), .ZN(n115) );
  INV_X1 U551 ( .A(n119), .ZN(n117) );
  NAND2_X1 U552 ( .A1(n568), .A2(n62), .ZN(n46) );
  AOI21_X1 U553 ( .B1(n74), .B2(n565), .A(n67), .ZN(n65) );
  XOR2_X1 U554 ( .A(n58), .B(n115), .Z(product[3]) );
  NAND2_X1 U555 ( .A1(n135), .A2(n114), .ZN(n58) );
  INV_X1 U556 ( .A(n113), .ZN(n135) );
  INV_X1 U557 ( .A(n122), .ZN(n120) );
  XNOR2_X1 U558 ( .A(n57), .B(n530), .ZN(product[4]) );
  NAND2_X1 U559 ( .A1(n577), .A2(n111), .ZN(n57) );
  INV_X1 U560 ( .A(n578), .ZN(n111) );
  NAND2_X1 U561 ( .A1(n176), .A2(n185), .ZN(n79) );
  OR2_X1 U562 ( .A1(n212), .A2(n217), .ZN(n566) );
  NAND2_X1 U563 ( .A1(n212), .A2(n217), .ZN(n95) );
  NAND2_X1 U564 ( .A1(n196), .A2(n203), .ZN(n86) );
  NAND2_X1 U565 ( .A1(n186), .A2(n195), .ZN(n83) );
  XNOR2_X1 U566 ( .A(n59), .B(n120), .ZN(product[2]) );
  NAND2_X1 U567 ( .A1(n567), .A2(n119), .ZN(n59) );
  NOR2_X1 U568 ( .A1(n218), .A2(n223), .ZN(n97) );
  OR2_X1 U569 ( .A1(n328), .A2(n314), .ZN(n567) );
  OR2_X1 U570 ( .A1(n151), .A2(n139), .ZN(n568) );
  OR2_X1 U571 ( .A1(n232), .A2(n233), .ZN(n577) );
  NAND2_X1 U572 ( .A1(n218), .A2(n223), .ZN(n98) );
  OR2_X1 U573 ( .A1(n224), .A2(n227), .ZN(n569) );
  AND2_X1 U574 ( .A1(n495), .A2(n122), .ZN(product[1]) );
  OR2_X1 U575 ( .A1(n580), .A2(n497), .ZN(n392) );
  OAI22_X1 U576 ( .A1(n6), .A2(n404), .B1(n403), .B2(n534), .ZN(n325) );
  OAI22_X1 U577 ( .A1(n554), .A2(n396), .B1(n395), .B2(n534), .ZN(n317) );
  OAI22_X1 U578 ( .A1(n39), .A2(n598), .B1(n337), .B2(n37), .ZN(n252) );
  OR2_X1 U579 ( .A1(n580), .A2(n598), .ZN(n337) );
  OAI22_X1 U580 ( .A1(n555), .A2(n400), .B1(n399), .B2(n534), .ZN(n321) );
  XNOR2_X1 U581 ( .A(n593), .B(n580), .ZN(n352) );
  OAI22_X1 U582 ( .A1(n555), .A2(n406), .B1(n405), .B2(n534), .ZN(n327) );
  XNOR2_X1 U583 ( .A(n585), .B(n580), .ZN(n391) );
  XNOR2_X1 U584 ( .A(n155), .B(n571), .ZN(n139) );
  XNOR2_X1 U585 ( .A(n153), .B(n141), .ZN(n571) );
  XNOR2_X1 U586 ( .A(n157), .B(n572), .ZN(n141) );
  XNOR2_X1 U587 ( .A(n145), .B(n143), .ZN(n572) );
  OAI22_X1 U588 ( .A1(n554), .A2(n408), .B1(n407), .B2(n534), .ZN(n329) );
  OAI22_X1 U589 ( .A1(n42), .A2(n600), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U590 ( .A1(n580), .A2(n600), .ZN(n332) );
  OAI22_X1 U591 ( .A1(n554), .A2(n398), .B1(n397), .B2(n534), .ZN(n319) );
  XNOR2_X1 U592 ( .A(n527), .B(n580), .ZN(n343) );
  XOR2_X1 U593 ( .A(n315), .B(n261), .Z(n150) );
  OAI22_X1 U594 ( .A1(n555), .A2(n394), .B1(n393), .B2(n534), .ZN(n315) );
  XNOR2_X1 U595 ( .A(n597), .B(n580), .ZN(n336) );
  AND2_X1 U596 ( .A1(n581), .A2(n553), .ZN(n278) );
  OAI22_X1 U597 ( .A1(n554), .A2(n401), .B1(n400), .B2(n534), .ZN(n322) );
  OAI22_X1 U598 ( .A1(n39), .A2(n336), .B1(n37), .B2(n335), .ZN(n263) );
  XNOR2_X1 U599 ( .A(n589), .B(n580), .ZN(n376) );
  INV_X1 U600 ( .A(n25), .ZN(n594) );
  AND2_X1 U601 ( .A1(n581), .A2(n237), .ZN(n264) );
  OAI22_X1 U602 ( .A1(n554), .A2(n397), .B1(n396), .B2(n534), .ZN(n318) );
  OAI22_X1 U603 ( .A1(n555), .A2(n405), .B1(n404), .B2(n534), .ZN(n326) );
  AND2_X1 U604 ( .A1(n581), .A2(n245), .ZN(n300) );
  AND2_X1 U605 ( .A1(n581), .A2(n556), .ZN(n288) );
  OAI22_X1 U606 ( .A1(n6), .A2(n403), .B1(n402), .B2(n534), .ZN(n324) );
  AND2_X1 U607 ( .A1(n581), .A2(n557), .ZN(n270) );
  OAI22_X1 U608 ( .A1(n555), .A2(n399), .B1(n398), .B2(n534), .ZN(n320) );
  OAI22_X1 U609 ( .A1(n554), .A2(n395), .B1(n394), .B2(n534), .ZN(n316) );
  AND2_X1 U610 ( .A1(n581), .A2(n235), .ZN(n260) );
  OAI22_X1 U611 ( .A1(n39), .A2(n335), .B1(n37), .B2(n334), .ZN(n262) );
  INV_X1 U612 ( .A(n7), .ZN(n587) );
  INV_X1 U613 ( .A(n41), .ZN(n235) );
  INV_X1 U614 ( .A(n37), .ZN(n237) );
  OAI22_X1 U615 ( .A1(n555), .A2(n402), .B1(n401), .B2(n534), .ZN(n323) );
  XNOR2_X1 U616 ( .A(n591), .B(n580), .ZN(n363) );
  AND2_X1 U617 ( .A1(n581), .A2(n247), .ZN(n314) );
  AND2_X1 U618 ( .A1(n581), .A2(n249), .ZN(product[0]) );
  OR2_X1 U619 ( .A1(n580), .A2(n509), .ZN(n364) );
  OR2_X1 U620 ( .A1(n580), .A2(n491), .ZN(n344) );
  OR2_X1 U621 ( .A1(n580), .A2(n594), .ZN(n353) );
  OR2_X1 U622 ( .A1(n580), .A2(n525), .ZN(n377) );
  XNOR2_X1 U623 ( .A(n595), .B(a[12]), .ZN(n37) );
  XNOR2_X1 U624 ( .A(n597), .B(a[14]), .ZN(n41) );
  OAI22_X1 U625 ( .A1(n39), .A2(n334), .B1(n37), .B2(n333), .ZN(n261) );
  XNOR2_X1 U626 ( .A(n597), .B(n422), .ZN(n333) );
  XNOR2_X1 U627 ( .A(n591), .B(b[9]), .ZN(n354) );
  XNOR2_X1 U628 ( .A(n589), .B(b[11]), .ZN(n365) );
  OAI22_X1 U629 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U630 ( .A(n599), .B(n424), .ZN(n330) );
  XNOR2_X1 U631 ( .A(n599), .B(n580), .ZN(n331) );
  XNOR2_X1 U632 ( .A(n597), .B(n424), .ZN(n335) );
  XNOR2_X1 U633 ( .A(n597), .B(n423), .ZN(n334) );
  XNOR2_X1 U634 ( .A(n583), .B(b[11]), .ZN(n397) );
  XNOR2_X1 U635 ( .A(n583), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U636 ( .A(n583), .B(b[13]), .ZN(n395) );
  XNOR2_X1 U637 ( .A(n583), .B(b[14]), .ZN(n394) );
  XOR2_X1 U638 ( .A(n593), .B(a[8]), .Z(n429) );
  XNOR2_X1 U639 ( .A(n535), .B(n418), .ZN(n345) );
  XNOR2_X1 U640 ( .A(n526), .B(n420), .ZN(n338) );
  XNOR2_X1 U641 ( .A(n585), .B(b[13]), .ZN(n378) );
  XNOR2_X1 U642 ( .A(n591), .B(n424), .ZN(n362) );
  XNOR2_X1 U643 ( .A(n527), .B(n424), .ZN(n342) );
  XNOR2_X1 U644 ( .A(n593), .B(n424), .ZN(n351) );
  XNOR2_X1 U645 ( .A(n526), .B(n423), .ZN(n341) );
  XNOR2_X1 U646 ( .A(n526), .B(n422), .ZN(n340) );
  XNOR2_X1 U647 ( .A(n527), .B(n421), .ZN(n339) );
  XNOR2_X1 U648 ( .A(n586), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U649 ( .A(n585), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U650 ( .A(n586), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U651 ( .A(n585), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U652 ( .A(n585), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U653 ( .A(n585), .B(n418), .ZN(n384) );
  XNOR2_X1 U654 ( .A(n586), .B(n419), .ZN(n385) );
  XNOR2_X1 U655 ( .A(n589), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U656 ( .A(n589), .B(n418), .ZN(n369) );
  XNOR2_X1 U657 ( .A(n589), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U658 ( .A(n589), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U659 ( .A(n535), .B(n422), .ZN(n349) );
  XNOR2_X1 U660 ( .A(n591), .B(n423), .ZN(n361) );
  XNOR2_X1 U661 ( .A(n591), .B(n422), .ZN(n360) );
  XNOR2_X1 U662 ( .A(n528), .B(n423), .ZN(n350) );
  XNOR2_X1 U663 ( .A(n591), .B(n420), .ZN(n358) );
  XNOR2_X1 U664 ( .A(n586), .B(n420), .ZN(n386) );
  XNOR2_X1 U665 ( .A(n528), .B(n420), .ZN(n347) );
  XNOR2_X1 U666 ( .A(n591), .B(n421), .ZN(n359) );
  XNOR2_X1 U667 ( .A(n535), .B(n421), .ZN(n348) );
  XNOR2_X1 U668 ( .A(n591), .B(n418), .ZN(n356) );
  XNOR2_X1 U669 ( .A(n535), .B(n419), .ZN(n346) );
  XNOR2_X1 U670 ( .A(n591), .B(n419), .ZN(n357) );
  NAND2_X1 U671 ( .A1(n427), .A2(n37), .ZN(n39) );
  XNOR2_X1 U672 ( .A(n591), .B(b[8]), .ZN(n355) );
  XNOR2_X1 U673 ( .A(n583), .B(b[15]), .ZN(n393) );
  NAND2_X1 U674 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U675 ( .A(n599), .B(a[14]), .Z(n426) );
  BUF_X1 U676 ( .A(n43), .Z(n581) );
  INV_X1 U677 ( .A(n584), .ZN(n582) );
  XOR2_X1 U678 ( .A(n597), .B(a[12]), .Z(n427) );
  INV_X1 U679 ( .A(n75), .ZN(n125) );
  NOR2_X1 U680 ( .A1(n75), .A2(n78), .ZN(n73) );
  NAND2_X1 U681 ( .A1(n164), .A2(n175), .ZN(n76) );
  INV_X1 U682 ( .A(n498), .ZN(n133) );
  AND2_X1 U683 ( .A1(n232), .A2(n233), .ZN(n578) );
  NAND2_X1 U684 ( .A1(n228), .A2(n231), .ZN(n106) );
  XNOR2_X1 U685 ( .A(n586), .B(n422), .ZN(n388) );
  XNOR2_X1 U686 ( .A(n586), .B(n423), .ZN(n389) );
  XNOR2_X1 U687 ( .A(n585), .B(n424), .ZN(n390) );
  XNOR2_X1 U688 ( .A(n585), .B(n421), .ZN(n387) );
  NOR2_X1 U689 ( .A1(n234), .A2(n257), .ZN(n113) );
  NAND2_X1 U690 ( .A1(n569), .A2(n103), .ZN(n55) );
  INV_X1 U691 ( .A(n103), .ZN(n101) );
  AOI21_X1 U692 ( .B1(n577), .B2(n530), .A(n578), .ZN(n579) );
  NAND2_X1 U693 ( .A1(n204), .A2(n211), .ZN(n90) );
  NOR2_X1 U694 ( .A1(n204), .A2(n211), .ZN(n89) );
  OAI22_X1 U695 ( .A1(n520), .A2(n346), .B1(n345), .B2(n532), .ZN(n271) );
  OAI22_X1 U696 ( .A1(n520), .A2(n350), .B1(n349), .B2(n532), .ZN(n275) );
  OAI22_X1 U697 ( .A1(n520), .A2(n347), .B1(n346), .B2(n532), .ZN(n272) );
  OAI22_X1 U698 ( .A1(n520), .A2(n351), .B1(n350), .B2(n532), .ZN(n276) );
  OAI22_X1 U699 ( .A1(n520), .A2(n349), .B1(n348), .B2(n532), .ZN(n274) );
  OAI22_X1 U700 ( .A1(n29), .A2(n594), .B1(n353), .B2(n532), .ZN(n254) );
  OAI22_X1 U701 ( .A1(n520), .A2(n348), .B1(n347), .B2(n532), .ZN(n273) );
  OAI22_X1 U702 ( .A1(n29), .A2(n352), .B1(n351), .B2(n532), .ZN(n277) );
  XNOR2_X1 U703 ( .A(n77), .B(n48), .ZN(product[13]) );
  XNOR2_X1 U704 ( .A(n70), .B(n47), .ZN(product[14]) );
  INV_X1 U705 ( .A(n505), .ZN(n127) );
  NOR2_X1 U706 ( .A1(n82), .A2(n523), .ZN(n80) );
  OAI21_X1 U707 ( .B1(n82), .B2(n86), .A(n83), .ZN(n81) );
  OAI22_X1 U708 ( .A1(n34), .A2(n339), .B1(n338), .B2(n32), .ZN(n265) );
  OAI22_X1 U709 ( .A1(n34), .A2(n340), .B1(n339), .B2(n32), .ZN(n266) );
  OAI22_X1 U710 ( .A1(n34), .A2(n342), .B1(n341), .B2(n32), .ZN(n268) );
  OAI22_X1 U711 ( .A1(n34), .A2(n341), .B1(n340), .B2(n32), .ZN(n267) );
  OAI22_X1 U712 ( .A1(n34), .A2(n343), .B1(n32), .B2(n342), .ZN(n269) );
  OAI22_X1 U713 ( .A1(n34), .A2(n491), .B1(n344), .B2(n32), .ZN(n253) );
  XNOR2_X1 U714 ( .A(n63), .B(n46), .ZN(product[15]) );
  XNOR2_X1 U715 ( .A(n55), .B(n519), .ZN(product[6]) );
  NOR2_X1 U716 ( .A1(n228), .A2(n231), .ZN(n105) );
  NAND2_X1 U717 ( .A1(n328), .A2(n314), .ZN(n119) );
  AOI21_X1 U718 ( .B1(n577), .B2(n112), .A(n578), .ZN(n107) );
  OAI21_X1 U719 ( .B1(n105), .B2(n107), .A(n106), .ZN(n104) );
  OAI22_X1 U720 ( .A1(n555), .A2(n407), .B1(n406), .B2(n534), .ZN(n328) );
  INV_X1 U721 ( .A(n1), .ZN(n584) );
  OAI22_X1 U722 ( .A1(n23), .A2(n358), .B1(n500), .B2(n357), .ZN(n282) );
  OAI22_X1 U723 ( .A1(n23), .A2(n356), .B1(n355), .B2(n506), .ZN(n280) );
  OAI22_X1 U724 ( .A1(n23), .A2(n357), .B1(n356), .B2(n21), .ZN(n281) );
  OAI22_X1 U725 ( .A1(n23), .A2(n360), .B1(n21), .B2(n359), .ZN(n284) );
  OAI22_X1 U726 ( .A1(n23), .A2(n509), .B1(n364), .B2(n21), .ZN(n255) );
  OAI22_X1 U727 ( .A1(n23), .A2(n362), .B1(n500), .B2(n361), .ZN(n286) );
  OAI22_X1 U728 ( .A1(n23), .A2(n361), .B1(n500), .B2(n360), .ZN(n285) );
  OAI22_X1 U729 ( .A1(n23), .A2(n355), .B1(n21), .B2(n354), .ZN(n279) );
  XNOR2_X1 U730 ( .A(n589), .B(n424), .ZN(n375) );
  OAI22_X1 U731 ( .A1(n23), .A2(n363), .B1(n21), .B2(n362), .ZN(n287) );
  XNOR2_X1 U732 ( .A(n589), .B(n423), .ZN(n374) );
  XNOR2_X1 U733 ( .A(n589), .B(n422), .ZN(n373) );
  XNOR2_X1 U734 ( .A(n589), .B(n421), .ZN(n372) );
  XNOR2_X1 U735 ( .A(n589), .B(n419), .ZN(n370) );
  XNOR2_X1 U736 ( .A(n589), .B(n420), .ZN(n371) );
  XOR2_X1 U737 ( .A(n56), .B(n579), .Z(product[5]) );
  OR2_X1 U738 ( .A1(n580), .A2(n552), .ZN(n409) );
  INV_X1 U739 ( .A(n510), .ZN(n583) );
  NAND2_X1 U740 ( .A1(n224), .A2(n227), .ZN(n103) );
  OAI21_X1 U741 ( .B1(n87), .B2(n523), .A(n86), .ZN(n84) );
  INV_X1 U742 ( .A(n13), .ZN(n590) );
  INV_X1 U743 ( .A(n73), .ZN(n71) );
  OAI22_X1 U744 ( .A1(n23), .A2(n359), .B1(n358), .B2(n21), .ZN(n283) );
  NAND2_X1 U745 ( .A1(n329), .A2(n258), .ZN(n122) );
  INV_X1 U746 ( .A(n88), .ZN(n87) );
  OAI22_X1 U747 ( .A1(n554), .A2(n552), .B1(n409), .B2(n534), .ZN(n258) );
  AOI21_X1 U748 ( .B1(n569), .B2(n104), .A(n101), .ZN(n99) );
  NAND2_X1 U749 ( .A1(n151), .A2(n139), .ZN(n62) );
  OAI22_X1 U750 ( .A1(n18), .A2(n370), .B1(n369), .B2(n573), .ZN(n293) );
  OAI22_X1 U751 ( .A1(n18), .A2(n367), .B1(n366), .B2(n573), .ZN(n290) );
  OAI22_X1 U752 ( .A1(n18), .A2(n375), .B1(n374), .B2(n573), .ZN(n298) );
  OAI22_X1 U753 ( .A1(n18), .A2(n373), .B1(n372), .B2(n573), .ZN(n296) );
  OAI22_X1 U754 ( .A1(n18), .A2(n372), .B1(n371), .B2(n573), .ZN(n295) );
  OAI22_X1 U755 ( .A1(n18), .A2(n368), .B1(n367), .B2(n573), .ZN(n291) );
  OAI22_X1 U756 ( .A1(n18), .A2(n374), .B1(n373), .B2(n573), .ZN(n297) );
  OAI22_X1 U757 ( .A1(n18), .A2(n376), .B1(n375), .B2(n573), .ZN(n299) );
  OAI22_X1 U758 ( .A1(n18), .A2(n525), .B1(n377), .B2(n573), .ZN(n256) );
  OAI22_X1 U759 ( .A1(n18), .A2(n371), .B1(n370), .B2(n573), .ZN(n294) );
  OAI22_X1 U760 ( .A1(n18), .A2(n369), .B1(n368), .B2(n573), .ZN(n292) );
  OAI22_X1 U761 ( .A1(n18), .A2(n366), .B1(n365), .B2(n573), .ZN(n289) );
  INV_X1 U762 ( .A(n573), .ZN(n245) );
  XNOR2_X1 U763 ( .A(n574), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U764 ( .A(n574), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U765 ( .A(n574), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U766 ( .A(n574), .B(n418), .ZN(n401) );
  XNOR2_X1 U767 ( .A(n574), .B(n419), .ZN(n402) );
  XNOR2_X1 U768 ( .A(n574), .B(n420), .ZN(n403) );
  XNOR2_X1 U769 ( .A(n574), .B(n422), .ZN(n405) );
  XNOR2_X1 U770 ( .A(n574), .B(n421), .ZN(n404) );
  XNOR2_X1 U771 ( .A(n574), .B(n580), .ZN(n408) );
  XNOR2_X1 U772 ( .A(n574), .B(n423), .ZN(n406) );
  XNOR2_X1 U773 ( .A(n574), .B(n424), .ZN(n407) );
  OAI21_X1 U774 ( .B1(n533), .B2(n78), .A(n79), .ZN(n77) );
  OAI21_X1 U775 ( .B1(n533), .B2(n71), .A(n72), .ZN(n70) );
  OAI21_X1 U776 ( .B1(n64), .B2(n493), .A(n65), .ZN(n63) );
  XOR2_X1 U777 ( .A(n550), .B(n54), .Z(product[7]) );
  OAI22_X1 U778 ( .A1(n559), .A2(n379), .B1(n378), .B2(n546), .ZN(n301) );
  OAI22_X1 U779 ( .A1(n559), .A2(n380), .B1(n379), .B2(n546), .ZN(n302) );
  OAI22_X1 U780 ( .A1(n559), .A2(n385), .B1(n384), .B2(n546), .ZN(n307) );
  OAI22_X1 U781 ( .A1(n12), .A2(n382), .B1(n381), .B2(n502), .ZN(n304) );
  OAI22_X1 U782 ( .A1(n12), .A2(n381), .B1(n380), .B2(n508), .ZN(n303) );
  NAND2_X1 U783 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U784 ( .A1(n529), .A2(n383), .B1(n575), .B2(n382), .ZN(n305) );
  OAI22_X1 U785 ( .A1(n529), .A2(n384), .B1(n383), .B2(n575), .ZN(n306) );
  OAI22_X1 U786 ( .A1(n529), .A2(n386), .B1(n385), .B2(n575), .ZN(n308) );
  OAI22_X1 U787 ( .A1(n12), .A2(n387), .B1(n386), .B2(n575), .ZN(n309) );
  OAI22_X1 U788 ( .A1(n12), .A2(n497), .B1(n392), .B2(n508), .ZN(n257) );
  OAI22_X1 U789 ( .A1(n529), .A2(n389), .B1(n388), .B2(n575), .ZN(n311) );
  OAI22_X1 U790 ( .A1(n12), .A2(n388), .B1(n387), .B2(n575), .ZN(n310) );
  OAI22_X1 U791 ( .A1(n12), .A2(n390), .B1(n389), .B2(n575), .ZN(n312) );
  INV_X1 U792 ( .A(n575), .ZN(n247) );
  OAI22_X1 U793 ( .A1(n12), .A2(n391), .B1(n390), .B2(n575), .ZN(n313) );
  INV_X1 U794 ( .A(n31), .ZN(n596) );
  INV_X1 U795 ( .A(n36), .ZN(n598) );
  INV_X1 U796 ( .A(n600), .ZN(n599) );
  INV_X1 U797 ( .A(n40), .ZN(n600) );
  XOR2_X1 U798 ( .A(n259), .B(n251), .Z(n148) );
  XOR2_X1 U799 ( .A(n289), .B(n279), .Z(n146) );
  XOR2_X1 U800 ( .A(n149), .B(n147), .Z(n144) );
  XOR2_X1 U801 ( .A(n159), .B(n150), .Z(n142) );
endmodule


module layer1_8_4_8_16_datapath_M8_N4_T16_P8_2_DW01_add_2 ( A, B, CI, SUM, CO
 );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n18,
         n19, n20, n21, n23, n25, n26, n27, n28, n30, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n46, n48, n49, n51, n53, n54, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n71, n72, n73,
         n74, n75, n77, n79, n80, n81, n82, n83, n85, n87, n88, n90, n93, n94,
         n98, n99, n100, n102, n104, n161, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178;

  OR2_X2 U126 ( .A1(A[10]), .A2(B[10]), .ZN(n178) );
  OR2_X1 U127 ( .A1(A[11]), .A2(B[11]), .ZN(n161) );
  AND2_X1 U128 ( .A1(n172), .A2(n90), .ZN(SUM[0]) );
  OR2_X1 U129 ( .A1(A[15]), .A2(B[15]), .ZN(n163) );
  AOI21_X2 U130 ( .B1(n175), .B2(n72), .A(n69), .ZN(n67) );
  XNOR2_X1 U131 ( .A(n41), .B(n164), .ZN(SUM[11]) );
  AND2_X1 U132 ( .A1(n161), .A2(n40), .ZN(n164) );
  AOI21_X1 U133 ( .B1(n56), .B2(n64), .A(n57), .ZN(n165) );
  AOI21_X1 U134 ( .B1(n178), .B2(n51), .A(n46), .ZN(n166) );
  AOI21_X1 U135 ( .B1(n56), .B2(n64), .A(n57), .ZN(n167) );
  NOR2_X2 U136 ( .A1(A[8]), .A2(B[8]), .ZN(n58) );
  OAI21_X1 U137 ( .B1(n43), .B2(n167), .A(n44), .ZN(n168) );
  NOR2_X1 U138 ( .A1(A[12]), .A2(B[12]), .ZN(n169) );
  NOR2_X1 U139 ( .A1(A[12]), .A2(B[12]), .ZN(n36) );
  AOI21_X1 U140 ( .B1(n168), .B2(n34), .A(n35), .ZN(n170) );
  AOI21_X1 U141 ( .B1(n42), .B2(n34), .A(n35), .ZN(n171) );
  OR2_X1 U142 ( .A1(A[0]), .A2(B[0]), .ZN(n172) );
  INV_X1 U143 ( .A(n64), .ZN(n63) );
  INV_X1 U144 ( .A(n165), .ZN(n54) );
  INV_X1 U145 ( .A(n48), .ZN(n46) );
  INV_X1 U146 ( .A(n71), .ZN(n69) );
  AOI21_X1 U147 ( .B1(n176), .B2(n80), .A(n77), .ZN(n75) );
  INV_X1 U148 ( .A(n79), .ZN(n77) );
  AOI21_X1 U149 ( .B1(n174), .B2(n88), .A(n85), .ZN(n83) );
  INV_X1 U150 ( .A(n87), .ZN(n85) );
  INV_X1 U151 ( .A(n28), .ZN(n30) );
  OAI21_X1 U152 ( .B1(n83), .B2(n81), .A(n82), .ZN(n80) );
  AOI21_X1 U153 ( .B1(n54), .B2(n173), .A(n51), .ZN(n49) );
  NAND2_X1 U154 ( .A1(n98), .A2(n59), .ZN(n8) );
  INV_X1 U155 ( .A(n90), .ZN(n88) );
  OAI21_X1 U156 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  INV_X1 U157 ( .A(n53), .ZN(n51) );
  INV_X1 U158 ( .A(n27), .ZN(n93) );
  NAND2_X1 U159 ( .A1(n173), .A2(n53), .ZN(n7) );
  NAND2_X1 U160 ( .A1(n176), .A2(n79), .ZN(n13) );
  NAND2_X1 U161 ( .A1(n99), .A2(n62), .ZN(n9) );
  INV_X1 U162 ( .A(n61), .ZN(n99) );
  NAND2_X1 U163 ( .A1(n104), .A2(n82), .ZN(n14) );
  INV_X1 U164 ( .A(n81), .ZN(n104) );
  NAND2_X1 U165 ( .A1(n100), .A2(n66), .ZN(n10) );
  INV_X1 U166 ( .A(n65), .ZN(n100) );
  NAND2_X1 U167 ( .A1(n102), .A2(n74), .ZN(n12) );
  INV_X1 U168 ( .A(n73), .ZN(n102) );
  NAND2_X1 U169 ( .A1(n175), .A2(n71), .ZN(n11) );
  NAND2_X1 U170 ( .A1(n174), .A2(n87), .ZN(n15) );
  INV_X1 U171 ( .A(n25), .ZN(n23) );
  NAND2_X1 U172 ( .A1(n37), .A2(n94), .ZN(n4) );
  XNOR2_X1 U173 ( .A(n54), .B(n7), .ZN(SUM[9]) );
  XOR2_X1 U174 ( .A(n63), .B(n9), .Z(SUM[7]) );
  XNOR2_X1 U175 ( .A(n13), .B(n80), .ZN(SUM[3]) );
  XNOR2_X1 U176 ( .A(n15), .B(n88), .ZN(SUM[1]) );
  NOR2_X1 U177 ( .A1(A[11]), .A2(B[11]), .ZN(n39) );
  NOR2_X1 U178 ( .A1(A[7]), .A2(B[7]), .ZN(n61) );
  NAND2_X1 U179 ( .A1(n93), .A2(n28), .ZN(n3) );
  OR2_X1 U180 ( .A1(A[9]), .A2(B[9]), .ZN(n173) );
  NOR2_X1 U181 ( .A1(A[2]), .A2(B[2]), .ZN(n81) );
  NAND2_X1 U182 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  XOR2_X1 U183 ( .A(n49), .B(n6), .Z(SUM[10]) );
  NAND2_X1 U184 ( .A1(A[11]), .A2(B[11]), .ZN(n40) );
  OR2_X1 U185 ( .A1(A[1]), .A2(B[1]), .ZN(n174) );
  NAND2_X1 U186 ( .A1(A[12]), .A2(B[12]), .ZN(n37) );
  XNOR2_X1 U187 ( .A(n60), .B(n8), .ZN(SUM[8]) );
  NOR2_X1 U188 ( .A1(A[4]), .A2(B[4]), .ZN(n73) );
  NOR2_X1 U189 ( .A1(A[6]), .A2(B[6]), .ZN(n65) );
  NAND2_X1 U190 ( .A1(A[7]), .A2(B[7]), .ZN(n62) );
  OR2_X1 U191 ( .A1(A[5]), .A2(B[5]), .ZN(n175) );
  NAND2_X1 U192 ( .A1(A[2]), .A2(B[2]), .ZN(n82) );
  OR2_X1 U193 ( .A1(A[3]), .A2(B[3]), .ZN(n176) );
  NAND2_X1 U194 ( .A1(A[15]), .A2(B[15]), .ZN(n18) );
  NAND2_X1 U195 ( .A1(A[5]), .A2(B[5]), .ZN(n71) );
  NAND2_X1 U196 ( .A1(A[1]), .A2(B[1]), .ZN(n87) );
  NAND2_X1 U197 ( .A1(A[0]), .A2(B[0]), .ZN(n90) );
  NAND2_X1 U198 ( .A1(A[4]), .A2(B[4]), .ZN(n74) );
  NAND2_X1 U199 ( .A1(A[6]), .A2(B[6]), .ZN(n66) );
  OR2_X1 U200 ( .A1(A[14]), .A2(B[14]), .ZN(n177) );
  NAND2_X1 U201 ( .A1(A[14]), .A2(B[14]), .ZN(n25) );
  XOR2_X1 U202 ( .A(n10), .B(n67), .Z(SUM[6]) );
  XNOR2_X1 U203 ( .A(n11), .B(n72), .ZN(SUM[5]) );
  XOR2_X1 U204 ( .A(n12), .B(n75), .Z(SUM[4]) );
  XOR2_X1 U205 ( .A(n14), .B(n83), .Z(SUM[2]) );
  INV_X1 U206 ( .A(n168), .ZN(n41) );
  NAND2_X1 U207 ( .A1(A[9]), .A2(B[9]), .ZN(n53) );
  NOR2_X1 U208 ( .A1(A[13]), .A2(B[13]), .ZN(n27) );
  NAND2_X1 U209 ( .A1(n163), .A2(n18), .ZN(n1) );
  OAI21_X1 U210 ( .B1(n41), .B2(n39), .A(n40), .ZN(n38) );
  OAI21_X1 U211 ( .B1(n36), .B2(n40), .A(n37), .ZN(n35) );
  NOR2_X1 U212 ( .A1(n169), .A2(n39), .ZN(n34) );
  INV_X1 U213 ( .A(n169), .ZN(n94) );
  INV_X1 U214 ( .A(n58), .ZN(n98) );
  NOR2_X1 U215 ( .A1(n58), .A2(n61), .ZN(n56) );
  OAI21_X1 U216 ( .B1(n58), .B2(n62), .A(n59), .ZN(n57) );
  NAND2_X1 U217 ( .A1(A[8]), .A2(B[8]), .ZN(n59) );
  AOI21_X1 U218 ( .B1(n177), .B2(n30), .A(n23), .ZN(n21) );
  NAND2_X1 U219 ( .A1(n177), .A2(n93), .ZN(n20) );
  NAND2_X1 U220 ( .A1(n177), .A2(n25), .ZN(n2) );
  NAND2_X1 U221 ( .A1(A[3]), .A2(B[3]), .ZN(n79) );
  OAI21_X1 U222 ( .B1(n75), .B2(n73), .A(n74), .ZN(n72) );
  OAI21_X1 U223 ( .B1(n67), .B2(n65), .A(n66), .ZN(n64) );
  XNOR2_X1 U224 ( .A(n19), .B(n1), .ZN(SUM[15]) );
  NAND2_X1 U225 ( .A1(n178), .A2(n48), .ZN(n6) );
  OAI21_X1 U226 ( .B1(n43), .B2(n167), .A(n166), .ZN(n42) );
  NAND2_X1 U227 ( .A1(n178), .A2(n173), .ZN(n43) );
  AOI21_X1 U228 ( .B1(n178), .B2(n51), .A(n46), .ZN(n44) );
  XNOR2_X1 U229 ( .A(n38), .B(n4), .ZN(SUM[12]) );
  XNOR2_X1 U230 ( .A(n26), .B(n2), .ZN(SUM[14]) );
  XOR2_X1 U231 ( .A(n170), .B(n3), .Z(SUM[13]) );
  OAI21_X1 U232 ( .B1(n171), .B2(n27), .A(n28), .ZN(n26) );
  OAI21_X1 U233 ( .B1(n170), .B2(n20), .A(n21), .ZN(n19) );
  NAND2_X1 U234 ( .A1(A[10]), .A2(B[10]), .ZN(n48) );
endmodule


module layer1_8_4_8_16_datapath_M8_N4_T16_P8_2 ( clk, clear_acc, data_out_x, 
        data_out, data_out_w, data_out_b, wr_en_y, m_valid, m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [3:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N27, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, n1, n2, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n87, n104, n113, n114, n115, n116, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n12), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n217), .CK(clk), .Q(n17) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n218), .CK(clk), .Q(n18) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n219), .CK(clk), .Q(n19) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n220), .CK(clk), .Q(n20) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n221), .CK(clk), .Q(n21) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n222), .CK(clk), .Q(n22) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n223), .CK(clk), .Q(n23) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n224), .CK(clk), .Q(n24) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n225), .CK(clk), .Q(n25) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n226), .CK(clk), .Q(n26) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n227), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n228), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n229), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n230), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n231), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n232), .CK(clk), .Q(n35) );
  DFF_X1 \f_reg[0]  ( .D(n85), .CK(clk), .Q(n58), .QN(n206) );
  DFF_X1 \f_reg[1]  ( .D(n84), .CK(clk), .Q(n56), .QN(n207) );
  DFF_X1 \f_reg[2]  ( .D(n83), .CK(clk), .Q(n54), .QN(n208) );
  DFF_X1 \f_reg[3]  ( .D(n82), .CK(clk), .Q(f[3]), .QN(n62) );
  DFF_X1 \f_reg[4]  ( .D(n81), .CK(clk), .Q(f[4]), .QN(n63) );
  DFF_X1 \f_reg[5]  ( .D(n80), .CK(clk), .Q(f[5]), .QN(n64) );
  DFF_X1 \f_reg[6]  ( .D(n79), .CK(clk), .Q(f[6]), .QN(n65) );
  DFF_X1 \f_reg[7]  ( .D(n78), .CK(clk), .Q(f[7]), .QN(n209) );
  DFF_X1 \f_reg[8]  ( .D(n77), .CK(clk), .Q(f[8]), .QN(n210) );
  DFF_X1 \f_reg[9]  ( .D(n76), .CK(clk), .Q(f[9]), .QN(n211) );
  DFF_X1 \f_reg[10]  ( .D(n75), .CK(clk), .Q(n46), .QN(n212) );
  DFF_X1 \f_reg[11]  ( .D(n74), .CK(clk), .Q(n44), .QN(n213) );
  DFF_X1 \f_reg[12]  ( .D(n73), .CK(clk), .Q(n42), .QN(n214) );
  DFF_X1 \f_reg[13]  ( .D(n72), .CK(clk), .Q(n40), .QN(n215) );
  DFF_X1 \f_reg[14]  ( .D(n1), .CK(clk), .Q(n39), .QN(n216) );
  DFF_X1 \f_reg[15]  ( .D(n6), .CK(clk), .Q(f[15]), .QN(n70) );
  DFF_X1 \data_out_reg[15]  ( .D(n104), .CK(clk), .Q(data_out[15]), .QN(n189)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n113), .CK(clk), .Q(data_out[14]), .QN(n188)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n114), .CK(clk), .Q(data_out[13]), .QN(n187)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n115), .CK(clk), .Q(data_out[12]), .QN(n186)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n116), .CK(clk), .Q(data_out[11]), .QN(n185)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n163), .CK(clk), .Q(data_out[10]), .QN(n184)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n164), .CK(clk), .Q(data_out[9]), .QN(n183) );
  DFF_X1 \data_out_reg[8]  ( .D(n165), .CK(clk), .Q(data_out[8]), .QN(n182) );
  DFF_X1 \data_out_reg[7]  ( .D(n166), .CK(clk), .Q(data_out[7]), .QN(n181) );
  DFF_X1 \data_out_reg[6]  ( .D(n167), .CK(clk), .Q(data_out[6]), .QN(n180) );
  DFF_X1 \data_out_reg[5]  ( .D(n168), .CK(clk), .Q(data_out[5]), .QN(n179) );
  DFF_X1 \data_out_reg[4]  ( .D(n169), .CK(clk), .Q(data_out[4]), .QN(n178) );
  DFF_X1 \data_out_reg[3]  ( .D(n170), .CK(clk), .Q(data_out[3]), .QN(n177) );
  DFF_X1 \data_out_reg[2]  ( .D(n171), .CK(clk), .Q(data_out[2]), .QN(n176) );
  DFF_X1 \data_out_reg[1]  ( .D(n172), .CK(clk), .Q(data_out[1]), .QN(n175) );
  DFF_X1 \data_out_reg[0]  ( .D(n173), .CK(clk), .Q(data_out[0]), .QN(n174) );
  layer1_8_4_8_16_datapath_M8_N4_T16_P8_2_DW_mult_tc_1 mult_183 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer1_8_4_8_16_datapath_M8_N4_T16_P8_2_DW01_add_2 add_184 ( .A({n196, n195, 
        n194, n193, n192, n191, n205, n204, n203, n202, n201, n200, n199, n198, 
        n197, n190}), .B({f[15], n39, n40, n42, n44, n46, f[9:3], n54, n56, 
        n58}), .CI(1'b0), .SUM(adder) );
  DFF_X2 delay_reg ( .D(N27), .CK(clk), .Q(n7), .QN(n233) );
  MUX2_X2 U3 ( .A(n22), .B(N39), .S(n233), .Z(n191) );
  MUX2_X1 U4 ( .A(N38), .B(n23), .S(n7), .Z(n205) );
  MUX2_X1 U5 ( .A(N43), .B(n18), .S(n7), .Z(n195) );
  NAND3_X1 U6 ( .A1(n4), .A2(n2), .A3(n5), .ZN(n1) );
  NAND2_X1 U8 ( .A1(data_out_b[14]), .A2(n12), .ZN(n2) );
  NAND2_X1 U9 ( .A1(adder[14]), .A2(n11), .ZN(n4) );
  NAND2_X1 U10 ( .A1(n60), .A2(n39), .ZN(n5) );
  MUX2_X2 U11 ( .A(n21), .B(N40), .S(n233), .Z(n192) );
  MUX2_X2 U12 ( .A(N41), .B(n20), .S(n7), .Z(n193) );
  NAND3_X1 U13 ( .A1(n9), .A2(n8), .A3(n10), .ZN(n6) );
  MUX2_X2 U14 ( .A(n19), .B(N42), .S(n233), .Z(n194) );
  NAND2_X1 U15 ( .A1(data_out_b[15]), .A2(n12), .ZN(n8) );
  NAND2_X1 U16 ( .A1(adder[15]), .A2(n11), .ZN(n9) );
  NAND2_X1 U17 ( .A1(n60), .A2(f[15]), .ZN(n10) );
  AND2_X2 U18 ( .A1(n38), .A2(n13), .ZN(n11) );
  INV_X1 U19 ( .A(n13), .ZN(n12) );
  INV_X1 U20 ( .A(n38), .ZN(n60) );
  INV_X1 U21 ( .A(clear_acc), .ZN(n13) );
  NAND2_X1 U22 ( .A1(n87), .A2(N27), .ZN(n235) );
  INV_X1 U23 ( .A(wr_en_y), .ZN(n87) );
  OAI22_X1 U24 ( .A1(n177), .A2(n235), .B1(n62), .B2(n234), .ZN(n170) );
  OAI22_X1 U25 ( .A1(n178), .A2(n235), .B1(n63), .B2(n234), .ZN(n169) );
  OAI22_X1 U26 ( .A1(n179), .A2(n235), .B1(n64), .B2(n234), .ZN(n168) );
  OAI22_X1 U27 ( .A1(n180), .A2(n235), .B1(n65), .B2(n234), .ZN(n167) );
  OAI22_X1 U28 ( .A1(n181), .A2(n235), .B1(n209), .B2(n234), .ZN(n166) );
  OAI22_X1 U29 ( .A1(n182), .A2(n235), .B1(n210), .B2(n234), .ZN(n165) );
  OAI22_X1 U30 ( .A1(n183), .A2(n235), .B1(n211), .B2(n234), .ZN(n164) );
  INV_X1 U31 ( .A(n16), .ZN(n34) );
  MUX2_X1 U32 ( .A(n29), .B(N32), .S(n233), .Z(n199) );
  AND3_X1 U33 ( .A1(sel[1]), .A2(sel[2]), .A3(sel[0]), .ZN(n15) );
  INV_X1 U34 ( .A(m_ready), .ZN(n14) );
  NAND2_X1 U35 ( .A1(m_valid), .A2(n14), .ZN(n36) );
  OAI21_X1 U36 ( .B1(sel[3]), .B2(n15), .A(n36), .ZN(N27) );
  NAND2_X1 U37 ( .A1(clear_acc_delay), .A2(n233), .ZN(n16) );
  MUX2_X1 U38 ( .A(n17), .B(N44), .S(n34), .Z(n217) );
  MUX2_X1 U39 ( .A(n17), .B(N44), .S(n233), .Z(n196) );
  MUX2_X1 U40 ( .A(n18), .B(N43), .S(n34), .Z(n218) );
  MUX2_X1 U41 ( .A(n19), .B(N42), .S(n34), .Z(n219) );
  MUX2_X1 U42 ( .A(n20), .B(N41), .S(n34), .Z(n220) );
  MUX2_X1 U43 ( .A(n21), .B(N40), .S(n34), .Z(n221) );
  MUX2_X1 U44 ( .A(n22), .B(N39), .S(n34), .Z(n222) );
  MUX2_X1 U45 ( .A(n23), .B(N38), .S(n34), .Z(n223) );
  MUX2_X1 U46 ( .A(n24), .B(N37), .S(n34), .Z(n224) );
  MUX2_X1 U47 ( .A(n24), .B(N37), .S(n233), .Z(n204) );
  MUX2_X1 U48 ( .A(n25), .B(N36), .S(n34), .Z(n225) );
  MUX2_X1 U49 ( .A(n25), .B(N36), .S(n233), .Z(n203) );
  MUX2_X1 U50 ( .A(n26), .B(N35), .S(n34), .Z(n226) );
  MUX2_X1 U51 ( .A(n26), .B(N35), .S(n233), .Z(n202) );
  MUX2_X1 U52 ( .A(n27), .B(N34), .S(n34), .Z(n227) );
  MUX2_X1 U53 ( .A(n27), .B(N34), .S(n233), .Z(n201) );
  MUX2_X1 U54 ( .A(n28), .B(N33), .S(n34), .Z(n228) );
  MUX2_X1 U55 ( .A(n28), .B(N33), .S(n233), .Z(n200) );
  MUX2_X1 U56 ( .A(n29), .B(N32), .S(n34), .Z(n229) );
  MUX2_X1 U57 ( .A(n32), .B(N31), .S(n34), .Z(n230) );
  MUX2_X1 U58 ( .A(n32), .B(N31), .S(n233), .Z(n198) );
  MUX2_X1 U59 ( .A(n33), .B(N30), .S(n34), .Z(n231) );
  MUX2_X1 U60 ( .A(n33), .B(N30), .S(n233), .Z(n197) );
  MUX2_X1 U61 ( .A(n35), .B(N29), .S(n34), .Z(n232) );
  MUX2_X1 U62 ( .A(n35), .B(N29), .S(n233), .Z(n190) );
  INV_X1 U63 ( .A(n36), .ZN(n37) );
  OAI21_X1 U64 ( .B1(n37), .B2(n7), .A(n13), .ZN(n38) );
  AOI222_X1 U65 ( .A1(data_out_b[13]), .A2(n12), .B1(adder[13]), .B2(n11), 
        .C1(n60), .C2(n40), .ZN(n41) );
  INV_X1 U66 ( .A(n41), .ZN(n72) );
  AOI222_X1 U67 ( .A1(data_out_b[12]), .A2(n12), .B1(adder[12]), .B2(n11), 
        .C1(n60), .C2(n42), .ZN(n43) );
  INV_X1 U68 ( .A(n43), .ZN(n73) );
  AOI222_X1 U69 ( .A1(data_out_b[11]), .A2(n12), .B1(adder[11]), .B2(n11), 
        .C1(n60), .C2(n44), .ZN(n45) );
  INV_X1 U70 ( .A(n45), .ZN(n74) );
  AOI222_X1 U71 ( .A1(data_out_b[10]), .A2(n12), .B1(adder[10]), .B2(n11), 
        .C1(n60), .C2(n46), .ZN(n47) );
  INV_X1 U72 ( .A(n47), .ZN(n75) );
  AOI222_X1 U73 ( .A1(data_out_b[8]), .A2(n12), .B1(adder[8]), .B2(n11), .C1(
        n60), .C2(f[8]), .ZN(n48) );
  INV_X1 U74 ( .A(n48), .ZN(n77) );
  AOI222_X1 U75 ( .A1(data_out_b[7]), .A2(n12), .B1(adder[7]), .B2(n11), .C1(
        n60), .C2(f[7]), .ZN(n49) );
  INV_X1 U76 ( .A(n49), .ZN(n78) );
  AOI222_X1 U77 ( .A1(data_out_b[6]), .A2(n12), .B1(adder[6]), .B2(n11), .C1(
        n60), .C2(f[6]), .ZN(n50) );
  INV_X1 U78 ( .A(n50), .ZN(n79) );
  AOI222_X1 U79 ( .A1(data_out_b[5]), .A2(n12), .B1(adder[5]), .B2(n11), .C1(
        n60), .C2(f[5]), .ZN(n51) );
  INV_X1 U80 ( .A(n51), .ZN(n80) );
  AOI222_X1 U81 ( .A1(data_out_b[4]), .A2(n12), .B1(adder[4]), .B2(n11), .C1(
        n60), .C2(f[4]), .ZN(n52) );
  INV_X1 U82 ( .A(n52), .ZN(n81) );
  AOI222_X1 U83 ( .A1(data_out_b[3]), .A2(n12), .B1(adder[3]), .B2(n11), .C1(
        n60), .C2(f[3]), .ZN(n53) );
  INV_X1 U84 ( .A(n53), .ZN(n82) );
  AOI222_X1 U85 ( .A1(data_out_b[2]), .A2(n12), .B1(adder[2]), .B2(n11), .C1(
        n60), .C2(n54), .ZN(n55) );
  INV_X1 U86 ( .A(n55), .ZN(n83) );
  AOI222_X1 U87 ( .A1(data_out_b[1]), .A2(n12), .B1(adder[1]), .B2(n11), .C1(
        n60), .C2(n56), .ZN(n57) );
  INV_X1 U88 ( .A(n57), .ZN(n84) );
  AOI222_X1 U89 ( .A1(data_out_b[0]), .A2(n12), .B1(adder[0]), .B2(n11), .C1(
        n60), .C2(n58), .ZN(n59) );
  INV_X1 U90 ( .A(n59), .ZN(n85) );
  AOI222_X1 U91 ( .A1(data_out_b[9]), .A2(n12), .B1(adder[9]), .B2(n11), .C1(
        n60), .C2(f[9]), .ZN(n61) );
  INV_X1 U92 ( .A(n61), .ZN(n76) );
  NOR4_X1 U93 ( .A1(n44), .A2(n42), .A3(n40), .A4(n39), .ZN(n69) );
  NOR4_X1 U94 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n46), .ZN(n68) );
  NAND4_X1 U95 ( .A1(n65), .A2(n64), .A3(n63), .A4(n62), .ZN(n66) );
  NOR4_X1 U96 ( .A1(n66), .A2(n58), .A3(n56), .A4(n54), .ZN(n67) );
  NAND3_X1 U97 ( .A1(n69), .A2(n68), .A3(n67), .ZN(n71) );
  NAND3_X1 U98 ( .A1(wr_en_y), .A2(n71), .A3(n70), .ZN(n234) );
  OAI22_X1 U99 ( .A1(n174), .A2(n235), .B1(n206), .B2(n234), .ZN(n173) );
  OAI22_X1 U100 ( .A1(n175), .A2(n235), .B1(n207), .B2(n234), .ZN(n172) );
  OAI22_X1 U101 ( .A1(n176), .A2(n235), .B1(n208), .B2(n234), .ZN(n171) );
  OAI22_X1 U102 ( .A1(n184), .A2(n235), .B1(n212), .B2(n234), .ZN(n163) );
  OAI22_X1 U103 ( .A1(n185), .A2(n235), .B1(n213), .B2(n234), .ZN(n116) );
  OAI22_X1 U104 ( .A1(n186), .A2(n235), .B1(n214), .B2(n234), .ZN(n115) );
  OAI22_X1 U105 ( .A1(n187), .A2(n235), .B1(n215), .B2(n234), .ZN(n114) );
  OAI22_X1 U106 ( .A1(n188), .A2(n235), .B1(n216), .B2(n234), .ZN(n113) );
  OAI22_X1 U107 ( .A1(n189), .A2(n235), .B1(n70), .B2(n234), .ZN(n104) );
endmodule


module layer1_8_4_8_16_datapath_M8_N4_T16_P8_1_DW_mult_tc_1 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n9, n12, n13, n16, n18, n19, n21, n23, n25, n27, n29, n31,
         n32, n34, n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n50,
         n52, n53, n54, n55, n56, n57, n58, n59, n62, n63, n64, n65, n67, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n87, n88, n89, n90, n91, n95, n96, n97, n98, n99, n101,
         n103, n104, n105, n106, n107, n111, n112, n113, n114, n115, n117,
         n119, n120, n122, n127, n131, n133, n135, n139, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n247, n249, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n418, n419, n420, n421, n422, n423, n424, n426, n427, n428, n430,
         n431, n432, n433, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U148 ( .A(n265), .B(n144), .Z(n145) );
  XOR2_X1 U150 ( .A(n271), .B(n146), .Z(n147) );
  XOR2_X1 U152 ( .A(n301), .B(n148), .Z(n149) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U162 ( .A(n170), .B(n172), .CI(n179), .CO(n165), .S(n166) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n263), .CI(n291), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n317), .B(n252), .CO(n173), .S(n174) );
  FA_X1 U167 ( .A(n180), .B(n187), .CI(n178), .CO(n175), .S(n176) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U169 ( .A(n193), .B(n282), .CI(n191), .CO(n179), .S(n180) );
  FA_X1 U170 ( .A(n268), .B(n292), .CI(n274), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U174 ( .A(n275), .B(n293), .CI(n194), .CO(n189), .S(n190) );
  HA_X1 U176 ( .A(n269), .B(n319), .CO(n193), .S(n194) );
  FA_X1 U177 ( .A(n205), .B(n200), .CI(n198), .CO(n195), .S(n196) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U179 ( .A(n276), .B(n294), .CI(n284), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n320), .B(n270), .CI(n306), .CO(n201), .S(n202) );
  FA_X1 U181 ( .A(n208), .B(n213), .CI(n206), .CO(n203), .S(n204) );
  FA_X1 U182 ( .A(n215), .B(n307), .CI(n210), .CO(n205), .S(n206) );
  FA_X1 U183 ( .A(n295), .B(n285), .CI(n254), .CO(n207), .S(n208) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U185 ( .A(n216), .B(n219), .CI(n214), .CO(n211), .S(n212) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n322), .B(n278), .CI(n308), .CO(n215), .S(n216) );
  FA_X1 U188 ( .A(n225), .B(n222), .CI(n220), .CO(n217), .S(n218) );
  FA_X1 U189 ( .A(n255), .B(n309), .CI(n297), .CO(n219), .S(n220) );
  HA_X1 U190 ( .A(n287), .B(n323), .CO(n221), .S(n222) );
  FA_X1 U192 ( .A(n324), .B(n288), .CI(n310), .CO(n225), .S(n226) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  HA_X1 U194 ( .A(n311), .B(n325), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n326), .B(n300), .CI(n312), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  XNOR2_X1 U414 ( .A(n578), .B(a[2]), .ZN(n432) );
  XOR2_X1 U415 ( .A(n199), .B(n201), .Z(n490) );
  XOR2_X1 U416 ( .A(n490), .B(n192), .Z(n188) );
  XOR2_X1 U417 ( .A(n197), .B(n190), .Z(n491) );
  XOR2_X1 U418 ( .A(n491), .B(n188), .Z(n186) );
  NAND2_X1 U419 ( .A1(n199), .A2(n201), .ZN(n492) );
  NAND2_X1 U420 ( .A1(n199), .A2(n192), .ZN(n493) );
  NAND2_X1 U421 ( .A1(n201), .A2(n192), .ZN(n494) );
  NAND3_X1 U422 ( .A1(n492), .A2(n493), .A3(n494), .ZN(n187) );
  NAND2_X1 U423 ( .A1(n197), .A2(n190), .ZN(n495) );
  NAND2_X1 U424 ( .A1(n197), .A2(n188), .ZN(n496) );
  NAND2_X1 U425 ( .A1(n190), .A2(n188), .ZN(n497) );
  NAND3_X1 U426 ( .A1(n495), .A2(n496), .A3(n497), .ZN(n185) );
  XOR2_X1 U427 ( .A(n283), .B(n253), .Z(n498) );
  XOR2_X1 U428 ( .A(n305), .B(n498), .Z(n192) );
  NAND2_X1 U429 ( .A1(n305), .A2(n283), .ZN(n499) );
  NAND2_X1 U430 ( .A1(n305), .A2(n253), .ZN(n500) );
  NAND2_X1 U431 ( .A1(n283), .A2(n253), .ZN(n501) );
  NAND3_X1 U432 ( .A1(n499), .A2(n500), .A3(n501), .ZN(n191) );
  FA_X1 U433 ( .A(n216), .B(n219), .CI(n214), .S(n502) );
  INV_X2 U434 ( .A(n508), .ZN(n526) );
  BUF_X1 U435 ( .A(n573), .Z(n548) );
  NOR2_X1 U436 ( .A1(n164), .A2(n175), .ZN(n75) );
  AOI21_X1 U437 ( .B1(n564), .B2(n112), .A(n537), .ZN(n107) );
  INV_X1 U438 ( .A(n541), .ZN(n27) );
  OR2_X1 U439 ( .A1(n329), .A2(n258), .ZN(n503) );
  OR2_X2 U440 ( .A1(n212), .A2(n217), .ZN(n561) );
  AND2_X1 U441 ( .A1(n502), .A2(n217), .ZN(n504) );
  OR2_X1 U442 ( .A1(n176), .A2(n185), .ZN(n505) );
  INV_X2 U443 ( .A(n578), .ZN(n577) );
  INV_X1 U444 ( .A(n523), .ZN(n37) );
  INV_X1 U445 ( .A(n32), .ZN(n506) );
  NAND2_X1 U446 ( .A1(n196), .A2(n203), .ZN(n507) );
  XNOR2_X1 U447 ( .A(n581), .B(a[6]), .ZN(n508) );
  CLKBUF_X3 U448 ( .A(n573), .Z(n509) );
  CLKBUF_X3 U449 ( .A(n573), .Z(n510) );
  XNOR2_X1 U450 ( .A(n509), .B(b[9]), .ZN(n511) );
  NAND2_X1 U451 ( .A1(n432), .A2(n569), .ZN(n512) );
  NAND2_X1 U452 ( .A1(n432), .A2(n569), .ZN(n513) );
  XNOR2_X1 U453 ( .A(n45), .B(n514), .ZN(product[12]) );
  AND2_X1 U454 ( .A1(n505), .A2(n79), .ZN(n514) );
  XNOR2_X1 U455 ( .A(n587), .B(a[10]), .ZN(n428) );
  AOI21_X1 U456 ( .B1(n563), .B2(n120), .A(n117), .ZN(n115) );
  XOR2_X1 U457 ( .A(n7), .B(a[4]), .Z(n542) );
  XOR2_X1 U458 ( .A(n527), .B(b[10]), .Z(n398) );
  XNOR2_X1 U459 ( .A(n166), .B(n515), .ZN(n164) );
  XNOR2_X1 U460 ( .A(n177), .B(n168), .ZN(n515) );
  OAI21_X1 U461 ( .B1(n91), .B2(n89), .A(n90), .ZN(n516) );
  INV_X1 U462 ( .A(n16), .ZN(n517) );
  OR2_X2 U463 ( .A1(n518), .A2(n541), .ZN(n29) );
  XNOR2_X1 U464 ( .A(n584), .B(a[8]), .ZN(n518) );
  NAND2_X1 U465 ( .A1(n166), .A2(n177), .ZN(n519) );
  NAND2_X1 U466 ( .A1(n166), .A2(n168), .ZN(n520) );
  NAND2_X1 U467 ( .A1(n177), .A2(n168), .ZN(n521) );
  NAND3_X1 U468 ( .A1(n519), .A2(n520), .A3(n521), .ZN(n163) );
  OR2_X1 U469 ( .A1(n164), .A2(n175), .ZN(n522) );
  OAI21_X1 U470 ( .B1(n507), .B2(n82), .A(n83), .ZN(n81) );
  OAI21_X1 U471 ( .B1(n113), .B2(n115), .A(n114), .ZN(n112) );
  XNOR2_X1 U472 ( .A(n581), .B(a[4]), .ZN(n431) );
  INV_X1 U473 ( .A(n581), .ZN(n579) );
  XNOR2_X1 U474 ( .A(n587), .B(a[12]), .ZN(n523) );
  INV_X2 U475 ( .A(n587), .ZN(n586) );
  NAND2_X1 U476 ( .A1(n428), .A2(n32), .ZN(n524) );
  XNOR2_X1 U477 ( .A(n516), .B(n525), .ZN(product[10]) );
  NAND2_X1 U478 ( .A1(n533), .A2(n507), .ZN(n525) );
  INV_X1 U479 ( .A(n540), .ZN(n21) );
  INV_X1 U480 ( .A(n1), .ZN(n527) );
  CLKBUF_X1 U481 ( .A(n584), .Z(n528) );
  BUF_X2 U482 ( .A(n9), .Z(n570) );
  AOI21_X1 U483 ( .B1(n531), .B2(n80), .A(n81), .ZN(n529) );
  AOI21_X1 U484 ( .B1(n80), .B2(n531), .A(n81), .ZN(n45) );
  XOR2_X1 U485 ( .A(n575), .B(a[2]), .Z(n9) );
  INV_X1 U486 ( .A(n1), .ZN(n575) );
  AOI21_X1 U487 ( .B1(n96), .B2(n561), .A(n504), .ZN(n530) );
  AOI21_X1 U488 ( .B1(n96), .B2(n561), .A(n504), .ZN(n91) );
  OAI21_X1 U489 ( .B1(n91), .B2(n89), .A(n90), .ZN(n531) );
  INV_X2 U490 ( .A(n542), .ZN(n532) );
  INV_X1 U491 ( .A(n542), .ZN(n16) );
  BUF_X2 U492 ( .A(n9), .Z(n569) );
  INV_X1 U493 ( .A(n578), .ZN(n576) );
  OR2_X1 U494 ( .A1(n196), .A2(n203), .ZN(n533) );
  OR2_X1 U495 ( .A1(n204), .A2(n211), .ZN(n534) );
  XNOR2_X1 U496 ( .A(n583), .B(a[6]), .ZN(n430) );
  XNOR2_X1 U497 ( .A(n527), .B(n249), .ZN(n433) );
  INV_X1 U498 ( .A(n533), .ZN(n535) );
  NOR2_X1 U499 ( .A1(n196), .A2(n203), .ZN(n85) );
  INV_X2 U500 ( .A(n249), .ZN(n571) );
  NOR2_X1 U501 ( .A1(n228), .A2(n231), .ZN(n536) );
  NOR2_X1 U502 ( .A1(n228), .A2(n231), .ZN(n105) );
  INV_X2 U503 ( .A(n538), .ZN(n32) );
  AND2_X1 U504 ( .A1(n232), .A2(n233), .ZN(n537) );
  XNOR2_X1 U505 ( .A(n585), .B(a[10]), .ZN(n538) );
  XNOR2_X1 U506 ( .A(n226), .B(n539), .ZN(n224) );
  XNOR2_X1 U507 ( .A(n298), .B(n229), .ZN(n539) );
  XNOR2_X1 U508 ( .A(n581), .B(a[6]), .ZN(n540) );
  XNOR2_X1 U509 ( .A(n583), .B(a[8]), .ZN(n541) );
  NAND2_X1 U510 ( .A1(n226), .A2(n298), .ZN(n543) );
  NAND2_X1 U511 ( .A1(n226), .A2(n229), .ZN(n544) );
  NAND2_X1 U512 ( .A1(n298), .A2(n229), .ZN(n545) );
  NAND3_X1 U513 ( .A1(n543), .A2(n544), .A3(n545), .ZN(n223) );
  OAI21_X1 U514 ( .B1(n536), .B2(n107), .A(n106), .ZN(n546) );
  OAI21_X1 U515 ( .B1(n105), .B2(n107), .A(n106), .ZN(n104) );
  NOR2_X1 U516 ( .A1(n186), .A2(n195), .ZN(n547) );
  NOR2_X1 U517 ( .A1(n186), .A2(n195), .ZN(n82) );
  INV_X2 U518 ( .A(n585), .ZN(n584) );
  AOI21_X1 U519 ( .B1(n546), .B2(n562), .A(n101), .ZN(n549) );
  NAND2_X1 U520 ( .A1(n433), .A2(n571), .ZN(n550) );
  NAND2_X1 U521 ( .A1(n433), .A2(n571), .ZN(n551) );
  INV_X1 U522 ( .A(n575), .ZN(n573) );
  NAND2_X1 U523 ( .A1(n433), .A2(n571), .ZN(n6) );
  NAND2_X1 U524 ( .A1(n430), .A2(n21), .ZN(n552) );
  NAND2_X1 U525 ( .A1(n430), .A2(n21), .ZN(n553) );
  NAND2_X1 U526 ( .A1(n430), .A2(n21), .ZN(n23) );
  OAI21_X1 U527 ( .B1(n549), .B2(n97), .A(n98), .ZN(n554) );
  NAND2_X1 U528 ( .A1(n431), .A2(n16), .ZN(n555) );
  NAND2_X1 U529 ( .A1(n431), .A2(n532), .ZN(n556) );
  NAND2_X1 U530 ( .A1(n431), .A2(n16), .ZN(n18) );
  INV_X2 U531 ( .A(n583), .ZN(n582) );
  CLKBUF_X1 U532 ( .A(n45), .Z(n557) );
  NAND2_X1 U533 ( .A1(n432), .A2(n569), .ZN(n558) );
  NAND2_X1 U534 ( .A1(n432), .A2(n569), .ZN(n559) );
  NAND2_X1 U535 ( .A1(n560), .A2(n69), .ZN(n47) );
  INV_X1 U536 ( .A(n73), .ZN(n71) );
  INV_X1 U537 ( .A(n69), .ZN(n67) );
  NAND2_X1 U538 ( .A1(n73), .A2(n560), .ZN(n64) );
  INV_X1 U539 ( .A(n74), .ZN(n72) );
  NOR2_X1 U540 ( .A1(n547), .A2(n85), .ZN(n80) );
  NAND2_X1 U541 ( .A1(n127), .A2(n83), .ZN(n50) );
  INV_X1 U542 ( .A(n547), .ZN(n127) );
  NAND2_X1 U543 ( .A1(n534), .A2(n90), .ZN(n52) );
  NAND2_X1 U544 ( .A1(n522), .A2(n76), .ZN(n48) );
  OR2_X1 U545 ( .A1(n152), .A2(n163), .ZN(n560) );
  OAI21_X1 U546 ( .B1(n75), .B2(n79), .A(n76), .ZN(n74) );
  NOR2_X1 U547 ( .A1(n75), .A2(n78), .ZN(n73) );
  NAND2_X1 U548 ( .A1(n152), .A2(n163), .ZN(n69) );
  NAND2_X1 U549 ( .A1(n561), .A2(n95), .ZN(n53) );
  NOR2_X1 U550 ( .A1(n176), .A2(n185), .ZN(n78) );
  NAND2_X1 U551 ( .A1(n131), .A2(n98), .ZN(n54) );
  INV_X1 U552 ( .A(n97), .ZN(n131) );
  NAND2_X1 U553 ( .A1(n176), .A2(n185), .ZN(n79) );
  NAND2_X1 U554 ( .A1(n564), .A2(n111), .ZN(n57) );
  INV_X1 U555 ( .A(n119), .ZN(n117) );
  INV_X1 U556 ( .A(n122), .ZN(n120) );
  XNOR2_X1 U557 ( .A(n63), .B(n46), .ZN(product[15]) );
  NAND2_X1 U558 ( .A1(n565), .A2(n62), .ZN(n46) );
  AOI21_X1 U559 ( .B1(n74), .B2(n560), .A(n67), .ZN(n65) );
  XNOR2_X1 U560 ( .A(n59), .B(n120), .ZN(product[2]) );
  NAND2_X1 U561 ( .A1(n563), .A2(n119), .ZN(n59) );
  NAND2_X1 U562 ( .A1(n164), .A2(n175), .ZN(n76) );
  NAND2_X1 U563 ( .A1(n186), .A2(n195), .ZN(n83) );
  NAND2_X1 U564 ( .A1(n502), .A2(n217), .ZN(n95) );
  NAND2_X1 U565 ( .A1(n204), .A2(n211), .ZN(n90) );
  INV_X1 U566 ( .A(n113), .ZN(n135) );
  NAND2_X1 U567 ( .A1(n133), .A2(n106), .ZN(n56) );
  INV_X1 U568 ( .A(n536), .ZN(n133) );
  INV_X1 U569 ( .A(n527), .ZN(n574) );
  OR2_X1 U570 ( .A1(n224), .A2(n227), .ZN(n562) );
  OR2_X1 U571 ( .A1(n328), .A2(n314), .ZN(n563) );
  OR2_X1 U572 ( .A1(n232), .A2(n233), .ZN(n564) );
  NAND2_X1 U573 ( .A1(n218), .A2(n223), .ZN(n98) );
  NAND2_X1 U574 ( .A1(n228), .A2(n231), .ZN(n106) );
  NAND2_X1 U575 ( .A1(n151), .A2(n139), .ZN(n62) );
  NAND2_X1 U576 ( .A1(n232), .A2(n233), .ZN(n111) );
  OR2_X1 U577 ( .A1(n151), .A2(n139), .ZN(n565) );
  AND2_X1 U578 ( .A1(n503), .A2(n122), .ZN(product[1]) );
  OR2_X1 U579 ( .A1(n43), .A2(n527), .ZN(n409) );
  OR2_X1 U580 ( .A1(n43), .A2(n578), .ZN(n392) );
  OAI22_X1 U581 ( .A1(n550), .A2(n406), .B1(n405), .B2(n571), .ZN(n327) );
  OAI22_X1 U582 ( .A1(n6), .A2(n408), .B1(n407), .B2(n571), .ZN(n329) );
  OAI22_X1 U583 ( .A1(n6), .A2(n400), .B1(n511), .B2(n571), .ZN(n321) );
  XNOR2_X1 U584 ( .A(n584), .B(n43), .ZN(n352) );
  OAI22_X1 U585 ( .A1(n42), .A2(n591), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U586 ( .A1(n43), .A2(n591), .ZN(n332) );
  OAI22_X1 U587 ( .A1(n404), .A2(n551), .B1(n403), .B2(n571), .ZN(n325) );
  XOR2_X1 U588 ( .A(n315), .B(n261), .Z(n150) );
  OAI22_X1 U589 ( .A1(n6), .A2(n394), .B1(n393), .B2(n571), .ZN(n315) );
  XNOR2_X1 U590 ( .A(n155), .B(n567), .ZN(n139) );
  XNOR2_X1 U591 ( .A(n153), .B(n141), .ZN(n567) );
  XNOR2_X1 U592 ( .A(n157), .B(n568), .ZN(n141) );
  XNOR2_X1 U593 ( .A(n145), .B(n143), .ZN(n568) );
  OR2_X1 U594 ( .A1(n572), .A2(n581), .ZN(n377) );
  AND2_X1 U595 ( .A1(n572), .A2(n517), .ZN(n300) );
  OAI22_X1 U596 ( .A1(n550), .A2(n405), .B1(n404), .B2(n571), .ZN(n326) );
  XNOR2_X1 U597 ( .A(n588), .B(n43), .ZN(n336) );
  XNOR2_X1 U598 ( .A(n580), .B(n572), .ZN(n376) );
  OAI22_X1 U599 ( .A1(n39), .A2(n336), .B1(n37), .B2(n335), .ZN(n263) );
  INV_X1 U600 ( .A(n19), .ZN(n583) );
  INV_X1 U601 ( .A(n25), .ZN(n585) );
  AND2_X1 U602 ( .A1(n572), .A2(n523), .ZN(n264) );
  OAI22_X1 U603 ( .A1(n550), .A2(n397), .B1(n396), .B2(n571), .ZN(n318) );
  AND2_X1 U604 ( .A1(n572), .A2(n508), .ZN(n288) );
  OAI22_X1 U605 ( .A1(n550), .A2(n403), .B1(n402), .B2(n571), .ZN(n324) );
  AND2_X1 U606 ( .A1(n572), .A2(n506), .ZN(n270) );
  OAI22_X1 U607 ( .A1(n399), .A2(n551), .B1(n398), .B2(n571), .ZN(n320) );
  AND2_X1 U608 ( .A1(n572), .A2(n235), .ZN(n260) );
  OAI22_X1 U609 ( .A1(n550), .A2(n395), .B1(n394), .B2(n571), .ZN(n316) );
  OAI22_X1 U610 ( .A1(n39), .A2(n335), .B1(n37), .B2(n334), .ZN(n262) );
  INV_X1 U611 ( .A(n13), .ZN(n581) );
  AND2_X1 U612 ( .A1(n572), .A2(n541), .ZN(n278) );
  OAI22_X1 U613 ( .A1(n6), .A2(n401), .B1(n400), .B2(n571), .ZN(n322) );
  INV_X1 U614 ( .A(n7), .ZN(n578) );
  INV_X1 U615 ( .A(n41), .ZN(n235) );
  OAI22_X1 U616 ( .A1(n551), .A2(n398), .B1(n397), .B2(n571), .ZN(n319) );
  XNOR2_X1 U617 ( .A(n586), .B(n43), .ZN(n343) );
  OAI22_X1 U618 ( .A1(n6), .A2(n402), .B1(n401), .B2(n571), .ZN(n323) );
  XNOR2_X1 U619 ( .A(n582), .B(n43), .ZN(n363) );
  OAI22_X1 U620 ( .A1(n550), .A2(n396), .B1(n395), .B2(n571), .ZN(n317) );
  OAI22_X1 U621 ( .A1(n39), .A2(n589), .B1(n337), .B2(n37), .ZN(n252) );
  OR2_X1 U622 ( .A1(n43), .A2(n589), .ZN(n337) );
  AND2_X1 U623 ( .A1(n572), .A2(n247), .ZN(n314) );
  AND2_X1 U624 ( .A1(n572), .A2(n249), .ZN(product[0]) );
  OR2_X1 U625 ( .A1(n43), .A2(n587), .ZN(n344) );
  OR2_X1 U626 ( .A1(n43), .A2(n583), .ZN(n364) );
  OR2_X1 U627 ( .A1(n43), .A2(n585), .ZN(n353) );
  XNOR2_X1 U628 ( .A(n588), .B(a[14]), .ZN(n41) );
  NAND2_X1 U629 ( .A1(n569), .A2(n432), .ZN(n12) );
  OAI22_X1 U630 ( .A1(n39), .A2(n334), .B1(n37), .B2(n333), .ZN(n261) );
  XNOR2_X1 U631 ( .A(n588), .B(n422), .ZN(n333) );
  XNOR2_X1 U632 ( .A(n580), .B(b[11]), .ZN(n365) );
  XNOR2_X1 U633 ( .A(n582), .B(b[9]), .ZN(n354) );
  OAI22_X1 U634 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U635 ( .A(n590), .B(n424), .ZN(n330) );
  XNOR2_X1 U636 ( .A(n590), .B(n43), .ZN(n331) );
  XNOR2_X1 U637 ( .A(n588), .B(n424), .ZN(n335) );
  XNOR2_X1 U638 ( .A(n574), .B(b[11]), .ZN(n397) );
  XNOR2_X1 U639 ( .A(n574), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U640 ( .A(n574), .B(b[13]), .ZN(n395) );
  XNOR2_X1 U641 ( .A(n574), .B(b[14]), .ZN(n394) );
  XNOR2_X1 U642 ( .A(n528), .B(n418), .ZN(n345) );
  XNOR2_X1 U643 ( .A(n586), .B(n420), .ZN(n338) );
  XNOR2_X1 U644 ( .A(n577), .B(b[13]), .ZN(n378) );
  NAND2_X1 U645 ( .A1(n427), .A2(n37), .ZN(n39) );
  XNOR2_X1 U646 ( .A(n582), .B(n424), .ZN(n362) );
  XNOR2_X1 U647 ( .A(n586), .B(n424), .ZN(n342) );
  XNOR2_X1 U648 ( .A(n584), .B(n424), .ZN(n351) );
  XNOR2_X1 U649 ( .A(n577), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U650 ( .A(n577), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U651 ( .A(n577), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U652 ( .A(n577), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U653 ( .A(n577), .B(n418), .ZN(n384) );
  XNOR2_X1 U654 ( .A(n577), .B(n419), .ZN(n385) );
  XNOR2_X1 U655 ( .A(n577), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U656 ( .A(n586), .B(n422), .ZN(n340) );
  XNOR2_X1 U657 ( .A(n586), .B(n421), .ZN(n339) );
  XNOR2_X1 U658 ( .A(n580), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U659 ( .A(n580), .B(n418), .ZN(n369) );
  XNOR2_X1 U660 ( .A(n580), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U661 ( .A(n580), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U662 ( .A(n582), .B(n422), .ZN(n360) );
  XNOR2_X1 U663 ( .A(n584), .B(n422), .ZN(n349) );
  XNOR2_X1 U664 ( .A(n582), .B(n421), .ZN(n359) );
  XNOR2_X1 U665 ( .A(n582), .B(n420), .ZN(n358) );
  XNOR2_X1 U666 ( .A(n584), .B(n420), .ZN(n347) );
  XNOR2_X1 U667 ( .A(n584), .B(n421), .ZN(n348) );
  XNOR2_X1 U668 ( .A(n582), .B(n418), .ZN(n356) );
  XNOR2_X1 U669 ( .A(n582), .B(n419), .ZN(n357) );
  XNOR2_X1 U670 ( .A(n528), .B(n419), .ZN(n346) );
  XNOR2_X1 U671 ( .A(n582), .B(b[8]), .ZN(n355) );
  XNOR2_X1 U672 ( .A(n574), .B(b[15]), .ZN(n393) );
  NAND2_X1 U673 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U674 ( .A(n590), .B(a[14]), .Z(n426) );
  XNOR2_X1 U675 ( .A(n588), .B(n423), .ZN(n334) );
  BUF_X1 U676 ( .A(n43), .Z(n572) );
  XNOR2_X1 U677 ( .A(n586), .B(n423), .ZN(n341) );
  XNOR2_X1 U678 ( .A(n584), .B(n423), .ZN(n350) );
  XNOR2_X1 U679 ( .A(n582), .B(n423), .ZN(n361) );
  OAI22_X1 U680 ( .A1(n524), .A2(n339), .B1(n338), .B2(n32), .ZN(n265) );
  OAI22_X1 U681 ( .A1(n34), .A2(n340), .B1(n339), .B2(n32), .ZN(n266) );
  OAI22_X1 U682 ( .A1(n34), .A2(n342), .B1(n341), .B2(n32), .ZN(n268) );
  OAI22_X1 U683 ( .A1(n524), .A2(n341), .B1(n340), .B2(n32), .ZN(n267) );
  OAI22_X1 U684 ( .A1(n524), .A2(n343), .B1(n342), .B2(n32), .ZN(n269) );
  OAI22_X1 U685 ( .A1(n34), .A2(n587), .B1(n344), .B2(n32), .ZN(n253) );
  NAND2_X1 U686 ( .A1(n428), .A2(n32), .ZN(n34) );
  XOR2_X1 U687 ( .A(n588), .B(a[12]), .Z(n427) );
  NAND2_X1 U688 ( .A1(n328), .A2(n314), .ZN(n119) );
  OAI22_X1 U689 ( .A1(n6), .A2(n407), .B1(n406), .B2(n571), .ZN(n328) );
  XNOR2_X1 U690 ( .A(n576), .B(n43), .ZN(n391) );
  XNOR2_X1 U691 ( .A(n576), .B(n420), .ZN(n386) );
  XNOR2_X1 U692 ( .A(n576), .B(n422), .ZN(n388) );
  XNOR2_X1 U693 ( .A(n576), .B(n424), .ZN(n390) );
  XNOR2_X1 U694 ( .A(n576), .B(n423), .ZN(n389) );
  XNOR2_X1 U695 ( .A(n576), .B(n421), .ZN(n387) );
  NOR2_X1 U696 ( .A1(n218), .A2(n223), .ZN(n97) );
  OAI21_X1 U697 ( .B1(n87), .B2(n535), .A(n507), .ZN(n84) );
  XNOR2_X1 U698 ( .A(n70), .B(n47), .ZN(product[14]) );
  NAND2_X1 U699 ( .A1(n329), .A2(n258), .ZN(n122) );
  OAI22_X1 U700 ( .A1(n551), .A2(n527), .B1(n409), .B2(n571), .ZN(n258) );
  NOR2_X1 U701 ( .A1(n234), .A2(n257), .ZN(n113) );
  NAND2_X1 U702 ( .A1(n562), .A2(n103), .ZN(n55) );
  NAND2_X1 U703 ( .A1(n224), .A2(n227), .ZN(n103) );
  NOR2_X1 U704 ( .A1(n204), .A2(n211), .ZN(n89) );
  OAI22_X1 U705 ( .A1(n29), .A2(n346), .B1(n345), .B2(n27), .ZN(n271) );
  OAI22_X1 U706 ( .A1(n29), .A2(n350), .B1(n349), .B2(n27), .ZN(n275) );
  OAI22_X1 U707 ( .A1(n29), .A2(n347), .B1(n346), .B2(n27), .ZN(n272) );
  OAI22_X1 U708 ( .A1(n29), .A2(n351), .B1(n350), .B2(n27), .ZN(n276) );
  OAI22_X1 U709 ( .A1(n29), .A2(n348), .B1(n347), .B2(n27), .ZN(n273) );
  OAI22_X1 U710 ( .A1(n29), .A2(n349), .B1(n348), .B2(n27), .ZN(n274) );
  OAI22_X1 U711 ( .A1(n29), .A2(n585), .B1(n353), .B2(n27), .ZN(n254) );
  OAI22_X1 U712 ( .A1(n29), .A2(n352), .B1(n351), .B2(n27), .ZN(n277) );
  XNOR2_X1 U713 ( .A(n77), .B(n48), .ZN(product[13]) );
  OAI22_X1 U714 ( .A1(n553), .A2(n358), .B1(n357), .B2(n526), .ZN(n282) );
  OAI22_X1 U715 ( .A1(n552), .A2(n356), .B1(n355), .B2(n526), .ZN(n280) );
  OAI22_X1 U716 ( .A1(n553), .A2(n362), .B1(n361), .B2(n526), .ZN(n286) );
  OAI22_X1 U717 ( .A1(n552), .A2(n357), .B1(n356), .B2(n526), .ZN(n281) );
  OAI22_X1 U718 ( .A1(n553), .A2(n360), .B1(n359), .B2(n526), .ZN(n284) );
  OAI22_X1 U719 ( .A1(n552), .A2(n583), .B1(n364), .B2(n526), .ZN(n255) );
  OAI22_X1 U720 ( .A1(n553), .A2(n361), .B1(n360), .B2(n526), .ZN(n285) );
  OAI22_X1 U721 ( .A1(n23), .A2(n363), .B1(n526), .B2(n362), .ZN(n287) );
  OAI22_X1 U722 ( .A1(n23), .A2(n359), .B1(n358), .B2(n21), .ZN(n283) );
  OAI22_X1 U723 ( .A1(n552), .A2(n355), .B1(n354), .B2(n526), .ZN(n279) );
  XOR2_X1 U724 ( .A(n58), .B(n115), .Z(product[3]) );
  XNOR2_X1 U725 ( .A(n579), .B(n424), .ZN(n375) );
  XNOR2_X1 U726 ( .A(n579), .B(n419), .ZN(n370) );
  XNOR2_X1 U727 ( .A(n579), .B(n423), .ZN(n374) );
  XNOR2_X1 U728 ( .A(n579), .B(n420), .ZN(n371) );
  XNOR2_X1 U729 ( .A(n579), .B(n422), .ZN(n373) );
  XNOR2_X1 U730 ( .A(n579), .B(n421), .ZN(n372) );
  XOR2_X1 U731 ( .A(n549), .B(n54), .Z(product[7]) );
  AOI21_X1 U732 ( .B1(n104), .B2(n562), .A(n101), .ZN(n99) );
  XNOR2_X1 U733 ( .A(n554), .B(n53), .ZN(product[8]) );
  OAI21_X1 U734 ( .B1(n99), .B2(n97), .A(n98), .ZN(n96) );
  INV_X1 U735 ( .A(n88), .ZN(n87) );
  OAI21_X1 U736 ( .B1(n530), .B2(n89), .A(n90), .ZN(n88) );
  XOR2_X1 U737 ( .A(n52), .B(n530), .Z(product[9]) );
  OAI22_X1 U738 ( .A1(n556), .A2(n370), .B1(n369), .B2(n532), .ZN(n293) );
  OAI22_X1 U739 ( .A1(n555), .A2(n367), .B1(n366), .B2(n532), .ZN(n290) );
  OAI22_X1 U740 ( .A1(n556), .A2(n368), .B1(n367), .B2(n532), .ZN(n291) );
  OAI22_X1 U741 ( .A1(n555), .A2(n372), .B1(n371), .B2(n532), .ZN(n295) );
  OAI22_X1 U742 ( .A1(n18), .A2(n369), .B1(n368), .B2(n532), .ZN(n292) );
  OAI22_X1 U743 ( .A1(n555), .A2(n375), .B1(n374), .B2(n532), .ZN(n298) );
  OAI22_X1 U744 ( .A1(n18), .A2(n371), .B1(n370), .B2(n532), .ZN(n294) );
  OAI22_X1 U745 ( .A1(n555), .A2(n373), .B1(n372), .B2(n532), .ZN(n296) );
  OAI22_X1 U746 ( .A1(n556), .A2(n581), .B1(n377), .B2(n532), .ZN(n256) );
  OAI22_X1 U747 ( .A1(n555), .A2(n376), .B1(n375), .B2(n532), .ZN(n299) );
  OAI22_X1 U748 ( .A1(n556), .A2(n366), .B1(n365), .B2(n532), .ZN(n289) );
  OAI22_X1 U749 ( .A1(n18), .A2(n374), .B1(n373), .B2(n532), .ZN(n297) );
  XNOR2_X1 U750 ( .A(n84), .B(n50), .ZN(product[11]) );
  INV_X1 U751 ( .A(n103), .ZN(n101) );
  XNOR2_X1 U752 ( .A(n55), .B(n546), .ZN(product[6]) );
  OAI21_X1 U753 ( .B1(n64), .B2(n557), .A(n65), .ZN(n63) );
  OAI21_X1 U754 ( .B1(n529), .B2(n78), .A(n79), .ZN(n77) );
  OAI21_X1 U755 ( .B1(n529), .B2(n71), .A(n72), .ZN(n70) );
  XOR2_X1 U756 ( .A(n56), .B(n107), .Z(product[5]) );
  XNOR2_X1 U757 ( .A(n57), .B(n112), .ZN(product[4]) );
  NAND2_X1 U758 ( .A1(n135), .A2(n114), .ZN(n58) );
  XNOR2_X1 U759 ( .A(n509), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U760 ( .A(n510), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U761 ( .A(n509), .B(n418), .ZN(n401) );
  XNOR2_X1 U762 ( .A(n548), .B(n420), .ZN(n403) );
  XNOR2_X1 U763 ( .A(n510), .B(n419), .ZN(n402) );
  XNOR2_X1 U764 ( .A(n548), .B(n421), .ZN(n404) );
  XNOR2_X1 U765 ( .A(n510), .B(n422), .ZN(n405) );
  XNOR2_X1 U766 ( .A(n510), .B(n423), .ZN(n406) );
  XNOR2_X1 U767 ( .A(n509), .B(n43), .ZN(n408) );
  XNOR2_X1 U768 ( .A(n548), .B(n424), .ZN(n407) );
  OAI22_X1 U769 ( .A1(n559), .A2(n379), .B1(n378), .B2(n570), .ZN(n301) );
  OAI22_X1 U770 ( .A1(n558), .A2(n380), .B1(n379), .B2(n570), .ZN(n302) );
  OAI22_X1 U771 ( .A1(n512), .A2(n385), .B1(n384), .B2(n570), .ZN(n307) );
  OAI22_X1 U772 ( .A1(n558), .A2(n382), .B1(n381), .B2(n570), .ZN(n304) );
  OAI22_X1 U773 ( .A1(n513), .A2(n381), .B1(n380), .B2(n570), .ZN(n303) );
  NAND2_X1 U774 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U775 ( .A1(n559), .A2(n383), .B1(n382), .B2(n570), .ZN(n305) );
  OAI22_X1 U776 ( .A1(n12), .A2(n384), .B1(n383), .B2(n570), .ZN(n306) );
  OAI22_X1 U777 ( .A1(n12), .A2(n386), .B1(n385), .B2(n570), .ZN(n308) );
  OAI22_X1 U778 ( .A1(n559), .A2(n387), .B1(n386), .B2(n570), .ZN(n309) );
  OAI22_X1 U779 ( .A1(n12), .A2(n578), .B1(n392), .B2(n570), .ZN(n257) );
  OAI22_X1 U780 ( .A1(n558), .A2(n389), .B1(n388), .B2(n570), .ZN(n311) );
  OAI22_X1 U781 ( .A1(n512), .A2(n388), .B1(n387), .B2(n570), .ZN(n310) );
  OAI22_X1 U782 ( .A1(n513), .A2(n390), .B1(n570), .B2(n389), .ZN(n312) );
  INV_X1 U783 ( .A(n570), .ZN(n247) );
  OAI22_X1 U784 ( .A1(n512), .A2(n391), .B1(n390), .B2(n570), .ZN(n313) );
  INV_X1 U785 ( .A(n581), .ZN(n580) );
  INV_X1 U786 ( .A(n31), .ZN(n587) );
  INV_X1 U787 ( .A(n589), .ZN(n588) );
  INV_X1 U788 ( .A(n36), .ZN(n589) );
  INV_X1 U789 ( .A(n591), .ZN(n590) );
  INV_X1 U790 ( .A(n40), .ZN(n591) );
  XOR2_X1 U791 ( .A(n259), .B(n251), .Z(n148) );
  XOR2_X1 U792 ( .A(n289), .B(n279), .Z(n146) );
  XOR2_X1 U793 ( .A(n149), .B(n147), .Z(n144) );
  XOR2_X1 U794 ( .A(n159), .B(n150), .Z(n142) );
endmodule


module layer1_8_4_8_16_datapath_M8_N4_T16_P8_1_DW01_add_2 ( A, B, CI, SUM, CO
 );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n7, n8, n9, n10, n11, n12, n13, n14, n15, n18,
         n19, n20, n21, n23, n25, n26, n27, n28, n30, n34, n35, n36, n37, n38,
         n39, n40, n42, n43, n44, n48, n49, n51, n53, n54, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n69, n71, n72, n73, n74, n75,
         n77, n79, n80, n81, n82, n83, n85, n87, n88, n90, n93, n94, n95, n98,
         n99, n100, n102, n104, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182;

  AND2_X1 U126 ( .A1(n174), .A2(n90), .ZN(SUM[0]) );
  XNOR2_X1 U127 ( .A(n49), .B(n162), .ZN(SUM[10]) );
  AND2_X1 U128 ( .A1(n181), .A2(n48), .ZN(n162) );
  AOI21_X1 U129 ( .B1(n56), .B2(n64), .A(n57), .ZN(n163) );
  AOI21_X1 U130 ( .B1(n56), .B2(n64), .A(n57), .ZN(n164) );
  NOR2_X1 U131 ( .A1(A[11]), .A2(B[11]), .ZN(n165) );
  XNOR2_X1 U132 ( .A(n42), .B(n5), .ZN(SUM[11]) );
  INV_X1 U133 ( .A(n42), .ZN(n166) );
  NOR2_X1 U134 ( .A1(A[8]), .A2(B[8]), .ZN(n167) );
  CLKBUF_X1 U135 ( .A(n27), .Z(n168) );
  AOI21_X1 U136 ( .B1(n181), .B2(n51), .A(n182), .ZN(n169) );
  OAI21_X1 U137 ( .B1(n43), .B2(n164), .A(n44), .ZN(n170) );
  NOR2_X1 U138 ( .A1(A[12]), .A2(B[12]), .ZN(n171) );
  NOR2_X1 U139 ( .A1(A[12]), .A2(B[12]), .ZN(n36) );
  OR2_X2 U140 ( .A1(A[10]), .A2(B[10]), .ZN(n181) );
  AOI21_X1 U141 ( .B1(n170), .B2(n34), .A(n35), .ZN(n172) );
  AOI21_X1 U142 ( .B1(n170), .B2(n34), .A(n35), .ZN(n173) );
  OR2_X1 U143 ( .A1(A[0]), .A2(B[0]), .ZN(n174) );
  INV_X1 U144 ( .A(n64), .ZN(n63) );
  INV_X1 U145 ( .A(n165), .ZN(n95) );
  OAI21_X1 U146 ( .B1(n75), .B2(n73), .A(n74), .ZN(n72) );
  AOI21_X1 U147 ( .B1(n180), .B2(n80), .A(n77), .ZN(n75) );
  INV_X1 U148 ( .A(n79), .ZN(n77) );
  OAI21_X1 U149 ( .B1(n67), .B2(n65), .A(n66), .ZN(n64) );
  AOI21_X1 U150 ( .B1(n175), .B2(n72), .A(n69), .ZN(n67) );
  INV_X1 U151 ( .A(n71), .ZN(n69) );
  NOR2_X1 U152 ( .A1(n167), .A2(n61), .ZN(n56) );
  OAI21_X1 U153 ( .B1(n58), .B2(n62), .A(n59), .ZN(n57) );
  OAI21_X1 U154 ( .B1(n83), .B2(n81), .A(n82), .ZN(n80) );
  AOI21_X1 U155 ( .B1(n54), .B2(n179), .A(n51), .ZN(n49) );
  INV_X1 U156 ( .A(n90), .ZN(n88) );
  OAI21_X1 U157 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  NAND2_X1 U158 ( .A1(n99), .A2(n62), .ZN(n9) );
  INV_X1 U159 ( .A(n61), .ZN(n99) );
  NAND2_X1 U160 ( .A1(n98), .A2(n59), .ZN(n8) );
  INV_X1 U161 ( .A(n167), .ZN(n98) );
  INV_X1 U162 ( .A(n27), .ZN(n93) );
  AOI21_X1 U163 ( .B1(n176), .B2(n88), .A(n85), .ZN(n83) );
  INV_X1 U164 ( .A(n87), .ZN(n85) );
  NAND2_X1 U165 ( .A1(n100), .A2(n66), .ZN(n10) );
  INV_X1 U166 ( .A(n65), .ZN(n100) );
  NAND2_X1 U167 ( .A1(n102), .A2(n74), .ZN(n12) );
  INV_X1 U168 ( .A(n73), .ZN(n102) );
  INV_X1 U169 ( .A(n171), .ZN(n94) );
  NAND2_X1 U170 ( .A1(n180), .A2(n79), .ZN(n13) );
  NAND2_X1 U171 ( .A1(n104), .A2(n82), .ZN(n14) );
  INV_X1 U172 ( .A(n81), .ZN(n104) );
  NAND2_X1 U173 ( .A1(n175), .A2(n71), .ZN(n11) );
  NAND2_X1 U174 ( .A1(n176), .A2(n87), .ZN(n15) );
  INV_X1 U175 ( .A(n25), .ZN(n23) );
  XNOR2_X1 U176 ( .A(n38), .B(n4), .ZN(SUM[12]) );
  NAND2_X1 U177 ( .A1(n94), .A2(n37), .ZN(n4) );
  XNOR2_X1 U178 ( .A(n54), .B(n7), .ZN(SUM[9]) );
  XOR2_X1 U179 ( .A(n63), .B(n9), .Z(SUM[7]) );
  XNOR2_X1 U180 ( .A(n11), .B(n72), .ZN(SUM[5]) );
  XNOR2_X1 U181 ( .A(n13), .B(n80), .ZN(SUM[3]) );
  XOR2_X1 U182 ( .A(n14), .B(n83), .Z(SUM[2]) );
  XNOR2_X1 U183 ( .A(n15), .B(n88), .ZN(SUM[1]) );
  NOR2_X1 U184 ( .A1(A[7]), .A2(B[7]), .ZN(n61) );
  NOR2_X1 U185 ( .A1(A[8]), .A2(B[8]), .ZN(n58) );
  NAND2_X1 U186 ( .A1(A[7]), .A2(B[7]), .ZN(n62) );
  NAND2_X1 U187 ( .A1(n93), .A2(n28), .ZN(n3) );
  NOR2_X1 U188 ( .A1(A[2]), .A2(B[2]), .ZN(n81) );
  OR2_X1 U189 ( .A1(A[5]), .A2(B[5]), .ZN(n175) );
  OR2_X1 U190 ( .A1(A[1]), .A2(B[1]), .ZN(n176) );
  OR2_X1 U191 ( .A1(A[14]), .A2(B[14]), .ZN(n177) );
  OR2_X1 U192 ( .A1(A[15]), .A2(B[15]), .ZN(n178) );
  NOR2_X1 U193 ( .A1(A[4]), .A2(B[4]), .ZN(n73) );
  NOR2_X1 U194 ( .A1(A[6]), .A2(B[6]), .ZN(n65) );
  OR2_X1 U195 ( .A1(A[9]), .A2(B[9]), .ZN(n179) );
  XNOR2_X1 U196 ( .A(n60), .B(n8), .ZN(SUM[8]) );
  NAND2_X1 U197 ( .A1(A[2]), .A2(B[2]), .ZN(n82) );
  OR2_X1 U198 ( .A1(A[3]), .A2(B[3]), .ZN(n180) );
  NAND2_X1 U199 ( .A1(A[1]), .A2(B[1]), .ZN(n87) );
  NAND2_X1 U200 ( .A1(A[5]), .A2(B[5]), .ZN(n71) );
  NAND2_X1 U201 ( .A1(A[0]), .A2(B[0]), .ZN(n90) );
  NAND2_X1 U202 ( .A1(A[4]), .A2(B[4]), .ZN(n74) );
  NAND2_X1 U203 ( .A1(A[6]), .A2(B[6]), .ZN(n66) );
  NAND2_X1 U204 ( .A1(A[9]), .A2(B[9]), .ZN(n53) );
  XOR2_X1 U205 ( .A(n10), .B(n67), .Z(SUM[6]) );
  XOR2_X1 U206 ( .A(n12), .B(n75), .Z(SUM[4]) );
  NAND2_X1 U207 ( .A1(A[8]), .A2(B[8]), .ZN(n59) );
  NAND2_X1 U208 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  INV_X1 U209 ( .A(n163), .ZN(n54) );
  INV_X1 U210 ( .A(n182), .ZN(n48) );
  NAND2_X1 U211 ( .A1(n179), .A2(n53), .ZN(n7) );
  INV_X1 U212 ( .A(n53), .ZN(n51) );
  NAND2_X1 U213 ( .A1(A[12]), .A2(B[12]), .ZN(n37) );
  NOR2_X1 U214 ( .A1(A[13]), .A2(B[13]), .ZN(n27) );
  INV_X1 U215 ( .A(n28), .ZN(n30) );
  AOI21_X1 U216 ( .B1(n181), .B2(n51), .A(n182), .ZN(n44) );
  NAND2_X1 U217 ( .A1(A[15]), .A2(B[15]), .ZN(n18) );
  AND2_X1 U218 ( .A1(A[10]), .A2(B[10]), .ZN(n182) );
  NAND2_X1 U219 ( .A1(A[3]), .A2(B[3]), .ZN(n79) );
  OAI21_X1 U220 ( .B1(n36), .B2(n40), .A(n37), .ZN(n35) );
  NAND2_X1 U221 ( .A1(n95), .A2(n40), .ZN(n5) );
  NAND2_X1 U222 ( .A1(A[11]), .A2(B[11]), .ZN(n40) );
  AOI21_X1 U223 ( .B1(n177), .B2(n30), .A(n23), .ZN(n21) );
  NAND2_X1 U224 ( .A1(n177), .A2(n93), .ZN(n20) );
  NAND2_X1 U225 ( .A1(n177), .A2(n25), .ZN(n2) );
  NAND2_X1 U226 ( .A1(A[14]), .A2(B[14]), .ZN(n25) );
  NOR2_X1 U227 ( .A1(A[11]), .A2(B[11]), .ZN(n39) );
  NAND2_X1 U228 ( .A1(n178), .A2(n18), .ZN(n1) );
  OAI21_X1 U229 ( .B1(n166), .B2(n165), .A(n40), .ZN(n38) );
  NOR2_X1 U230 ( .A1(n171), .A2(n39), .ZN(n34) );
  OAI21_X1 U231 ( .B1(n43), .B2(n164), .A(n169), .ZN(n42) );
  NAND2_X1 U232 ( .A1(n181), .A2(n179), .ZN(n43) );
  XNOR2_X1 U233 ( .A(n19), .B(n1), .ZN(SUM[15]) );
  XNOR2_X1 U234 ( .A(n26), .B(n2), .ZN(SUM[14]) );
  XOR2_X1 U235 ( .A(n172), .B(n3), .Z(SUM[13]) );
  OAI21_X1 U236 ( .B1(n173), .B2(n168), .A(n28), .ZN(n26) );
  OAI21_X1 U237 ( .B1(n172), .B2(n20), .A(n21), .ZN(n19) );
endmodule


module layer1_8_4_8_16_datapath_M8_N4_T16_P8_1 ( clk, clear_acc, data_out_x, 
        data_out, data_out_w, data_out_b, wr_en_y, m_valid, m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [3:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N27, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, n1, n2, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n87, n104, n113, n114, n115, n116, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n21), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n227), .CK(clk), .Q(n26) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n228), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n229), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n230), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n231), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n232), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n233), .CK(clk), .Q(n34) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n234), .CK(clk), .Q(n35) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n235), .CK(clk), .Q(n36) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n236), .CK(clk), .Q(n37) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n237), .CK(clk), .Q(n38) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n238), .CK(clk), .Q(n39) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n239), .CK(clk), .Q(n40) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n240), .CK(clk), .Q(n41) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n241), .CK(clk), .Q(n42) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n242), .CK(clk), .Q(n44) );
  DFF_X1 \f_reg[0]  ( .D(n115), .CK(clk), .Q(n65), .QN(n216) );
  DFF_X1 \f_reg[1]  ( .D(n114), .CK(clk), .Q(n63), .QN(n217) );
  DFF_X1 \f_reg[2]  ( .D(n113), .CK(clk), .Q(n61), .QN(n218) );
  DFF_X1 \f_reg[3]  ( .D(n104), .CK(clk), .Q(f[3]), .QN(n69) );
  DFF_X1 \f_reg[4]  ( .D(n87), .CK(clk), .Q(f[4]), .QN(n70) );
  DFF_X1 \f_reg[5]  ( .D(n85), .CK(clk), .Q(f[5]), .QN(n71) );
  DFF_X1 \f_reg[6]  ( .D(n84), .CK(clk), .Q(f[6]), .QN(n72) );
  DFF_X1 \f_reg[7]  ( .D(n83), .CK(clk), .Q(f[7]), .QN(n219) );
  DFF_X1 \f_reg[8]  ( .D(n82), .CK(clk), .Q(f[8]), .QN(n220) );
  DFF_X1 \f_reg[9]  ( .D(n81), .CK(clk), .Q(f[9]), .QN(n221) );
  DFF_X1 \f_reg[10]  ( .D(n80), .CK(clk), .Q(n53), .QN(n222) );
  DFF_X1 \f_reg[11]  ( .D(n79), .CK(clk), .Q(n51), .QN(n223) );
  DFF_X1 \f_reg[12]  ( .D(n6), .CK(clk), .Q(n50), .QN(n224) );
  DFF_X1 \f_reg[13]  ( .D(n1), .CK(clk), .Q(n49), .QN(n225) );
  DFF_X1 \f_reg[14]  ( .D(n7), .CK(clk), .Q(n48), .QN(n226) );
  DFF_X1 \f_reg[15]  ( .D(n11), .CK(clk), .Q(f[15]), .QN(n77) );
  DFF_X1 \data_out_reg[15]  ( .D(n168), .CK(clk), .Q(data_out[15]), .QN(n199)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n169), .CK(clk), .Q(data_out[14]), .QN(n198)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n170), .CK(clk), .Q(data_out[13]), .QN(n197)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n171), .CK(clk), .Q(data_out[12]), .QN(n196)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n172), .CK(clk), .Q(data_out[11]), .QN(n195)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n173), .CK(clk), .Q(data_out[10]), .QN(n194)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n174), .CK(clk), .Q(data_out[9]), .QN(n193) );
  DFF_X1 \data_out_reg[8]  ( .D(n175), .CK(clk), .Q(data_out[8]), .QN(n192) );
  DFF_X1 \data_out_reg[7]  ( .D(n176), .CK(clk), .Q(data_out[7]), .QN(n191) );
  DFF_X1 \data_out_reg[6]  ( .D(n177), .CK(clk), .Q(data_out[6]), .QN(n190) );
  DFF_X1 \data_out_reg[5]  ( .D(n178), .CK(clk), .Q(data_out[5]), .QN(n189) );
  DFF_X1 \data_out_reg[4]  ( .D(n179), .CK(clk), .Q(data_out[4]), .QN(n188) );
  DFF_X1 \data_out_reg[3]  ( .D(n180), .CK(clk), .Q(data_out[3]), .QN(n187) );
  DFF_X1 \data_out_reg[2]  ( .D(n181), .CK(clk), .Q(data_out[2]), .QN(n186) );
  DFF_X1 \data_out_reg[1]  ( .D(n182), .CK(clk), .Q(data_out[1]), .QN(n185) );
  DFF_X1 \data_out_reg[0]  ( .D(n183), .CK(clk), .Q(data_out[0]), .QN(n184) );
  layer1_8_4_8_16_datapath_M8_N4_T16_P8_1_DW_mult_tc_1 mult_183 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer1_8_4_8_16_datapath_M8_N4_T16_P8_1_DW01_add_2 add_184 ( .A({n206, n205, 
        n204, n203, n202, n201, n215, n214, n213, n212, n211, n210, n209, n208, 
        n207, n200}), .B({f[15], n48, n49, n50, n51, n53, f[9:3], n61, n63, 
        n65}), .CI(1'b0), .SUM(adder) );
  DFF_X2 delay_reg ( .D(N27), .CK(clk), .Q(n12), .QN(n243) );
  MUX2_X1 U3 ( .A(N39), .B(n33), .S(n12), .Z(n201) );
  MUX2_X2 U4 ( .A(N41), .B(n29), .S(n12), .Z(n203) );
  NAND3_X1 U5 ( .A1(n4), .A2(n2), .A3(n5), .ZN(n1) );
  NAND2_X1 U6 ( .A1(data_out_b[13]), .A2(n21), .ZN(n2) );
  NAND2_X1 U8 ( .A1(adder[13]), .A2(n19), .ZN(n4) );
  NAND2_X1 U9 ( .A1(n67), .A2(n49), .ZN(n5) );
  MUX2_X2 U10 ( .A(n32), .B(N40), .S(n243), .Z(n202) );
  NAND3_X1 U11 ( .A1(n9), .A2(n8), .A3(n10), .ZN(n6) );
  MUX2_X2 U12 ( .A(N43), .B(n27), .S(n12), .Z(n205) );
  MUX2_X2 U13 ( .A(n28), .B(N42), .S(n243), .Z(n204) );
  MUX2_X2 U14 ( .A(n35), .B(N37), .S(n243), .Z(n214) );
  NAND3_X1 U15 ( .A1(n14), .A2(n13), .A3(n15), .ZN(n7) );
  NAND2_X1 U16 ( .A1(data_out_b[12]), .A2(n21), .ZN(n8) );
  NAND2_X1 U17 ( .A1(adder[12]), .A2(n19), .ZN(n9) );
  NAND2_X1 U18 ( .A1(n67), .A2(n50), .ZN(n10) );
  NAND3_X1 U19 ( .A1(n17), .A2(n16), .A3(n18), .ZN(n11) );
  NAND2_X1 U20 ( .A1(data_out_b[14]), .A2(n21), .ZN(n13) );
  NAND2_X1 U21 ( .A1(adder[14]), .A2(n19), .ZN(n14) );
  NAND2_X1 U22 ( .A1(n67), .A2(n48), .ZN(n15) );
  NAND2_X1 U23 ( .A1(data_out_b[15]), .A2(n21), .ZN(n16) );
  NAND2_X1 U24 ( .A1(adder[15]), .A2(n19), .ZN(n17) );
  NAND2_X1 U25 ( .A1(n67), .A2(f[15]), .ZN(n18) );
  AND2_X2 U26 ( .A1(n47), .A2(n22), .ZN(n19) );
  INV_X1 U27 ( .A(n22), .ZN(n21) );
  INV_X1 U28 ( .A(n47), .ZN(n67) );
  INV_X1 U29 ( .A(clear_acc), .ZN(n22) );
  NAND2_X1 U30 ( .A1(n116), .A2(N27), .ZN(n245) );
  INV_X1 U31 ( .A(wr_en_y), .ZN(n116) );
  OAI22_X1 U32 ( .A1(n187), .A2(n245), .B1(n69), .B2(n244), .ZN(n180) );
  OAI22_X1 U33 ( .A1(n188), .A2(n245), .B1(n70), .B2(n244), .ZN(n179) );
  OAI22_X1 U34 ( .A1(n189), .A2(n245), .B1(n71), .B2(n244), .ZN(n178) );
  OAI22_X1 U35 ( .A1(n190), .A2(n245), .B1(n72), .B2(n244), .ZN(n177) );
  OAI22_X1 U36 ( .A1(n191), .A2(n245), .B1(n219), .B2(n244), .ZN(n176) );
  OAI22_X1 U37 ( .A1(n192), .A2(n245), .B1(n220), .B2(n244), .ZN(n175) );
  OAI22_X1 U38 ( .A1(n193), .A2(n245), .B1(n221), .B2(n244), .ZN(n174) );
  INV_X1 U39 ( .A(n25), .ZN(n43) );
  MUX2_X1 U40 ( .A(n36), .B(N36), .S(n243), .Z(n213) );
  CLKBUF_X1 U41 ( .A(N42), .Z(n20) );
  AND3_X1 U42 ( .A1(sel[1]), .A2(sel[2]), .A3(sel[0]), .ZN(n24) );
  INV_X1 U43 ( .A(m_ready), .ZN(n23) );
  NAND2_X1 U44 ( .A1(m_valid), .A2(n23), .ZN(n45) );
  OAI21_X1 U45 ( .B1(sel[3]), .B2(n24), .A(n45), .ZN(N27) );
  NAND2_X1 U46 ( .A1(clear_acc_delay), .A2(n243), .ZN(n25) );
  MUX2_X1 U47 ( .A(n26), .B(N44), .S(n43), .Z(n227) );
  MUX2_X1 U48 ( .A(n26), .B(N44), .S(n243), .Z(n206) );
  MUX2_X1 U49 ( .A(n27), .B(N43), .S(n43), .Z(n228) );
  MUX2_X1 U50 ( .A(n28), .B(n20), .S(n43), .Z(n229) );
  MUX2_X1 U51 ( .A(n29), .B(N41), .S(n43), .Z(n230) );
  MUX2_X1 U52 ( .A(n32), .B(N40), .S(n43), .Z(n231) );
  MUX2_X1 U53 ( .A(n33), .B(N39), .S(n43), .Z(n232) );
  MUX2_X1 U54 ( .A(n34), .B(N38), .S(n43), .Z(n233) );
  MUX2_X1 U55 ( .A(n34), .B(N38), .S(n243), .Z(n215) );
  MUX2_X1 U56 ( .A(n35), .B(N37), .S(n43), .Z(n234) );
  MUX2_X1 U57 ( .A(n36), .B(N36), .S(n43), .Z(n235) );
  MUX2_X1 U58 ( .A(n37), .B(N35), .S(n43), .Z(n236) );
  MUX2_X1 U59 ( .A(n37), .B(N35), .S(n243), .Z(n212) );
  MUX2_X1 U60 ( .A(n38), .B(N34), .S(n43), .Z(n237) );
  MUX2_X1 U61 ( .A(n38), .B(N34), .S(n243), .Z(n211) );
  MUX2_X1 U62 ( .A(n39), .B(N33), .S(n43), .Z(n238) );
  MUX2_X1 U63 ( .A(n39), .B(N33), .S(n243), .Z(n210) );
  MUX2_X1 U64 ( .A(n40), .B(N32), .S(n43), .Z(n239) );
  MUX2_X1 U65 ( .A(n40), .B(N32), .S(n243), .Z(n209) );
  MUX2_X1 U66 ( .A(n41), .B(N31), .S(n43), .Z(n240) );
  MUX2_X1 U67 ( .A(n41), .B(N31), .S(n243), .Z(n208) );
  MUX2_X1 U68 ( .A(n42), .B(N30), .S(n43), .Z(n241) );
  MUX2_X1 U69 ( .A(n42), .B(N30), .S(n243), .Z(n207) );
  MUX2_X1 U70 ( .A(n44), .B(N29), .S(n43), .Z(n242) );
  MUX2_X1 U71 ( .A(n44), .B(N29), .S(n243), .Z(n200) );
  INV_X1 U72 ( .A(n45), .ZN(n46) );
  OAI21_X1 U73 ( .B1(n46), .B2(n12), .A(n22), .ZN(n47) );
  AOI222_X1 U74 ( .A1(data_out_b[11]), .A2(n21), .B1(adder[11]), .B2(n19), 
        .C1(n67), .C2(n51), .ZN(n52) );
  INV_X1 U75 ( .A(n52), .ZN(n79) );
  AOI222_X1 U76 ( .A1(data_out_b[10]), .A2(n21), .B1(adder[10]), .B2(n19), 
        .C1(n67), .C2(n53), .ZN(n54) );
  INV_X1 U77 ( .A(n54), .ZN(n80) );
  AOI222_X1 U78 ( .A1(data_out_b[8]), .A2(n21), .B1(adder[8]), .B2(n19), .C1(
        n67), .C2(f[8]), .ZN(n55) );
  INV_X1 U79 ( .A(n55), .ZN(n82) );
  AOI222_X1 U80 ( .A1(data_out_b[7]), .A2(n21), .B1(adder[7]), .B2(n19), .C1(
        n67), .C2(f[7]), .ZN(n56) );
  INV_X1 U81 ( .A(n56), .ZN(n83) );
  AOI222_X1 U82 ( .A1(data_out_b[6]), .A2(n21), .B1(adder[6]), .B2(n19), .C1(
        n67), .C2(f[6]), .ZN(n57) );
  INV_X1 U83 ( .A(n57), .ZN(n84) );
  AOI222_X1 U84 ( .A1(data_out_b[5]), .A2(n21), .B1(adder[5]), .B2(n19), .C1(
        n67), .C2(f[5]), .ZN(n58) );
  INV_X1 U85 ( .A(n58), .ZN(n85) );
  AOI222_X1 U86 ( .A1(data_out_b[4]), .A2(n21), .B1(adder[4]), .B2(n19), .C1(
        n67), .C2(f[4]), .ZN(n59) );
  INV_X1 U87 ( .A(n59), .ZN(n87) );
  AOI222_X1 U88 ( .A1(data_out_b[3]), .A2(n21), .B1(adder[3]), .B2(n19), .C1(
        n67), .C2(f[3]), .ZN(n60) );
  INV_X1 U89 ( .A(n60), .ZN(n104) );
  AOI222_X1 U90 ( .A1(data_out_b[2]), .A2(n21), .B1(adder[2]), .B2(n19), .C1(
        n67), .C2(n61), .ZN(n62) );
  INV_X1 U91 ( .A(n62), .ZN(n113) );
  AOI222_X1 U92 ( .A1(data_out_b[1]), .A2(n21), .B1(adder[1]), .B2(n19), .C1(
        n67), .C2(n63), .ZN(n64) );
  INV_X1 U93 ( .A(n64), .ZN(n114) );
  AOI222_X1 U94 ( .A1(data_out_b[0]), .A2(n21), .B1(adder[0]), .B2(n19), .C1(
        n67), .C2(n65), .ZN(n66) );
  INV_X1 U95 ( .A(n66), .ZN(n115) );
  AOI222_X1 U96 ( .A1(data_out_b[9]), .A2(n21), .B1(adder[9]), .B2(n19), .C1(
        n67), .C2(f[9]), .ZN(n68) );
  INV_X1 U97 ( .A(n68), .ZN(n81) );
  NOR4_X1 U98 ( .A1(n51), .A2(n50), .A3(n49), .A4(n48), .ZN(n76) );
  NOR4_X1 U99 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n53), .ZN(n75) );
  NAND4_X1 U100 ( .A1(n72), .A2(n71), .A3(n70), .A4(n69), .ZN(n73) );
  NOR4_X1 U101 ( .A1(n73), .A2(n65), .A3(n63), .A4(n61), .ZN(n74) );
  NAND3_X1 U102 ( .A1(n76), .A2(n75), .A3(n74), .ZN(n78) );
  NAND3_X1 U103 ( .A1(wr_en_y), .A2(n78), .A3(n77), .ZN(n244) );
  OAI22_X1 U104 ( .A1(n184), .A2(n245), .B1(n216), .B2(n244), .ZN(n183) );
  OAI22_X1 U105 ( .A1(n185), .A2(n245), .B1(n217), .B2(n244), .ZN(n182) );
  OAI22_X1 U106 ( .A1(n186), .A2(n245), .B1(n218), .B2(n244), .ZN(n181) );
  OAI22_X1 U107 ( .A1(n194), .A2(n245), .B1(n222), .B2(n244), .ZN(n173) );
  OAI22_X1 U108 ( .A1(n195), .A2(n245), .B1(n223), .B2(n244), .ZN(n172) );
  OAI22_X1 U109 ( .A1(n196), .A2(n245), .B1(n224), .B2(n244), .ZN(n171) );
  OAI22_X1 U110 ( .A1(n197), .A2(n245), .B1(n225), .B2(n244), .ZN(n170) );
  OAI22_X1 U111 ( .A1(n198), .A2(n245), .B1(n226), .B2(n244), .ZN(n169) );
  OAI22_X1 U112 ( .A1(n199), .A2(n245), .B1(n77), .B2(n244), .ZN(n168) );
endmodule


module layer1_8_4_8_16_ctrlpath_M8_N4_T16_P8 ( clk, reset, s_valid, s_ready, 
        m_valid, m_ready, clear_acc, wr_en_x, wr_en_y, sel, addr_x, addr_w_0, 
        addr_b_0, addr_w_1, addr_b_1, addr_w_2, addr_b_2, addr_w_3, addr_b_3, 
        addr_w_4, addr_b_4, addr_w_5, addr_b_5, addr_w_6, addr_b_6, addr_w_7, 
        addr_b_7 );
  output [3:0] sel;
  output [2:0] addr_x;
  output [2:0] addr_w_0;
  output [0:0] addr_b_0;
  output [2:0] addr_w_1;
  output [0:0] addr_b_1;
  output [2:0] addr_w_2;
  output [0:0] addr_b_2;
  output [2:0] addr_w_3;
  output [0:0] addr_b_3;
  output [2:0] addr_w_4;
  output [0:0] addr_b_4;
  output [2:0] addr_w_5;
  output [0:0] addr_b_5;
  output [2:0] addr_w_6;
  output [0:0] addr_b_6;
  output [2:0] addr_w_7;
  output [0:0] addr_b_7;
  input clk, reset, s_valid, m_ready;
  output s_ready, m_valid, clear_acc, wr_en_x, wr_en_y;
  wire   N11, clear_acc_delay, n35, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n97, n99, n100, n101, n104, n105, n106,
         n107, n150, n151, n153, n154, n156, n158, n159, n160, n161, n167,
         n168, n169, n170, n171, n172, n173, n175, n176, n179, n180, n181,
         n182, n183, n184, n185, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n2, n3, n4, n5, n6,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n98, n102, n103, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138;
  wire   [3:0] state;

  DFF_X1 wr_en_y_reg ( .D(n223), .CK(clk), .Q(wr_en_y) );
  NAND3_X1 U144 ( .A1(addr_x[0]), .A2(n63), .A3(n119), .ZN(n156) );
  NAND3_X1 U146 ( .A1(sel[0]), .A2(n100), .A3(n126), .ZN(n171) );
  NAND3_X1 U147 ( .A1(n120), .A2(n16), .A3(n126), .ZN(n173) );
  NAND3_X1 U149 ( .A1(n175), .A2(n121), .A3(n179), .ZN(n176) );
  DFF_X1 clear_acc_delay_reg ( .D(n9), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \addr_b_7_reg[0]  ( .D(n209), .CK(clk), .Q(addr_b_7[0]), .QN(n72) );
  DFF_X1 \addr_b_6_reg[0]  ( .D(n208), .CK(clk), .Q(addr_b_6[0]), .QN(n71) );
  DFF_X1 \addr_b_5_reg[0]  ( .D(n207), .CK(clk), .Q(addr_b_5[0]), .QN(n70) );
  DFF_X1 \addr_b_4_reg[0]  ( .D(n214), .CK(clk), .Q(addr_b_4[0]), .QN(n69) );
  DFF_X1 \addr_b_3_reg[0]  ( .D(n213), .CK(clk), .Q(addr_b_3[0]), .QN(n68) );
  DFF_X1 \addr_b_2_reg[0]  ( .D(n212), .CK(clk), .Q(addr_b_2[0]), .QN(n67) );
  DFF_X1 \addr_b_1_reg[0]  ( .D(n211), .CK(clk), .Q(addr_b_1[0]), .QN(n66) );
  DFF_X1 \addr_b_0_reg[0]  ( .D(n210), .CK(clk), .Q(addr_b_0[0]), .QN(n65) );
  DFF_X1 clear_acc_reg ( .D(n136), .CK(clk), .Q(clear_acc), .QN(n35) );
  DFF_X1 m_valid_reg ( .D(n221), .CK(clk), .Q(m_valid), .QN(n97) );
  DFF_X1 \sel_count_reg[0]  ( .D(n222), .CK(clk), .Q(sel[0]), .QN(n101) );
  DFF_X1 \state_reg[1]  ( .D(n124), .CK(clk), .Q(state[1]), .QN(n60) );
  DFF_X1 \state_reg[0]  ( .D(N11), .CK(clk), .Q(state[0]), .QN(n61) );
  DFF_X1 \sel_count_reg[1]  ( .D(n219), .CK(clk), .Q(sel[1]), .QN(n100) );
  DFF_X1 \sel_count_reg[2]  ( .D(n218), .CK(clk), .Q(sel[2]), .QN(n99) );
  DFF_X1 \sel_count_reg[3]  ( .D(n220), .CK(clk), .Q(sel[3]), .QN(n16) );
  DFF_X1 \addr_w2_7_reg[0]  ( .D(n194), .CK(clk), .Q(addr_w_7[0]), .QN(n25) );
  DFF_X1 \addr_w2_6_reg[0]  ( .D(n196), .CK(clk), .Q(addr_w_6[0]), .QN(n33) );
  DFF_X1 \addr_w2_5_reg[0]  ( .D(n192), .CK(clk), .Q(addr_w_5[0]), .QN(n42) );
  DFF_X1 \addr_w2_4_reg[0]  ( .D(n198), .CK(clk), .Q(addr_w_4[0]), .QN(n50) );
  DFF_X1 \addr_w2_3_reg[0]  ( .D(n200), .CK(clk), .Q(addr_w_3[0]), .QN(n58) );
  DFF_X1 \addr_w2_2_reg[0]  ( .D(n202), .CK(clk), .Q(addr_w_2[0]), .QN(n80) );
  DFF_X1 \addr_w2_0_reg[0]  ( .D(n206), .CK(clk), .Q(addr_w_0[0]), .QN(n98) );
  DFF_X1 \addr_w2_1_reg[0]  ( .D(n204), .CK(clk), .Q(addr_w_1[0]), .QN(n88) );
  DFF_X1 \addr_x_reg[0]  ( .D(n216), .CK(clk), .Q(addr_x[0]), .QN(n64) );
  DFF_X1 \addr_w2_7_reg[1]  ( .D(n193), .CK(clk), .Q(addr_w_7[1]), .QN(n27) );
  DFF_X1 \addr_w2_6_reg[1]  ( .D(n195), .CK(clk), .Q(addr_w_6[1]), .QN(n36) );
  DFF_X1 \addr_w2_5_reg[1]  ( .D(n191), .CK(clk), .Q(addr_w_5[1]), .QN(n44) );
  DFF_X1 \addr_w2_0_reg[1]  ( .D(n205), .CK(clk), .Q(addr_w_0[1]), .QN(n103)
         );
  DFF_X1 \addr_w2_4_reg[1]  ( .D(n197), .CK(clk), .Q(addr_w_4[1]), .QN(n52) );
  DFF_X1 \addr_w2_3_reg[1]  ( .D(n199), .CK(clk), .Q(addr_w_3[1]), .QN(n74) );
  DFF_X1 \addr_w2_2_reg[1]  ( .D(n201), .CK(clk), .Q(addr_w_2[1]), .QN(n82) );
  DFF_X1 \addr_w2_1_reg[1]  ( .D(n203), .CK(clk), .Q(addr_w_1[1]), .QN(n90) );
  DFF_X1 \addr_w2_7_reg[2]  ( .D(n129), .CK(clk), .Q(addr_w_7[2]), .QN(n30) );
  DFF_X1 \addr_w2_6_reg[2]  ( .D(n130), .CK(clk), .Q(addr_w_6[2]), .QN(n39) );
  DFF_X1 \addr_w2_5_reg[2]  ( .D(n128), .CK(clk), .Q(addr_w_5[2]), .QN(n47) );
  DFF_X1 \addr_w2_0_reg[2]  ( .D(n135), .CK(clk), .Q(addr_w_0[2]), .QN(n110)
         );
  DFF_X1 \addr_w2_4_reg[2]  ( .D(n131), .CK(clk), .Q(addr_w_4[2]), .QN(n55) );
  DFF_X1 \addr_w2_3_reg[2]  ( .D(n132), .CK(clk), .Q(addr_w_3[2]), .QN(n77) );
  DFF_X1 \addr_w2_2_reg[2]  ( .D(n133), .CK(clk), .Q(addr_w_2[2]), .QN(n85) );
  DFF_X1 \addr_w2_1_reg[2]  ( .D(n134), .CK(clk), .Q(addr_w_1[2]), .QN(n93) );
  DFF_X1 \addr_x_reg[1]  ( .D(n215), .CK(clk), .Q(addr_x[1]), .QN(n63) );
  DFF_X1 \addr_x_reg[2]  ( .D(n217), .CK(clk), .Q(addr_x[2]), .QN(n62) );
  SDFF_X2 \state_reg[2]  ( .D(1'b0), .SI(n4), .SE(n121), .CK(clk), .Q(state[2]), .QN(n59) );
  AND4_X2 U3 ( .A1(m_ready), .A2(m_valid), .A3(n120), .A4(n16), .ZN(n3) );
  CLKBUF_X1 U4 ( .A(m_ready), .Z(n2) );
  AND4_X1 U5 ( .A1(m_ready), .A2(m_valid), .A3(n120), .A4(n16), .ZN(n181) );
  CLKBUF_X1 U6 ( .A(n104), .Z(n4) );
  AOI21_X1 U7 ( .B1(n187), .B2(n12), .A(n10), .ZN(n5) );
  OR3_X1 U8 ( .A1(n167), .A2(n104), .A3(n138), .ZN(n6) );
  NOR2_X1 U10 ( .A1(n35), .A2(n8), .ZN(n9) );
  INV_X1 U11 ( .A(n12), .ZN(n8) );
  OAI221_X1 U12 ( .B1(n181), .B2(n151), .C1(addr_x[2]), .C2(n183), .A(n188), 
        .ZN(n10) );
  NAND4_X4 U13 ( .A1(n151), .A2(n121), .A3(n112), .A4(n116), .ZN(n96) );
  BUF_X1 U14 ( .A(n112), .Z(n14) );
  CLKBUF_X1 U15 ( .A(n112), .Z(n15) );
  INV_X1 U16 ( .A(n11), .ZN(n136) );
  NOR3_X1 U17 ( .A1(n223), .A2(n150), .A3(n12), .ZN(n182) );
  NOR2_X1 U18 ( .A1(n180), .A2(n184), .ZN(n179) );
  OAI21_X1 U19 ( .B1(n10), .B2(n223), .A(n121), .ZN(n105) );
  INV_X1 U20 ( .A(n175), .ZN(n126) );
  AND3_X1 U21 ( .A1(n116), .A2(n121), .A3(n17), .ZN(n11) );
  NOR2_X1 U22 ( .A1(n184), .A2(n189), .ZN(n188) );
  NOR3_X1 U23 ( .A1(n190), .A2(state[0]), .A3(n138), .ZN(n189) );
  NAND2_X1 U24 ( .A1(n59), .A2(n60), .ZN(n190) );
  NOR3_X1 U25 ( .A1(n60), .A2(state[0]), .A3(n59), .ZN(n184) );
  NAND2_X1 U26 ( .A1(clear_acc_delay), .A2(n121), .ZN(n153) );
  OAI21_X1 U27 ( .B1(n63), .B2(n64), .A(n62), .ZN(n187) );
  NOR3_X1 U28 ( .A1(state[0]), .A2(state[2]), .A3(n60), .ZN(n180) );
  INV_X1 U29 ( .A(n154), .ZN(n137) );
  AOI211_X1 U30 ( .C1(state[1]), .C2(state[0]), .A(clear_acc_delay), .B(reset), 
        .ZN(n154) );
  NAND4_X1 U31 ( .A1(n179), .A2(m_valid), .A3(n2), .A4(n121), .ZN(n175) );
  OAI21_X1 U32 ( .B1(sel[1]), .B2(n175), .A(n170), .ZN(n169) );
  OAI22_X1 U33 ( .A1(n101), .A2(n176), .B1(sel[0]), .B2(n175), .ZN(n222) );
  OAI21_X1 U34 ( .B1(addr_x[0]), .B2(n123), .A(n159), .ZN(n158) );
  OAI22_X1 U35 ( .A1(n137), .A2(n69), .B1(addr_b_4[0]), .B2(n153), .ZN(n214)
         );
  OAI22_X1 U36 ( .A1(n137), .A2(n68), .B1(addr_b_3[0]), .B2(n153), .ZN(n213)
         );
  OAI22_X1 U37 ( .A1(n137), .A2(n67), .B1(addr_b_2[0]), .B2(n153), .ZN(n212)
         );
  OAI22_X1 U38 ( .A1(n137), .A2(n66), .B1(addr_b_1[0]), .B2(n153), .ZN(n211)
         );
  OAI22_X1 U39 ( .A1(n137), .A2(n65), .B1(addr_b_0[0]), .B2(n153), .ZN(n210)
         );
  OAI22_X1 U40 ( .A1(n137), .A2(n72), .B1(addr_b_7[0]), .B2(n153), .ZN(n209)
         );
  OAI22_X1 U41 ( .A1(n137), .A2(n71), .B1(addr_b_6[0]), .B2(n153), .ZN(n208)
         );
  OAI22_X1 U42 ( .A1(n137), .A2(n70), .B1(addr_b_5[0]), .B2(n153), .ZN(n207)
         );
  OAI22_X1 U43 ( .A1(n64), .A2(n159), .B1(addr_x[0]), .B2(n123), .ZN(n216) );
  AND2_X1 U44 ( .A1(n61), .A2(n13), .ZN(n12) );
  AOI21_X1 U45 ( .B1(n126), .B2(n99), .A(n169), .ZN(n172) );
  NAND4_X1 U46 ( .A1(n119), .A2(addr_x[1]), .A3(addr_x[0]), .A4(n62), .ZN(n161) );
  AOI21_X1 U47 ( .B1(n119), .B2(n63), .A(n158), .ZN(n160) );
  AND2_X1 U48 ( .A1(n13), .A2(state[0]), .ZN(n223) );
  OAI21_X1 U49 ( .B1(n170), .B2(n100), .A(n171), .ZN(n219) );
  OAI21_X1 U50 ( .B1(n4), .B2(n105), .A(n106), .ZN(s_ready) );
  NOR2_X1 U51 ( .A1(state[0]), .A2(reset), .ZN(n107) );
  NOR2_X1 U52 ( .A1(state[1]), .A2(n59), .ZN(n13) );
  NOR2_X1 U53 ( .A1(reset), .A2(n167), .ZN(N11) );
  OR3_X1 U54 ( .A1(n100), .A2(n99), .A3(n101), .ZN(n114) );
  AOI21_X1 U55 ( .B1(n101), .B2(n126), .A(n127), .ZN(n170) );
  INV_X1 U56 ( .A(n176), .ZN(n127) );
  OAI21_X1 U57 ( .B1(n125), .B2(n99), .A(n168), .ZN(n218) );
  NAND4_X1 U58 ( .A1(n126), .A2(sel[1]), .A3(sel[0]), .A4(n99), .ZN(n168) );
  INV_X1 U59 ( .A(n169), .ZN(n125) );
  OR2_X1 U60 ( .A1(n183), .A2(n62), .ZN(n116) );
  INV_X1 U61 ( .A(s_valid), .ZN(n138) );
  OAI21_X1 U62 ( .B1(n122), .B2(n63), .A(n156), .ZN(n215) );
  INV_X1 U63 ( .A(n158), .ZN(n122) );
  INV_X1 U64 ( .A(reset), .ZN(n121) );
  AOI21_X1 U65 ( .B1(n187), .B2(n12), .A(n185), .ZN(n167) );
  OAI221_X1 U66 ( .B1(n3), .B2(n151), .C1(addr_x[2]), .C2(n183), .A(n188), 
        .ZN(n185) );
  NOR3_X1 U67 ( .A1(n5), .A2(n138), .A3(n104), .ZN(wr_en_x) );
  INV_X1 U68 ( .A(n105), .ZN(n124) );
  NAND3_X1 U69 ( .A1(state[2]), .A2(state[0]), .A3(state[1]), .ZN(n151) );
  OAI211_X1 U70 ( .C1(n3), .C2(n151), .A(n179), .B(n182), .ZN(n104) );
  NAND3_X1 U71 ( .A1(n59), .A2(state[0]), .A3(state[1]), .ZN(n183) );
  OAI21_X1 U72 ( .B1(n160), .B2(n62), .A(n161), .ZN(n217) );
  INV_X1 U73 ( .A(n180), .ZN(n17) );
  OAI211_X1 U74 ( .C1(n16), .C2(n172), .A(n173), .B(n121), .ZN(n220) );
  NAND2_X1 U75 ( .A1(n114), .A2(n16), .ZN(n23) );
  NAND2_X1 U76 ( .A1(wr_en_y), .A2(n23), .ZN(n22) );
  INV_X1 U77 ( .A(n23), .ZN(n20) );
  INV_X1 U78 ( .A(n2), .ZN(n19) );
  OAI21_X1 U79 ( .B1(n20), .B2(n19), .A(m_valid), .ZN(n21) );
  AOI21_X1 U80 ( .B1(n22), .B2(n21), .A(reset), .ZN(n221) );
  OAI211_X1 U81 ( .C1(n97), .C2(m_ready), .A(n12), .B(n23), .ZN(n115) );
  INV_X1 U82 ( .A(n115), .ZN(n24) );
  NAND2_X1 U83 ( .A1(n24), .A2(n121), .ZN(n112) );
  OAI22_X1 U84 ( .A1(n25), .A2(n96), .B1(addr_w_7[0]), .B2(n112), .ZN(n194) );
  OAI21_X1 U85 ( .B1(n14), .B2(addr_w_7[0]), .A(n96), .ZN(n29) );
  NOR2_X1 U86 ( .A1(n14), .A2(n25), .ZN(n26) );
  MUX2_X1 U87 ( .A(n29), .B(n26), .S(n27), .Z(n193) );
  AND2_X1 U88 ( .A1(n30), .A2(addr_w_7[0]), .ZN(n28) );
  AOI22_X1 U89 ( .A1(n28), .A2(addr_w_7[1]), .B1(addr_w_7[2]), .B2(n27), .ZN(
        n32) );
  INV_X1 U90 ( .A(n29), .ZN(n31) );
  OAI22_X1 U91 ( .A1(n32), .A2(n15), .B1(n31), .B2(n30), .ZN(n129) );
  OAI22_X1 U92 ( .A1(n33), .A2(n96), .B1(addr_w_6[0]), .B2(n15), .ZN(n196) );
  OAI21_X1 U93 ( .B1(n14), .B2(addr_w_6[0]), .A(n96), .ZN(n38) );
  NOR2_X1 U94 ( .A1(n14), .A2(n33), .ZN(n34) );
  MUX2_X1 U95 ( .A(n38), .B(n34), .S(n36), .Z(n195) );
  AND2_X1 U96 ( .A1(n39), .A2(addr_w_6[0]), .ZN(n37) );
  AOI22_X1 U97 ( .A1(n37), .A2(addr_w_6[1]), .B1(addr_w_6[2]), .B2(n36), .ZN(
        n41) );
  INV_X1 U98 ( .A(n38), .ZN(n40) );
  OAI22_X1 U99 ( .A1(n41), .A2(n15), .B1(n40), .B2(n39), .ZN(n130) );
  OAI22_X1 U100 ( .A1(n42), .A2(n96), .B1(addr_w_5[0]), .B2(n14), .ZN(n192) );
  OAI21_X1 U101 ( .B1(n14), .B2(addr_w_5[0]), .A(n96), .ZN(n46) );
  NOR2_X1 U102 ( .A1(n14), .A2(n42), .ZN(n43) );
  MUX2_X1 U103 ( .A(n46), .B(n43), .S(n44), .Z(n191) );
  AND2_X1 U104 ( .A1(n47), .A2(addr_w_5[0]), .ZN(n45) );
  AOI22_X1 U105 ( .A1(n45), .A2(addr_w_5[1]), .B1(addr_w_5[2]), .B2(n44), .ZN(
        n49) );
  INV_X1 U106 ( .A(n46), .ZN(n48) );
  OAI22_X1 U107 ( .A1(n49), .A2(n15), .B1(n48), .B2(n47), .ZN(n128) );
  OAI22_X1 U108 ( .A1(n50), .A2(n96), .B1(addr_w_4[0]), .B2(n112), .ZN(n198)
         );
  OAI21_X1 U109 ( .B1(n14), .B2(addr_w_4[0]), .A(n96), .ZN(n54) );
  NOR2_X1 U110 ( .A1(n14), .A2(n50), .ZN(n51) );
  MUX2_X1 U111 ( .A(n54), .B(n51), .S(n52), .Z(n197) );
  AND2_X1 U112 ( .A1(n55), .A2(addr_w_4[0]), .ZN(n53) );
  AOI22_X1 U113 ( .A1(n53), .A2(addr_w_4[1]), .B1(addr_w_4[2]), .B2(n52), .ZN(
        n57) );
  INV_X1 U114 ( .A(n54), .ZN(n56) );
  OAI22_X1 U115 ( .A1(n57), .A2(n15), .B1(n56), .B2(n55), .ZN(n131) );
  OAI22_X1 U116 ( .A1(n58), .A2(n96), .B1(addr_w_3[0]), .B2(n112), .ZN(n200)
         );
  OAI21_X1 U117 ( .B1(n14), .B2(addr_w_3[0]), .A(n96), .ZN(n76) );
  NOR2_X1 U118 ( .A1(n14), .A2(n58), .ZN(n73) );
  MUX2_X1 U119 ( .A(n76), .B(n73), .S(n74), .Z(n199) );
  AND2_X1 U120 ( .A1(n77), .A2(addr_w_3[0]), .ZN(n75) );
  AOI22_X1 U121 ( .A1(n75), .A2(addr_w_3[1]), .B1(addr_w_3[2]), .B2(n74), .ZN(
        n79) );
  INV_X1 U122 ( .A(n76), .ZN(n78) );
  OAI22_X1 U123 ( .A1(n79), .A2(n15), .B1(n78), .B2(n77), .ZN(n132) );
  OAI22_X1 U124 ( .A1(n80), .A2(n96), .B1(addr_w_2[0]), .B2(n14), .ZN(n202) );
  OAI21_X1 U125 ( .B1(n14), .B2(addr_w_2[0]), .A(n96), .ZN(n84) );
  NOR2_X1 U126 ( .A1(n14), .A2(n80), .ZN(n81) );
  MUX2_X1 U127 ( .A(n84), .B(n81), .S(n82), .Z(n201) );
  AND2_X1 U128 ( .A1(n85), .A2(addr_w_2[0]), .ZN(n83) );
  AOI22_X1 U129 ( .A1(n83), .A2(addr_w_2[1]), .B1(addr_w_2[2]), .B2(n82), .ZN(
        n87) );
  INV_X1 U130 ( .A(n84), .ZN(n86) );
  OAI22_X1 U131 ( .A1(n87), .A2(n15), .B1(n86), .B2(n85), .ZN(n133) );
  OAI22_X1 U132 ( .A1(n88), .A2(n96), .B1(addr_w_1[0]), .B2(n15), .ZN(n204) );
  OAI21_X1 U133 ( .B1(n15), .B2(addr_w_1[0]), .A(n96), .ZN(n92) );
  NOR2_X1 U134 ( .A1(n14), .A2(n88), .ZN(n89) );
  MUX2_X1 U135 ( .A(n92), .B(n89), .S(n90), .Z(n203) );
  AND2_X1 U136 ( .A1(n93), .A2(addr_w_1[0]), .ZN(n91) );
  AOI22_X1 U137 ( .A1(n91), .A2(addr_w_1[1]), .B1(addr_w_1[2]), .B2(n90), .ZN(
        n95) );
  INV_X1 U138 ( .A(n92), .ZN(n94) );
  OAI22_X1 U139 ( .A1(n95), .A2(n15), .B1(n94), .B2(n93), .ZN(n134) );
  OAI22_X1 U140 ( .A1(n98), .A2(n96), .B1(addr_w_0[0]), .B2(n15), .ZN(n206) );
  OAI21_X1 U141 ( .B1(n14), .B2(addr_w_0[0]), .A(n96), .ZN(n109) );
  NOR2_X1 U142 ( .A1(n14), .A2(n98), .ZN(n102) );
  MUX2_X1 U143 ( .A(n109), .B(n102), .S(n103), .Z(n205) );
  AND2_X1 U145 ( .A1(n110), .A2(addr_w_0[0]), .ZN(n108) );
  AOI22_X1 U148 ( .A1(n108), .A2(addr_w_0[1]), .B1(addr_w_0[2]), .B2(n103), 
        .ZN(n113) );
  INV_X1 U150 ( .A(n109), .ZN(n111) );
  OAI22_X1 U151 ( .A1(n113), .A2(n15), .B1(n111), .B2(n110), .ZN(n135) );
  INV_X1 U152 ( .A(n114), .ZN(n120) );
  NAND2_X1 U153 ( .A1(n115), .A2(n6), .ZN(n117) );
  NAND2_X1 U154 ( .A1(n117), .A2(n121), .ZN(n123) );
  INV_X1 U155 ( .A(n123), .ZN(n119) );
  INV_X1 U156 ( .A(n116), .ZN(n150) );
  INV_X1 U157 ( .A(n117), .ZN(n118) );
  NAND3_X1 U158 ( .A1(n11), .A2(n151), .A3(n118), .ZN(n159) );
  NAND3_X1 U159 ( .A1(n60), .A2(n107), .A3(n59), .ZN(n106) );
endmodule


module layer1_8_4_8_16 ( clk, reset, s_valid, m_ready, data_in, m_valid, 
        s_ready, data_out );
  input [15:0] data_in;
  output [15:0] data_out;
  input clk, reset, s_valid, m_ready;
  output m_valid, s_ready;
  wire   wr_en_x, \addr_b_0[0] , \addr_b_1[0] , \addr_b_2[0] , \addr_b_3[0] ,
         \addr_b_4[0] , \addr_b_5[0] , \addr_b_6[0] , \addr_b_7[0] , clear_acc,
         wr_en_y, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131;
  wire   [15:0] data_out_x;
  wire   [2:0] addr_x;
  wire   [2:0] addr_w_0;
  wire   [15:0] data_out_w_0;
  wire   [15:0] data_out_b_0;
  wire   [2:0] addr_w_1;
  wire   [15:0] data_out_w_1;
  wire   [15:0] data_out_b_1;
  wire   [2:0] addr_w_2;
  wire   [15:0] data_out_w_2;
  wire   [15:0] data_out_b_2;
  wire   [2:0] addr_w_3;
  wire   [15:0] data_out_w_3;
  wire   [15:0] data_out_b_3;
  wire   [2:0] addr_w_4;
  wire   [15:0] data_out_w_4;
  wire   [15:0] data_out_b_4;
  wire   [2:0] addr_w_5;
  wire   [15:0] data_out_w_5;
  wire   [15:0] data_out_b_5;
  wire   [2:0] addr_w_6;
  wire   [15:0] data_out_w_6;
  wire   [15:0] data_out_b_6;
  wire   [2:0] addr_w_7;
  wire   [15:0] data_out_w_7;
  wire   [15:0] data_out_b_7;
  wire   [15:0] data_out_0;
  wire   [3:0] sel;
  wire   [15:0] data_out_1;
  wire   [15:0] data_out_2;
  wire   [15:0] data_out_3;
  wire   [15:0] data_out_4;
  wire   [15:0] data_out_5;
  wire   [15:0] data_out_6;
  wire   [15:0] data_out_7;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22;

  memory_WIDTH16_SIZE4_LOGSIZE3 mem_x ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_x), .addr(addr_x), .wr_en(wr_en_x) );
  layer1_8_4_8_16_W_rom_0 mem_w_0 ( .clk(clk), .addr(addr_w_0), .z({
        data_out_w_0[15:2], SYNOPSYS_UNCONNECTED__0, data_out_w_0[0]}) );
  layer1_8_4_8_16_B_rom_0 mem_b_0 ( .clk(clk), .addr(\addr_b_0[0] ) );
  layer1_8_4_8_16_W_rom_1 mem_w_1 ( .clk(clk), .addr(addr_w_1), .z({
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, data_out_w_1[6:0]}) );
  layer1_8_4_8_16_B_rom_1 mem_b_1 ( .clk(clk), .addr(\addr_b_1[0] ) );
  layer1_8_4_8_16_W_rom_2 mem_w_2 ( .clk(clk), .addr(addr_w_2), .z(
        data_out_w_2) );
  layer1_8_4_8_16_B_rom_2 mem_b_2 ( .clk(clk), .addr(\addr_b_2[0] ) );
  layer1_8_4_8_16_W_rom_3 mem_w_3 ( .clk(clk), .addr(addr_w_3), .z({
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, data_out_w_3[6:2], SYNOPSYS_UNCONNECTED__19, 
        data_out_w_3[0]}) );
  layer1_8_4_8_16_B_rom_3 mem_b_3 ( .clk(clk), .addr(\addr_b_3[0] ) );
  layer1_8_4_8_16_W_rom_4 mem_w_4 ( .clk(clk), .addr(addr_w_4), .z(
        data_out_w_4) );
  layer1_8_4_8_16_B_rom_4 mem_b_4 ( .clk(clk), .addr(\addr_b_4[0] ) );
  layer1_8_4_8_16_W_rom_5 mem_w_5 ( .clk(clk), .addr(addr_w_5), .z({
        data_out_w_5[15:4], SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        data_out_w_5[1:0]}) );
  layer1_8_4_8_16_B_rom_5 mem_b_5 ( .clk(clk), .addr(\addr_b_5[0] ) );
  layer1_8_4_8_16_W_rom_6 mem_w_6 ( .clk(clk), .addr(addr_w_6), .z(
        data_out_w_6) );
  layer1_8_4_8_16_B_rom_6 mem_b_6 ( .clk(clk), .addr(\addr_b_6[0] ) );
  layer1_8_4_8_16_W_rom_7 mem_w_7 ( .clk(clk), .addr(addr_w_7), .z({
        data_out_w_7[15:3], SYNOPSYS_UNCONNECTED__22, data_out_w_7[1:0]}) );
  layer1_8_4_8_16_B_rom_7 mem_b_7 ( .clk(clk), .addr(\addr_b_7[0] ) );
  layer1_8_4_8_16_datapath_M8_N4_T16_P8_0 d_0 ( .clk(clk), .clear_acc(
        clear_acc), .data_out_x({data_out_x[15:14], n3, n5, data_out_x[11:9], 
        n9, data_out_x[7], n108, n113, n7, data_out_x[3], n17, data_out_x[1], 
        n110}), .data_out(data_out_0), .data_out_w({data_out_w_0[15:2], 1'b0, 
        data_out_w_0[0]}), .data_out_b({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1}), 
        .wr_en_y(wr_en_y), .m_valid(m_valid), .m_ready(m_ready), .sel(sel) );
  layer1_8_4_8_16_datapath_M8_N4_T16_P8_7 d_1 ( .clk(clk), .clear_acc(
        clear_acc), .data_out_x({data_out_x[15:14], n4, n5, n1, 
        data_out_x[10:9], n12, data_out_x[7], n19, data_out_x[5], n7, n112, 
        n16, n111, n15}), .data_out(data_out_1), .data_out_w({1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, data_out_w_1[6:0]}), .data_out_b({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b0}), .wr_en_y(wr_en_y), .m_valid(m_valid), 
        .m_ready(m_ready), .sel(sel) );
  layer1_8_4_8_16_datapath_M8_N4_T16_P8_6 d_2 ( .clk(clk), .clear_acc(
        clear_acc), .data_out_x({data_out_x[15:14], n4, n5, data_out_x[11:9], 
        n12, data_out_x[7], n14, data_out_x[5], n7, n11, n16, n111, n15}), 
        .data_out(data_out_2), .data_out_w(data_out_w_2), .data_out_b({1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 
        1'b0, 1'b1, 1'b0}), .wr_en_y(wr_en_y), .m_valid(m_valid), .m_ready(
        m_ready), .sel(sel) );
  layer1_8_4_8_16_datapath_M8_N4_T16_P8_5 d_3 ( .clk(clk), .clear_acc(
        clear_acc), .data_out_x({data_out_x[15:14], n4, n5, data_out_x[11:9], 
        n12, data_out_x[7], n19, data_out_x[5], n8, data_out_x[3], n10, 
        data_out_x[1], n110}), .data_out(data_out_3), .data_out_w({1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, data_out_w_3[6:2], 1'b0, 
        data_out_w_3[0]}), .data_out_b({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0}), 
        .wr_en_y(wr_en_y), .m_valid(m_valid), .m_ready(m_ready), .sel(sel) );
  layer1_8_4_8_16_datapath_M8_N4_T16_P8_4 d_4 ( .clk(clk), .clear_acc(
        clear_acc), .data_out_x({data_out_x[15:14], n4, n5, data_out_x[11:9], 
        n9, data_out_x[7], n108, data_out_x[5], n8, n112, n16, data_out_x[1], 
        n15}), .data_out(data_out_4), .data_out_w(data_out_w_4), .data_out_b({
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 
        1'b1, 1'b0, 1'b0, 1'b0}), .wr_en_y(wr_en_y), .m_valid(m_valid), 
        .m_ready(m_ready), .sel(sel) );
  layer1_8_4_8_16_datapath_M8_N4_T16_P8_3 d_5 ( .clk(clk), .clear_acc(
        clear_acc), .data_out_x({data_out_x[15:14], n3, n5, data_out_x[11:9], 
        n9, data_out_x[7], n13, n113, n6, data_out_x[3], n10, data_out_x[1], 
        n15}), .data_out(data_out_5), .data_out_w({data_out_w_5[15:4], 1'b0, 
        1'b1, data_out_w_5[1:0]}), .data_out_b({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1}), 
        .wr_en_y(wr_en_y), .m_valid(m_valid), .m_ready(m_ready), .sel(sel) );
  layer1_8_4_8_16_datapath_M8_N4_T16_P8_2 d_6 ( .clk(clk), .clear_acc(
        clear_acc), .data_out_x({data_out_x[15:14], n4, data_out_x[12:9], n12, 
        data_out_x[7], n14, data_out_x[5], n6, data_out_x[3], n17, 
        data_out_x[1], n110}), .data_out(data_out_6), .data_out_w(data_out_w_6), .data_out_b({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 
        1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1}), .wr_en_y(wr_en_y), .m_valid(
        m_valid), .m_ready(m_ready), .sel(sel) );
  layer1_8_4_8_16_datapath_M8_N4_T16_P8_1 d_7 ( .clk(clk), .clear_acc(
        clear_acc), .data_out_x({data_out_x[15:14], n4, n5, n2, 
        data_out_x[10:9], n9, data_out_x[7], n19, n113, n8, n11, n16, n18, 
        n110}), .data_out(data_out_7), .data_out_w({data_out_w_7[15:3], 1'b1, 
        data_out_w_7[1:0]}), .data_out_b({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1}), 
        .wr_en_y(wr_en_y), .m_valid(m_valid), .m_ready(m_ready), .sel(sel) );
  layer1_8_4_8_16_ctrlpath_M8_N4_T16_P8 c ( .clk(clk), .reset(reset), 
        .s_valid(s_valid), .s_ready(s_ready), .m_valid(m_valid), .m_ready(
        m_ready), .clear_acc(clear_acc), .wr_en_x(wr_en_x), .wr_en_y(wr_en_y), 
        .sel(sel), .addr_x(addr_x), .addr_w_0(addr_w_0), .addr_b_0(
        \addr_b_0[0] ), .addr_w_1(addr_w_1), .addr_b_1(\addr_b_1[0] ), 
        .addr_w_2(addr_w_2), .addr_b_2(\addr_b_2[0] ), .addr_w_3(addr_w_3), 
        .addr_b_3(\addr_b_3[0] ), .addr_w_4(addr_w_4), .addr_b_4(\addr_b_4[0] ), .addr_w_5(addr_w_5), .addr_b_5(\addr_b_5[0] ), .addr_w_6(addr_w_6), 
        .addr_b_6(\addr_b_6[0] ), .addr_w_7(addr_w_7), .addr_b_7(\addr_b_7[0] ) );
  CLKBUF_X1 U1 ( .A(data_out_x[11]), .Z(n1) );
  BUF_X2 U2 ( .A(data_out_x[3]), .Z(n112) );
  BUF_X2 U3 ( .A(data_out_x[6]), .Z(n13) );
  BUF_X4 U4 ( .A(data_out_x[0]), .Z(n15) );
  BUF_X2 U5 ( .A(data_out_x[8]), .Z(n12) );
  CLKBUF_X3 U6 ( .A(data_out_x[8]), .Z(n9) );
  BUF_X1 U7 ( .A(data_out_x[5]), .Z(n113) );
  BUF_X2 U8 ( .A(data_out_x[6]), .Z(n19) );
  BUF_X1 U9 ( .A(data_out_x[1]), .Z(n18) );
  BUF_X2 U10 ( .A(data_out_x[4]), .Z(n6) );
  CLKBUF_X1 U11 ( .A(data_out_x[11]), .Z(n2) );
  CLKBUF_X1 U12 ( .A(data_out_x[13]), .Z(n3) );
  BUF_X2 U13 ( .A(data_out_x[13]), .Z(n4) );
  CLKBUF_X3 U14 ( .A(data_out_x[2]), .Z(n16) );
  BUF_X4 U15 ( .A(data_out_x[12]), .Z(n5) );
  CLKBUF_X3 U16 ( .A(data_out_x[4]), .Z(n7) );
  CLKBUF_X3 U17 ( .A(data_out_x[4]), .Z(n8) );
  BUF_X1 U18 ( .A(data_out_x[3]), .Z(n11) );
  BUF_X2 U19 ( .A(data_out_x[2]), .Z(n17) );
  BUF_X2 U20 ( .A(data_out_x[2]), .Z(n10) );
  BUF_X1 U21 ( .A(data_out_x[6]), .Z(n14) );
  BUF_X2 U22 ( .A(data_out_x[6]), .Z(n108) );
  BUF_X1 U23 ( .A(data_out_x[1]), .Z(n111) );
  NOR3_X4 U24 ( .A1(sel[1]), .A2(sel[2]), .A3(sel[0]), .ZN(n32) );
  NOR3_X4 U25 ( .A1(sel[1]), .A2(sel[2]), .A3(n130), .ZN(n31) );
  INV_X1 U26 ( .A(sel[3]), .ZN(n109) );
  AND3_X1 U27 ( .A1(sel[0]), .A2(n131), .A3(sel[2]), .ZN(n27) );
  AND3_X1 U28 ( .A1(sel[1]), .A2(sel[0]), .A3(sel[2]), .ZN(n25) );
  AND3_X1 U29 ( .A1(sel[1]), .A2(n130), .A3(sel[2]), .ZN(n26) );
  AND3_X1 U30 ( .A1(n130), .A2(n131), .A3(sel[2]), .ZN(n28) );
  AOI22_X1 U31 ( .A1(data_out_1[0]), .A2(n31), .B1(data_out_0[0]), .B2(n32), 
        .ZN(n104) );
  AOI22_X1 U32 ( .A1(data_out_1[1]), .A2(n31), .B1(data_out_0[1]), .B2(n32), 
        .ZN(n69) );
  AOI22_X1 U33 ( .A1(data_out_1[2]), .A2(n31), .B1(data_out_0[2]), .B2(n32), 
        .ZN(n64) );
  AOI22_X1 U34 ( .A1(data_out_1[3]), .A2(n31), .B1(data_out_0[3]), .B2(n32), 
        .ZN(n59) );
  AOI22_X1 U35 ( .A1(data_out_1[4]), .A2(n31), .B1(data_out_0[4]), .B2(n32), 
        .ZN(n54) );
  AOI22_X1 U36 ( .A1(data_out_1[5]), .A2(n31), .B1(data_out_0[5]), .B2(n32), 
        .ZN(n49) );
  AOI22_X1 U37 ( .A1(data_out_1[6]), .A2(n31), .B1(data_out_0[6]), .B2(n32), 
        .ZN(n44) );
  AOI22_X1 U38 ( .A1(data_out_1[7]), .A2(n31), .B1(data_out_0[7]), .B2(n32), 
        .ZN(n39) );
  AOI22_X1 U39 ( .A1(data_out_1[8]), .A2(n31), .B1(data_out_0[8]), .B2(n32), 
        .ZN(n34) );
  AOI22_X1 U40 ( .A1(data_out_1[9]), .A2(n31), .B1(data_out_0[9]), .B2(n32), 
        .ZN(n21) );
  AOI22_X1 U41 ( .A1(data_out_1[10]), .A2(n31), .B1(data_out_0[10]), .B2(n32), 
        .ZN(n99) );
  AOI22_X1 U42 ( .A1(data_out_1[11]), .A2(n31), .B1(data_out_0[11]), .B2(n32), 
        .ZN(n94) );
  AOI22_X1 U43 ( .A1(data_out_1[12]), .A2(n31), .B1(data_out_0[12]), .B2(n32), 
        .ZN(n89) );
  AOI22_X1 U44 ( .A1(data_out_1[13]), .A2(n31), .B1(data_out_0[13]), .B2(n32), 
        .ZN(n84) );
  AOI22_X1 U45 ( .A1(data_out_1[14]), .A2(n31), .B1(data_out_0[14]), .B2(n32), 
        .ZN(n79) );
  AOI22_X1 U46 ( .A1(data_out_1[15]), .A2(n31), .B1(data_out_0[15]), .B2(n32), 
        .ZN(n74) );
  OAI22_X1 U47 ( .A1(n109), .A2(n129), .B1(sel[3]), .B2(n103), .ZN(data_out[0]) );
  INV_X1 U48 ( .A(data_out_7[0]), .ZN(n129) );
  AND4_X1 U49 ( .A1(n104), .A2(n105), .A3(n106), .A4(n107), .ZN(n103) );
  OAI22_X1 U50 ( .A1(n109), .A2(n128), .B1(sel[3]), .B2(n68), .ZN(data_out[1])
         );
  INV_X1 U51 ( .A(data_out_7[1]), .ZN(n128) );
  AND4_X1 U52 ( .A1(n69), .A2(n70), .A3(n71), .A4(n72), .ZN(n68) );
  OAI22_X1 U53 ( .A1(n109), .A2(n127), .B1(sel[3]), .B2(n63), .ZN(data_out[2])
         );
  INV_X1 U54 ( .A(data_out_7[2]), .ZN(n127) );
  AND4_X1 U55 ( .A1(n64), .A2(n65), .A3(n66), .A4(n67), .ZN(n63) );
  OAI22_X1 U56 ( .A1(n109), .A2(n126), .B1(sel[3]), .B2(n58), .ZN(data_out[3])
         );
  INV_X1 U57 ( .A(data_out_7[3]), .ZN(n126) );
  AND4_X1 U58 ( .A1(n59), .A2(n60), .A3(n61), .A4(n62), .ZN(n58) );
  OAI22_X1 U59 ( .A1(n109), .A2(n125), .B1(sel[3]), .B2(n53), .ZN(data_out[4])
         );
  INV_X1 U60 ( .A(data_out_7[4]), .ZN(n125) );
  AND4_X1 U61 ( .A1(n54), .A2(n55), .A3(n56), .A4(n57), .ZN(n53) );
  OAI22_X1 U62 ( .A1(n109), .A2(n124), .B1(sel[3]), .B2(n48), .ZN(data_out[5])
         );
  INV_X1 U63 ( .A(data_out_7[5]), .ZN(n124) );
  AND4_X1 U64 ( .A1(n49), .A2(n50), .A3(n51), .A4(n52), .ZN(n48) );
  OAI22_X1 U65 ( .A1(n109), .A2(n123), .B1(sel[3]), .B2(n43), .ZN(data_out[6])
         );
  INV_X1 U66 ( .A(data_out_7[6]), .ZN(n123) );
  AND4_X1 U67 ( .A1(n44), .A2(n45), .A3(n46), .A4(n47), .ZN(n43) );
  OAI22_X1 U68 ( .A1(n109), .A2(n122), .B1(sel[3]), .B2(n38), .ZN(data_out[7])
         );
  INV_X1 U69 ( .A(data_out_7[7]), .ZN(n122) );
  AND4_X1 U70 ( .A1(n39), .A2(n40), .A3(n41), .A4(n42), .ZN(n38) );
  OAI22_X1 U71 ( .A1(n109), .A2(n121), .B1(sel[3]), .B2(n33), .ZN(data_out[8])
         );
  INV_X1 U72 ( .A(data_out_7[8]), .ZN(n121) );
  AND4_X1 U73 ( .A1(n34), .A2(n35), .A3(n36), .A4(n37), .ZN(n33) );
  OAI22_X1 U74 ( .A1(n120), .A2(n109), .B1(sel[3]), .B2(n20), .ZN(data_out[9])
         );
  INV_X1 U75 ( .A(data_out_7[9]), .ZN(n120) );
  AND4_X1 U76 ( .A1(n21), .A2(n22), .A3(n23), .A4(n24), .ZN(n20) );
  OAI22_X1 U77 ( .A1(n109), .A2(n119), .B1(sel[3]), .B2(n98), .ZN(data_out[10]) );
  INV_X1 U78 ( .A(data_out_7[10]), .ZN(n119) );
  AND4_X1 U79 ( .A1(n99), .A2(n100), .A3(n101), .A4(n102), .ZN(n98) );
  OAI22_X1 U80 ( .A1(n109), .A2(n118), .B1(sel[3]), .B2(n93), .ZN(data_out[11]) );
  INV_X1 U81 ( .A(data_out_7[11]), .ZN(n118) );
  AND4_X1 U82 ( .A1(n94), .A2(n95), .A3(n96), .A4(n97), .ZN(n93) );
  OAI22_X1 U83 ( .A1(n109), .A2(n117), .B1(sel[3]), .B2(n88), .ZN(data_out[12]) );
  INV_X1 U84 ( .A(data_out_7[12]), .ZN(n117) );
  AND4_X1 U85 ( .A1(n89), .A2(n90), .A3(n91), .A4(n92), .ZN(n88) );
  OAI22_X1 U86 ( .A1(n109), .A2(n116), .B1(sel[3]), .B2(n83), .ZN(data_out[13]) );
  INV_X1 U87 ( .A(data_out_7[13]), .ZN(n116) );
  AND4_X1 U88 ( .A1(n84), .A2(n85), .A3(n86), .A4(n87), .ZN(n83) );
  OAI22_X1 U89 ( .A1(n109), .A2(n115), .B1(sel[3]), .B2(n78), .ZN(data_out[14]) );
  INV_X1 U90 ( .A(data_out_7[14]), .ZN(n115) );
  AND4_X1 U91 ( .A1(n79), .A2(n80), .A3(n81), .A4(n82), .ZN(n78) );
  OAI22_X1 U92 ( .A1(n109), .A2(n114), .B1(sel[3]), .B2(n73), .ZN(data_out[15]) );
  INV_X1 U93 ( .A(data_out_7[15]), .ZN(n114) );
  AND4_X1 U94 ( .A1(n74), .A2(n75), .A3(n76), .A4(n77), .ZN(n73) );
  AOI22_X1 U95 ( .A1(data_out_3[0]), .A2(n29), .B1(data_out_2[0]), .B2(n30), 
        .ZN(n105) );
  AOI22_X1 U96 ( .A1(data_out_3[1]), .A2(n29), .B1(data_out_2[1]), .B2(n30), 
        .ZN(n70) );
  AOI22_X1 U97 ( .A1(data_out_3[2]), .A2(n29), .B1(data_out_2[2]), .B2(n30), 
        .ZN(n65) );
  AOI22_X1 U98 ( .A1(data_out_3[3]), .A2(n29), .B1(data_out_2[3]), .B2(n30), 
        .ZN(n60) );
  AOI22_X1 U99 ( .A1(data_out_3[4]), .A2(n29), .B1(data_out_2[4]), .B2(n30), 
        .ZN(n55) );
  AOI22_X1 U100 ( .A1(data_out_3[5]), .A2(n29), .B1(data_out_2[5]), .B2(n30), 
        .ZN(n50) );
  AOI22_X1 U101 ( .A1(data_out_3[6]), .A2(n29), .B1(data_out_2[6]), .B2(n30), 
        .ZN(n45) );
  AOI22_X1 U102 ( .A1(data_out_3[7]), .A2(n29), .B1(data_out_2[7]), .B2(n30), 
        .ZN(n40) );
  AOI22_X1 U103 ( .A1(data_out_3[8]), .A2(n29), .B1(data_out_2[8]), .B2(n30), 
        .ZN(n35) );
  AOI22_X1 U104 ( .A1(data_out_3[9]), .A2(n29), .B1(data_out_2[9]), .B2(n30), 
        .ZN(n22) );
  AOI22_X1 U105 ( .A1(data_out_3[10]), .A2(n29), .B1(data_out_2[10]), .B2(n30), 
        .ZN(n100) );
  AOI22_X1 U106 ( .A1(data_out_3[11]), .A2(n29), .B1(data_out_2[11]), .B2(n30), 
        .ZN(n95) );
  AOI22_X1 U107 ( .A1(data_out_3[12]), .A2(n29), .B1(data_out_2[12]), .B2(n30), 
        .ZN(n90) );
  AOI22_X1 U108 ( .A1(data_out_3[13]), .A2(n29), .B1(data_out_2[13]), .B2(n30), 
        .ZN(n85) );
  AOI22_X1 U109 ( .A1(data_out_3[14]), .A2(n29), .B1(data_out_2[14]), .B2(n30), 
        .ZN(n80) );
  AOI22_X1 U110 ( .A1(data_out_3[15]), .A2(n29), .B1(data_out_2[15]), .B2(n30), 
        .ZN(n75) );
  AOI22_X1 U111 ( .A1(data_out_7[0]), .A2(n25), .B1(data_out_6[0]), .B2(n26), 
        .ZN(n107) );
  AOI22_X1 U112 ( .A1(data_out_7[1]), .A2(n25), .B1(data_out_6[1]), .B2(n26), 
        .ZN(n72) );
  AOI22_X1 U113 ( .A1(data_out_7[2]), .A2(n25), .B1(data_out_6[2]), .B2(n26), 
        .ZN(n67) );
  AOI22_X1 U114 ( .A1(data_out_7[3]), .A2(n25), .B1(data_out_6[3]), .B2(n26), 
        .ZN(n62) );
  AOI22_X1 U115 ( .A1(data_out_7[4]), .A2(n25), .B1(data_out_6[4]), .B2(n26), 
        .ZN(n57) );
  AOI22_X1 U116 ( .A1(data_out_7[5]), .A2(n25), .B1(data_out_6[5]), .B2(n26), 
        .ZN(n52) );
  AOI22_X1 U117 ( .A1(data_out_7[6]), .A2(n25), .B1(data_out_6[6]), .B2(n26), 
        .ZN(n47) );
  AOI22_X1 U118 ( .A1(data_out_7[7]), .A2(n25), .B1(data_out_6[7]), .B2(n26), 
        .ZN(n42) );
  AOI22_X1 U119 ( .A1(data_out_7[8]), .A2(n25), .B1(data_out_6[8]), .B2(n26), 
        .ZN(n37) );
  AOI22_X1 U120 ( .A1(data_out_7[9]), .A2(n25), .B1(data_out_6[9]), .B2(n26), 
        .ZN(n24) );
  AOI22_X1 U121 ( .A1(data_out_7[10]), .A2(n25), .B1(data_out_6[10]), .B2(n26), 
        .ZN(n102) );
  AOI22_X1 U122 ( .A1(data_out_7[11]), .A2(n25), .B1(data_out_6[11]), .B2(n26), 
        .ZN(n97) );
  AOI22_X1 U123 ( .A1(data_out_7[12]), .A2(n25), .B1(data_out_6[12]), .B2(n26), 
        .ZN(n92) );
  AOI22_X1 U124 ( .A1(data_out_7[13]), .A2(n25), .B1(data_out_6[13]), .B2(n26), 
        .ZN(n87) );
  AOI22_X1 U125 ( .A1(data_out_7[14]), .A2(n25), .B1(data_out_6[14]), .B2(n26), 
        .ZN(n82) );
  AOI22_X1 U126 ( .A1(data_out_7[15]), .A2(n25), .B1(data_out_6[15]), .B2(n26), 
        .ZN(n77) );
  AOI22_X1 U127 ( .A1(data_out_5[0]), .A2(n27), .B1(data_out_4[0]), .B2(n28), 
        .ZN(n106) );
  AOI22_X1 U128 ( .A1(data_out_5[1]), .A2(n27), .B1(data_out_4[1]), .B2(n28), 
        .ZN(n71) );
  AOI22_X1 U129 ( .A1(data_out_5[2]), .A2(n27), .B1(data_out_4[2]), .B2(n28), 
        .ZN(n66) );
  AOI22_X1 U130 ( .A1(data_out_5[3]), .A2(n27), .B1(data_out_4[3]), .B2(n28), 
        .ZN(n61) );
  AOI22_X1 U131 ( .A1(data_out_5[4]), .A2(n27), .B1(data_out_4[4]), .B2(n28), 
        .ZN(n56) );
  AOI22_X1 U132 ( .A1(data_out_5[5]), .A2(n27), .B1(data_out_4[5]), .B2(n28), 
        .ZN(n51) );
  AOI22_X1 U133 ( .A1(data_out_5[6]), .A2(n27), .B1(data_out_4[6]), .B2(n28), 
        .ZN(n46) );
  AOI22_X1 U134 ( .A1(data_out_5[7]), .A2(n27), .B1(data_out_4[7]), .B2(n28), 
        .ZN(n41) );
  AOI22_X1 U135 ( .A1(data_out_5[8]), .A2(n27), .B1(data_out_4[8]), .B2(n28), 
        .ZN(n36) );
  AOI22_X1 U136 ( .A1(data_out_5[9]), .A2(n27), .B1(data_out_4[9]), .B2(n28), 
        .ZN(n23) );
  AOI22_X1 U137 ( .A1(data_out_5[10]), .A2(n27), .B1(data_out_4[10]), .B2(n28), 
        .ZN(n101) );
  AOI22_X1 U138 ( .A1(data_out_5[11]), .A2(n27), .B1(data_out_4[11]), .B2(n28), 
        .ZN(n96) );
  AOI22_X1 U139 ( .A1(data_out_5[12]), .A2(n27), .B1(data_out_4[12]), .B2(n28), 
        .ZN(n91) );
  AOI22_X1 U140 ( .A1(data_out_5[13]), .A2(n27), .B1(data_out_4[13]), .B2(n28), 
        .ZN(n86) );
  AOI22_X1 U141 ( .A1(data_out_5[14]), .A2(n27), .B1(data_out_4[14]), .B2(n28), 
        .ZN(n81) );
  AOI22_X1 U142 ( .A1(data_out_5[15]), .A2(n27), .B1(data_out_4[15]), .B2(n28), 
        .ZN(n76) );
  INV_X1 U143 ( .A(sel[0]), .ZN(n130) );
  INV_X1 U144 ( .A(sel[1]), .ZN(n131) );
  BUF_X4 U145 ( .A(data_out_x[0]), .Z(n110) );
  NOR3_X4 U146 ( .A1(n130), .A2(sel[2]), .A3(n131), .ZN(n29) );
  NOR3_X4 U147 ( .A1(sel[0]), .A2(sel[2]), .A3(n131), .ZN(n30) );
endmodule


module memory_WIDTH16_SIZE8_LOGSIZE4 ( clk, data_in, data_out, addr, wr_en );
  input [15:0] data_in;
  output [15:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][15] , \mem[7][14] , \mem[7][13] , \mem[7][12] ,
         \mem[7][11] , \mem[7][10] , \mem[7][9] , \mem[7][8] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][15] , \mem[6][14] , \mem[6][13] ,
         \mem[6][12] , \mem[6][11] , \mem[6][10] , \mem[6][9] , \mem[6][8] ,
         \mem[6][7] , \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] ,
         \mem[6][2] , \mem[6][1] , \mem[6][0] , \mem[5][15] , \mem[5][14] ,
         \mem[5][13] , \mem[5][12] , \mem[5][11] , \mem[5][10] , \mem[5][9] ,
         \mem[5][8] , \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] ,
         \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][15] ,
         \mem[4][14] , \mem[4][13] , \mem[4][12] , \mem[4][11] , \mem[4][10] ,
         \mem[4][9] , \mem[4][8] , \mem[4][7] , \mem[4][6] , \mem[4][5] ,
         \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] , \mem[4][0] ,
         \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] ,
         \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][15] , \mem[1][14] , \mem[1][13] ,
         \mem[1][12] , \mem[1][11] , \mem[1][10] , \mem[1][9] , \mem[1][8] ,
         \mem[1][7] , \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] ,
         \mem[1][2] , \mem[1][1] , \mem[1][0] , \mem[0][15] , \mem[0][14] ,
         \mem[0][13] , \mem[0][12] , \mem[0][11] , \mem[0][10] , \mem[0][9] ,
         \mem[0][8] , \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] ,
         \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N28, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n1, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[15]  ( .D(N13), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \data_out_reg[14]  ( .D(N14), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[12]  ( .D(N16), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[10]  ( .D(N18), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[8]  ( .D(N20), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[7]  ( .D(N21), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N22), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N23), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N24), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[3]  ( .D(N25), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[2]  ( .D(N26), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N28), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[7][15]  ( .D(n287), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n286), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n285), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n284), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n283), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n282), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n281), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n280), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n279), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n278), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n277), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n276), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n275), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n274), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n273), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n272), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n271), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n270), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n269), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n268), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n267), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n266), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n265), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n264), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n263), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n262), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n261), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n260), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n259), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n258), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n257), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n256), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n255), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n254), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n253), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n252), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n251), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n250), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n249), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n248), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n247), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n246), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n245), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n244), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n243), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n242), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n241), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n240), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n239), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n238), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n237), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n236), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n235), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n234), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n233), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n232), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n231), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n230), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n229), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n228), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n227), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n226), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n225), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n224), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n223), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n222), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n221), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n220), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n219), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n218), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n217), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n216), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n215), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n214), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n213), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n212), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n211), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n210), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n209), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n208), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n207), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n206), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n205), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n204), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n203), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n202), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n201), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n200), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n199), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n198), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n197), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n196), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n195), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n194), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n193), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n192), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n191), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n190), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n189), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n188), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n187), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n186), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n185), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n184), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n183), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n182), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n181), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n180), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n179), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n178), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n177), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n176), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n167), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n166), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n165), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n164), .CK(clk), .Q(\mem[0][4] ) );
  NAND3_X1 U282 ( .A1(n398), .A2(n399), .A3(n38), .ZN(n21) );
  NAND3_X1 U283 ( .A1(n38), .A2(n399), .A3(N10), .ZN(n39) );
  NAND3_X1 U284 ( .A1(n38), .A2(n398), .A3(N11), .ZN(n56) );
  NAND3_X1 U285 ( .A1(N10), .A2(n38), .A3(N11), .ZN(n73) );
  NAND3_X1 U286 ( .A1(n398), .A2(n399), .A3(n108), .ZN(n91) );
  NAND3_X1 U287 ( .A1(N10), .A2(n399), .A3(n108), .ZN(n109) );
  NAND3_X1 U288 ( .A1(N11), .A2(n398), .A3(n108), .ZN(n126) );
  NAND3_X1 U289 ( .A1(N11), .A2(N10), .A3(n108), .ZN(n143) );
  DFF_X1 \data_out_reg[9]  ( .D(N19), .CK(clk), .QN(n1) );
  DFF_X1 \mem_reg[0][14]  ( .D(n174), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n173), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n172), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n171), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n170), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n169), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n168), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n175), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n163), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n162), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n161), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n160), .CK(clk), .Q(\mem[0][0] ) );
  SDFF_X1 \data_out_reg[1]  ( .D(n14), .SI(n11), .SE(N12), .CK(clk), .Q(
        data_out[1]) );
  DFF_X2 \data_out_reg[11]  ( .D(N17), .CK(clk), .Q(data_out[11]) );
  DFF_X2 \data_out_reg[13]  ( .D(N15), .CK(clk), .Q(data_out[13]) );
  INV_X2 U3 ( .A(n1), .ZN(data_out[9]) );
  BUF_X1 U4 ( .A(n21), .Z(n395) );
  BUF_X1 U5 ( .A(n56), .Z(n390) );
  BUF_X1 U6 ( .A(n39), .Z(n393) );
  BUF_X1 U7 ( .A(n73), .Z(n387) );
  BUF_X1 U8 ( .A(n91), .Z(n384) );
  BUF_X1 U9 ( .A(n126), .Z(n378) );
  BUF_X1 U10 ( .A(n109), .Z(n381) );
  BUF_X1 U11 ( .A(n143), .Z(n375) );
  BUF_X1 U12 ( .A(N10), .Z(n372) );
  BUF_X1 U13 ( .A(N10), .Z(n373) );
  BUF_X1 U14 ( .A(n21), .Z(n396) );
  BUF_X1 U15 ( .A(n39), .Z(n392) );
  BUF_X1 U16 ( .A(n109), .Z(n380) );
  BUF_X1 U17 ( .A(n143), .Z(n374) );
  BUF_X1 U18 ( .A(n126), .Z(n377) );
  BUF_X1 U19 ( .A(n91), .Z(n383) );
  BUF_X1 U20 ( .A(n73), .Z(n386) );
  BUF_X1 U21 ( .A(n56), .Z(n389) );
  CLKBUF_X1 U22 ( .A(n39), .Z(n394) );
  CLKBUF_X1 U23 ( .A(n109), .Z(n382) );
  CLKBUF_X1 U24 ( .A(n143), .Z(n376) );
  CLKBUF_X1 U25 ( .A(n126), .Z(n379) );
  CLKBUF_X1 U26 ( .A(n91), .Z(n385) );
  CLKBUF_X1 U27 ( .A(n73), .Z(n388) );
  CLKBUF_X1 U28 ( .A(n56), .Z(n391) );
  BUF_X1 U29 ( .A(N10), .Z(n369) );
  BUF_X1 U30 ( .A(N10), .Z(n370) );
  BUF_X1 U31 ( .A(N10), .Z(n371) );
  BUF_X1 U32 ( .A(N11), .Z(n367) );
  BUF_X1 U33 ( .A(N11), .Z(n368) );
  CLKBUF_X1 U34 ( .A(n21), .Z(n397) );
  BUF_X1 U35 ( .A(N11), .Z(n366) );
  INV_X1 U36 ( .A(data_in[0]), .ZN(n415) );
  INV_X1 U37 ( .A(data_in[1]), .ZN(n414) );
  INV_X1 U38 ( .A(data_in[2]), .ZN(n413) );
  INV_X1 U39 ( .A(data_in[3]), .ZN(n412) );
  INV_X1 U40 ( .A(data_in[4]), .ZN(n411) );
  INV_X1 U41 ( .A(data_in[5]), .ZN(n410) );
  INV_X1 U42 ( .A(data_in[6]), .ZN(n409) );
  INV_X1 U43 ( .A(data_in[7]), .ZN(n408) );
  INV_X1 U44 ( .A(data_in[8]), .ZN(n407) );
  INV_X1 U45 ( .A(data_in[9]), .ZN(n406) );
  INV_X1 U46 ( .A(data_in[10]), .ZN(n405) );
  INV_X1 U47 ( .A(data_in[11]), .ZN(n404) );
  INV_X1 U48 ( .A(data_in[12]), .ZN(n403) );
  INV_X1 U49 ( .A(data_in[13]), .ZN(n402) );
  INV_X1 U50 ( .A(data_in[14]), .ZN(n401) );
  INV_X1 U51 ( .A(data_in[15]), .ZN(n400) );
  NOR2_X1 U52 ( .A1(n90), .A2(N12), .ZN(n38) );
  NOR2_X1 U53 ( .A1(n416), .A2(n90), .ZN(n108) );
  INV_X1 U54 ( .A(N12), .ZN(n416) );
  OAI21_X1 U55 ( .B1(n408), .B2(n376), .A(n151), .ZN(n279) );
  NAND2_X1 U56 ( .A1(\mem[7][7] ), .A2(n375), .ZN(n151) );
  OAI21_X1 U57 ( .B1(n407), .B2(n379), .A(n135), .ZN(n264) );
  NAND2_X1 U58 ( .A1(\mem[6][8] ), .A2(n377), .ZN(n135) );
  OAI21_X1 U59 ( .B1(n406), .B2(n379), .A(n136), .ZN(n265) );
  NAND2_X1 U60 ( .A1(\mem[6][9] ), .A2(n377), .ZN(n136) );
  OAI21_X1 U61 ( .B1(n402), .B2(n379), .A(n140), .ZN(n269) );
  NAND2_X1 U62 ( .A1(\mem[6][13] ), .A2(n377), .ZN(n140) );
  OAI21_X1 U63 ( .B1(n401), .B2(n379), .A(n141), .ZN(n270) );
  NAND2_X1 U64 ( .A1(\mem[6][14] ), .A2(n377), .ZN(n141) );
  OAI21_X1 U65 ( .B1(n405), .B2(n379), .A(n137), .ZN(n266) );
  NAND2_X1 U66 ( .A1(\mem[6][10] ), .A2(n377), .ZN(n137) );
  OAI21_X1 U67 ( .B1(n404), .B2(n379), .A(n138), .ZN(n267) );
  NAND2_X1 U68 ( .A1(\mem[6][11] ), .A2(n377), .ZN(n138) );
  OAI21_X1 U69 ( .B1(n403), .B2(n379), .A(n139), .ZN(n268) );
  NAND2_X1 U70 ( .A1(\mem[6][12] ), .A2(n377), .ZN(n139) );
  OAI21_X1 U71 ( .B1(n408), .B2(n391), .A(n64), .ZN(n199) );
  NAND2_X1 U72 ( .A1(\mem[2][7] ), .A2(n390), .ZN(n64) );
  OAI21_X1 U73 ( .B1(n397), .B2(n407), .A(n30), .ZN(n168) );
  NAND2_X1 U74 ( .A1(\mem[0][8] ), .A2(n395), .ZN(n30) );
  OAI21_X1 U75 ( .B1(n397), .B2(n406), .A(n31), .ZN(n169) );
  NAND2_X1 U76 ( .A1(\mem[0][9] ), .A2(n395), .ZN(n31) );
  OAI21_X1 U77 ( .B1(n397), .B2(n402), .A(n35), .ZN(n173) );
  NAND2_X1 U78 ( .A1(\mem[0][13] ), .A2(n395), .ZN(n35) );
  OAI21_X1 U79 ( .B1(n397), .B2(n401), .A(n36), .ZN(n174) );
  NAND2_X1 U80 ( .A1(\mem[0][14] ), .A2(n395), .ZN(n36) );
  OAI21_X1 U81 ( .B1(n397), .B2(n405), .A(n32), .ZN(n170) );
  NAND2_X1 U82 ( .A1(\mem[0][10] ), .A2(n395), .ZN(n32) );
  OAI21_X1 U83 ( .B1(n397), .B2(n404), .A(n33), .ZN(n171) );
  NAND2_X1 U84 ( .A1(\mem[0][11] ), .A2(n395), .ZN(n33) );
  OAI21_X1 U85 ( .B1(n397), .B2(n403), .A(n34), .ZN(n172) );
  NAND2_X1 U86 ( .A1(\mem[0][12] ), .A2(n395), .ZN(n34) );
  INV_X1 U87 ( .A(N11), .ZN(n399) );
  INV_X1 U88 ( .A(N10), .ZN(n398) );
  OAI21_X1 U89 ( .B1(n411), .B2(n375), .A(n148), .ZN(n276) );
  NAND2_X1 U90 ( .A1(\mem[7][4] ), .A2(n375), .ZN(n148) );
  OAI21_X1 U91 ( .B1(n410), .B2(n375), .A(n149), .ZN(n277) );
  NAND2_X1 U92 ( .A1(\mem[7][5] ), .A2(n375), .ZN(n149) );
  OAI21_X1 U93 ( .B1(n409), .B2(n375), .A(n150), .ZN(n278) );
  NAND2_X1 U94 ( .A1(\mem[7][6] ), .A2(n375), .ZN(n150) );
  OAI21_X1 U95 ( .B1(n415), .B2(n378), .A(n127), .ZN(n256) );
  NAND2_X1 U96 ( .A1(\mem[6][0] ), .A2(n377), .ZN(n127) );
  OAI21_X1 U97 ( .B1(n414), .B2(n378), .A(n128), .ZN(n257) );
  NAND2_X1 U98 ( .A1(\mem[6][1] ), .A2(n377), .ZN(n128) );
  OAI21_X1 U99 ( .B1(n413), .B2(n378), .A(n129), .ZN(n258) );
  NAND2_X1 U100 ( .A1(\mem[6][2] ), .A2(n377), .ZN(n129) );
  OAI21_X1 U101 ( .B1(n412), .B2(n378), .A(n130), .ZN(n259) );
  NAND2_X1 U102 ( .A1(\mem[6][3] ), .A2(n377), .ZN(n130) );
  OAI21_X1 U103 ( .B1(n400), .B2(n378), .A(n142), .ZN(n271) );
  NAND2_X1 U104 ( .A1(\mem[6][15] ), .A2(n377), .ZN(n142) );
  OAI21_X1 U105 ( .B1(n411), .B2(n390), .A(n61), .ZN(n196) );
  NAND2_X1 U106 ( .A1(\mem[2][4] ), .A2(n390), .ZN(n61) );
  OAI21_X1 U107 ( .B1(n410), .B2(n390), .A(n62), .ZN(n197) );
  NAND2_X1 U108 ( .A1(\mem[2][5] ), .A2(n390), .ZN(n62) );
  OAI21_X1 U109 ( .B1(n409), .B2(n390), .A(n63), .ZN(n198) );
  NAND2_X1 U110 ( .A1(\mem[2][6] ), .A2(n390), .ZN(n63) );
  OAI21_X1 U111 ( .B1(n396), .B2(n415), .A(n22), .ZN(n160) );
  NAND2_X1 U112 ( .A1(\mem[0][0] ), .A2(n395), .ZN(n22) );
  OAI21_X1 U113 ( .B1(n396), .B2(n414), .A(n23), .ZN(n161) );
  NAND2_X1 U114 ( .A1(\mem[0][1] ), .A2(n395), .ZN(n23) );
  OAI21_X1 U115 ( .B1(n396), .B2(n413), .A(n24), .ZN(n162) );
  NAND2_X1 U116 ( .A1(\mem[0][2] ), .A2(n395), .ZN(n24) );
  OAI21_X1 U117 ( .B1(n396), .B2(n412), .A(n25), .ZN(n163) );
  NAND2_X1 U118 ( .A1(\mem[0][3] ), .A2(n395), .ZN(n25) );
  OAI21_X1 U119 ( .B1(n396), .B2(n400), .A(n37), .ZN(n175) );
  NAND2_X1 U120 ( .A1(\mem[0][15] ), .A2(n395), .ZN(n37) );
  NAND2_X1 U121 ( .A1(wr_en), .A2(n417), .ZN(n90) );
  INV_X1 U122 ( .A(addr[3]), .ZN(n417) );
  OAI21_X1 U123 ( .B1(n408), .B2(n382), .A(n117), .ZN(n247) );
  NAND2_X1 U124 ( .A1(\mem[5][7] ), .A2(n381), .ZN(n117) );
  OAI21_X1 U125 ( .B1(n411), .B2(n381), .A(n114), .ZN(n244) );
  NAND2_X1 U126 ( .A1(\mem[5][4] ), .A2(n381), .ZN(n114) );
  OAI21_X1 U127 ( .B1(n410), .B2(n381), .A(n115), .ZN(n245) );
  NAND2_X1 U128 ( .A1(\mem[5][5] ), .A2(n381), .ZN(n115) );
  OAI21_X1 U129 ( .B1(n409), .B2(n381), .A(n116), .ZN(n246) );
  NAND2_X1 U130 ( .A1(\mem[5][6] ), .A2(n381), .ZN(n116) );
  OAI21_X1 U131 ( .B1(n408), .B2(n388), .A(n81), .ZN(n215) );
  NAND2_X1 U132 ( .A1(\mem[3][7] ), .A2(n387), .ZN(n81) );
  OAI21_X1 U133 ( .B1(n411), .B2(n387), .A(n78), .ZN(n212) );
  NAND2_X1 U134 ( .A1(\mem[3][4] ), .A2(n387), .ZN(n78) );
  OAI21_X1 U135 ( .B1(n410), .B2(n387), .A(n79), .ZN(n213) );
  NAND2_X1 U136 ( .A1(\mem[3][5] ), .A2(n387), .ZN(n79) );
  OAI21_X1 U137 ( .B1(n409), .B2(n387), .A(n80), .ZN(n214) );
  NAND2_X1 U138 ( .A1(\mem[3][6] ), .A2(n387), .ZN(n80) );
  OAI21_X1 U139 ( .B1(n408), .B2(n379), .A(n134), .ZN(n263) );
  NAND2_X1 U140 ( .A1(\mem[6][7] ), .A2(n378), .ZN(n134) );
  OAI21_X1 U141 ( .B1(n411), .B2(n378), .A(n131), .ZN(n260) );
  NAND2_X1 U142 ( .A1(\mem[6][4] ), .A2(n378), .ZN(n131) );
  OAI21_X1 U143 ( .B1(n410), .B2(n378), .A(n132), .ZN(n261) );
  NAND2_X1 U144 ( .A1(\mem[6][5] ), .A2(n378), .ZN(n132) );
  OAI21_X1 U145 ( .B1(n409), .B2(n378), .A(n133), .ZN(n262) );
  NAND2_X1 U146 ( .A1(\mem[6][6] ), .A2(n378), .ZN(n133) );
  OAI21_X1 U147 ( .B1(n408), .B2(n394), .A(n47), .ZN(n183) );
  NAND2_X1 U148 ( .A1(\mem[1][7] ), .A2(n393), .ZN(n47) );
  OAI21_X1 U149 ( .B1(n411), .B2(n393), .A(n44), .ZN(n180) );
  NAND2_X1 U150 ( .A1(\mem[1][4] ), .A2(n393), .ZN(n44) );
  OAI21_X1 U151 ( .B1(n410), .B2(n393), .A(n45), .ZN(n181) );
  NAND2_X1 U152 ( .A1(\mem[1][5] ), .A2(n393), .ZN(n45) );
  OAI21_X1 U153 ( .B1(n409), .B2(n393), .A(n46), .ZN(n182) );
  NAND2_X1 U154 ( .A1(\mem[1][6] ), .A2(n393), .ZN(n46) );
  OAI21_X1 U155 ( .B1(n408), .B2(n385), .A(n99), .ZN(n231) );
  NAND2_X1 U156 ( .A1(\mem[4][7] ), .A2(n384), .ZN(n99) );
  OAI21_X1 U157 ( .B1(n411), .B2(n384), .A(n96), .ZN(n228) );
  NAND2_X1 U158 ( .A1(\mem[4][4] ), .A2(n384), .ZN(n96) );
  OAI21_X1 U159 ( .B1(n410), .B2(n384), .A(n97), .ZN(n229) );
  NAND2_X1 U160 ( .A1(\mem[4][5] ), .A2(n384), .ZN(n97) );
  OAI21_X1 U161 ( .B1(n409), .B2(n384), .A(n98), .ZN(n230) );
  NAND2_X1 U162 ( .A1(\mem[4][6] ), .A2(n384), .ZN(n98) );
  OAI21_X1 U163 ( .B1(n407), .B2(n382), .A(n118), .ZN(n248) );
  NAND2_X1 U164 ( .A1(\mem[5][8] ), .A2(n380), .ZN(n118) );
  OAI21_X1 U165 ( .B1(n406), .B2(n382), .A(n119), .ZN(n249) );
  NAND2_X1 U166 ( .A1(\mem[5][9] ), .A2(n380), .ZN(n119) );
  OAI21_X1 U167 ( .B1(n402), .B2(n382), .A(n123), .ZN(n253) );
  NAND2_X1 U168 ( .A1(\mem[5][13] ), .A2(n380), .ZN(n123) );
  OAI21_X1 U169 ( .B1(n401), .B2(n382), .A(n124), .ZN(n254) );
  NAND2_X1 U170 ( .A1(\mem[5][14] ), .A2(n380), .ZN(n124) );
  OAI21_X1 U171 ( .B1(n415), .B2(n381), .A(n110), .ZN(n240) );
  NAND2_X1 U172 ( .A1(\mem[5][0] ), .A2(n380), .ZN(n110) );
  OAI21_X1 U173 ( .B1(n414), .B2(n381), .A(n111), .ZN(n241) );
  NAND2_X1 U174 ( .A1(\mem[5][1] ), .A2(n380), .ZN(n111) );
  OAI21_X1 U175 ( .B1(n413), .B2(n381), .A(n112), .ZN(n242) );
  NAND2_X1 U176 ( .A1(\mem[5][2] ), .A2(n380), .ZN(n112) );
  OAI21_X1 U177 ( .B1(n412), .B2(n381), .A(n113), .ZN(n243) );
  NAND2_X1 U178 ( .A1(\mem[5][3] ), .A2(n380), .ZN(n113) );
  OAI21_X1 U179 ( .B1(n405), .B2(n382), .A(n120), .ZN(n250) );
  NAND2_X1 U180 ( .A1(\mem[5][10] ), .A2(n380), .ZN(n120) );
  OAI21_X1 U181 ( .B1(n404), .B2(n382), .A(n121), .ZN(n251) );
  NAND2_X1 U182 ( .A1(\mem[5][11] ), .A2(n380), .ZN(n121) );
  OAI21_X1 U183 ( .B1(n403), .B2(n382), .A(n122), .ZN(n252) );
  NAND2_X1 U184 ( .A1(\mem[5][12] ), .A2(n380), .ZN(n122) );
  OAI21_X1 U185 ( .B1(n400), .B2(n381), .A(n125), .ZN(n255) );
  NAND2_X1 U186 ( .A1(\mem[5][15] ), .A2(n380), .ZN(n125) );
  OAI21_X1 U187 ( .B1(n407), .B2(n388), .A(n82), .ZN(n216) );
  NAND2_X1 U188 ( .A1(\mem[3][8] ), .A2(n386), .ZN(n82) );
  OAI21_X1 U189 ( .B1(n406), .B2(n388), .A(n83), .ZN(n217) );
  NAND2_X1 U190 ( .A1(\mem[3][9] ), .A2(n386), .ZN(n83) );
  OAI21_X1 U191 ( .B1(n402), .B2(n388), .A(n87), .ZN(n221) );
  NAND2_X1 U192 ( .A1(\mem[3][13] ), .A2(n386), .ZN(n87) );
  OAI21_X1 U193 ( .B1(n401), .B2(n388), .A(n88), .ZN(n222) );
  NAND2_X1 U194 ( .A1(\mem[3][14] ), .A2(n386), .ZN(n88) );
  OAI21_X1 U195 ( .B1(n415), .B2(n387), .A(n74), .ZN(n208) );
  NAND2_X1 U196 ( .A1(\mem[3][0] ), .A2(n386), .ZN(n74) );
  OAI21_X1 U197 ( .B1(n414), .B2(n387), .A(n75), .ZN(n209) );
  NAND2_X1 U198 ( .A1(\mem[3][1] ), .A2(n386), .ZN(n75) );
  OAI21_X1 U199 ( .B1(n413), .B2(n387), .A(n76), .ZN(n210) );
  NAND2_X1 U200 ( .A1(\mem[3][2] ), .A2(n386), .ZN(n76) );
  OAI21_X1 U201 ( .B1(n412), .B2(n387), .A(n77), .ZN(n211) );
  NAND2_X1 U202 ( .A1(\mem[3][3] ), .A2(n386), .ZN(n77) );
  OAI21_X1 U203 ( .B1(n405), .B2(n388), .A(n84), .ZN(n218) );
  NAND2_X1 U204 ( .A1(\mem[3][10] ), .A2(n386), .ZN(n84) );
  OAI21_X1 U205 ( .B1(n404), .B2(n388), .A(n85), .ZN(n219) );
  NAND2_X1 U206 ( .A1(\mem[3][11] ), .A2(n386), .ZN(n85) );
  OAI21_X1 U207 ( .B1(n403), .B2(n388), .A(n86), .ZN(n220) );
  NAND2_X1 U208 ( .A1(\mem[3][12] ), .A2(n386), .ZN(n86) );
  OAI21_X1 U209 ( .B1(n400), .B2(n387), .A(n89), .ZN(n223) );
  NAND2_X1 U210 ( .A1(\mem[3][15] ), .A2(n386), .ZN(n89) );
  OAI21_X1 U211 ( .B1(n407), .B2(n376), .A(n152), .ZN(n280) );
  NAND2_X1 U212 ( .A1(\mem[7][8] ), .A2(n374), .ZN(n152) );
  OAI21_X1 U213 ( .B1(n406), .B2(n376), .A(n153), .ZN(n281) );
  NAND2_X1 U214 ( .A1(\mem[7][9] ), .A2(n374), .ZN(n153) );
  OAI21_X1 U215 ( .B1(n402), .B2(n376), .A(n157), .ZN(n285) );
  NAND2_X1 U216 ( .A1(\mem[7][13] ), .A2(n374), .ZN(n157) );
  OAI21_X1 U217 ( .B1(n401), .B2(n376), .A(n158), .ZN(n286) );
  NAND2_X1 U218 ( .A1(\mem[7][14] ), .A2(n374), .ZN(n158) );
  OAI21_X1 U219 ( .B1(n415), .B2(n375), .A(n144), .ZN(n272) );
  NAND2_X1 U220 ( .A1(\mem[7][0] ), .A2(n374), .ZN(n144) );
  OAI21_X1 U221 ( .B1(n414), .B2(n375), .A(n145), .ZN(n273) );
  NAND2_X1 U222 ( .A1(\mem[7][1] ), .A2(n374), .ZN(n145) );
  OAI21_X1 U223 ( .B1(n413), .B2(n375), .A(n146), .ZN(n274) );
  NAND2_X1 U224 ( .A1(\mem[7][2] ), .A2(n374), .ZN(n146) );
  OAI21_X1 U225 ( .B1(n412), .B2(n375), .A(n147), .ZN(n275) );
  NAND2_X1 U226 ( .A1(\mem[7][3] ), .A2(n374), .ZN(n147) );
  OAI21_X1 U227 ( .B1(n405), .B2(n376), .A(n154), .ZN(n282) );
  NAND2_X1 U228 ( .A1(\mem[7][10] ), .A2(n374), .ZN(n154) );
  OAI21_X1 U229 ( .B1(n404), .B2(n376), .A(n155), .ZN(n283) );
  NAND2_X1 U230 ( .A1(\mem[7][11] ), .A2(n374), .ZN(n155) );
  OAI21_X1 U231 ( .B1(n403), .B2(n376), .A(n156), .ZN(n284) );
  NAND2_X1 U232 ( .A1(\mem[7][12] ), .A2(n374), .ZN(n156) );
  OAI21_X1 U233 ( .B1(n400), .B2(n375), .A(n159), .ZN(n287) );
  NAND2_X1 U234 ( .A1(\mem[7][15] ), .A2(n374), .ZN(n159) );
  OAI21_X1 U235 ( .B1(n407), .B2(n394), .A(n48), .ZN(n184) );
  NAND2_X1 U236 ( .A1(\mem[1][8] ), .A2(n392), .ZN(n48) );
  OAI21_X1 U237 ( .B1(n406), .B2(n394), .A(n49), .ZN(n185) );
  NAND2_X1 U238 ( .A1(\mem[1][9] ), .A2(n392), .ZN(n49) );
  OAI21_X1 U239 ( .B1(n402), .B2(n394), .A(n53), .ZN(n189) );
  NAND2_X1 U240 ( .A1(\mem[1][13] ), .A2(n392), .ZN(n53) );
  OAI21_X1 U241 ( .B1(n401), .B2(n394), .A(n54), .ZN(n190) );
  NAND2_X1 U242 ( .A1(\mem[1][14] ), .A2(n392), .ZN(n54) );
  OAI21_X1 U243 ( .B1(n415), .B2(n393), .A(n40), .ZN(n176) );
  NAND2_X1 U244 ( .A1(\mem[1][0] ), .A2(n392), .ZN(n40) );
  OAI21_X1 U245 ( .B1(n414), .B2(n393), .A(n41), .ZN(n177) );
  NAND2_X1 U246 ( .A1(\mem[1][1] ), .A2(n392), .ZN(n41) );
  OAI21_X1 U247 ( .B1(n413), .B2(n393), .A(n42), .ZN(n178) );
  NAND2_X1 U248 ( .A1(\mem[1][2] ), .A2(n392), .ZN(n42) );
  OAI21_X1 U249 ( .B1(n412), .B2(n393), .A(n43), .ZN(n179) );
  NAND2_X1 U250 ( .A1(\mem[1][3] ), .A2(n392), .ZN(n43) );
  OAI21_X1 U251 ( .B1(n405), .B2(n394), .A(n50), .ZN(n186) );
  NAND2_X1 U252 ( .A1(\mem[1][10] ), .A2(n392), .ZN(n50) );
  OAI21_X1 U253 ( .B1(n404), .B2(n394), .A(n51), .ZN(n187) );
  NAND2_X1 U254 ( .A1(\mem[1][11] ), .A2(n392), .ZN(n51) );
  OAI21_X1 U255 ( .B1(n403), .B2(n394), .A(n52), .ZN(n188) );
  NAND2_X1 U256 ( .A1(\mem[1][12] ), .A2(n392), .ZN(n52) );
  OAI21_X1 U257 ( .B1(n400), .B2(n393), .A(n55), .ZN(n191) );
  NAND2_X1 U258 ( .A1(\mem[1][15] ), .A2(n392), .ZN(n55) );
  OAI21_X1 U259 ( .B1(n407), .B2(n391), .A(n65), .ZN(n200) );
  NAND2_X1 U260 ( .A1(\mem[2][8] ), .A2(n389), .ZN(n65) );
  OAI21_X1 U261 ( .B1(n406), .B2(n391), .A(n66), .ZN(n201) );
  NAND2_X1 U262 ( .A1(\mem[2][9] ), .A2(n389), .ZN(n66) );
  OAI21_X1 U263 ( .B1(n402), .B2(n391), .A(n70), .ZN(n205) );
  NAND2_X1 U264 ( .A1(\mem[2][13] ), .A2(n389), .ZN(n70) );
  OAI21_X1 U265 ( .B1(n401), .B2(n391), .A(n71), .ZN(n206) );
  NAND2_X1 U266 ( .A1(\mem[2][14] ), .A2(n389), .ZN(n71) );
  OAI21_X1 U267 ( .B1(n415), .B2(n390), .A(n57), .ZN(n192) );
  NAND2_X1 U268 ( .A1(\mem[2][0] ), .A2(n389), .ZN(n57) );
  OAI21_X1 U269 ( .B1(n414), .B2(n390), .A(n58), .ZN(n193) );
  NAND2_X1 U270 ( .A1(\mem[2][1] ), .A2(n389), .ZN(n58) );
  OAI21_X1 U271 ( .B1(n413), .B2(n390), .A(n59), .ZN(n194) );
  NAND2_X1 U272 ( .A1(\mem[2][2] ), .A2(n389), .ZN(n59) );
  OAI21_X1 U273 ( .B1(n412), .B2(n390), .A(n60), .ZN(n195) );
  NAND2_X1 U274 ( .A1(\mem[2][3] ), .A2(n389), .ZN(n60) );
  OAI21_X1 U275 ( .B1(n405), .B2(n391), .A(n67), .ZN(n202) );
  NAND2_X1 U276 ( .A1(\mem[2][10] ), .A2(n389), .ZN(n67) );
  OAI21_X1 U277 ( .B1(n404), .B2(n391), .A(n68), .ZN(n203) );
  NAND2_X1 U278 ( .A1(\mem[2][11] ), .A2(n389), .ZN(n68) );
  OAI21_X1 U279 ( .B1(n403), .B2(n391), .A(n69), .ZN(n204) );
  NAND2_X1 U280 ( .A1(\mem[2][12] ), .A2(n389), .ZN(n69) );
  OAI21_X1 U281 ( .B1(n400), .B2(n390), .A(n72), .ZN(n207) );
  NAND2_X1 U290 ( .A1(\mem[2][15] ), .A2(n389), .ZN(n72) );
  OAI21_X1 U291 ( .B1(n396), .B2(n411), .A(n26), .ZN(n164) );
  NAND2_X1 U292 ( .A1(\mem[0][4] ), .A2(n396), .ZN(n26) );
  OAI21_X1 U293 ( .B1(n396), .B2(n410), .A(n27), .ZN(n165) );
  NAND2_X1 U294 ( .A1(\mem[0][5] ), .A2(n396), .ZN(n27) );
  OAI21_X1 U295 ( .B1(n396), .B2(n409), .A(n28), .ZN(n166) );
  NAND2_X1 U296 ( .A1(\mem[0][6] ), .A2(n396), .ZN(n28) );
  OAI21_X1 U297 ( .B1(n396), .B2(n408), .A(n29), .ZN(n167) );
  NAND2_X1 U298 ( .A1(\mem[0][7] ), .A2(n396), .ZN(n29) );
  OAI21_X1 U299 ( .B1(n407), .B2(n385), .A(n100), .ZN(n232) );
  NAND2_X1 U300 ( .A1(\mem[4][8] ), .A2(n383), .ZN(n100) );
  OAI21_X1 U301 ( .B1(n406), .B2(n385), .A(n101), .ZN(n233) );
  NAND2_X1 U302 ( .A1(\mem[4][9] ), .A2(n383), .ZN(n101) );
  OAI21_X1 U303 ( .B1(n402), .B2(n385), .A(n105), .ZN(n237) );
  NAND2_X1 U304 ( .A1(\mem[4][13] ), .A2(n383), .ZN(n105) );
  OAI21_X1 U305 ( .B1(n401), .B2(n385), .A(n106), .ZN(n238) );
  NAND2_X1 U306 ( .A1(\mem[4][14] ), .A2(n383), .ZN(n106) );
  OAI21_X1 U307 ( .B1(n415), .B2(n384), .A(n92), .ZN(n224) );
  NAND2_X1 U308 ( .A1(\mem[4][0] ), .A2(n383), .ZN(n92) );
  OAI21_X1 U309 ( .B1(n414), .B2(n384), .A(n93), .ZN(n225) );
  NAND2_X1 U310 ( .A1(\mem[4][1] ), .A2(n383), .ZN(n93) );
  OAI21_X1 U311 ( .B1(n413), .B2(n384), .A(n94), .ZN(n226) );
  NAND2_X1 U312 ( .A1(\mem[4][2] ), .A2(n383), .ZN(n94) );
  OAI21_X1 U313 ( .B1(n412), .B2(n384), .A(n95), .ZN(n227) );
  NAND2_X1 U314 ( .A1(\mem[4][3] ), .A2(n383), .ZN(n95) );
  OAI21_X1 U315 ( .B1(n405), .B2(n385), .A(n102), .ZN(n234) );
  NAND2_X1 U316 ( .A1(\mem[4][10] ), .A2(n383), .ZN(n102) );
  OAI21_X1 U317 ( .B1(n404), .B2(n385), .A(n103), .ZN(n235) );
  NAND2_X1 U318 ( .A1(\mem[4][11] ), .A2(n383), .ZN(n103) );
  OAI21_X1 U319 ( .B1(n403), .B2(n385), .A(n104), .ZN(n236) );
  NAND2_X1 U320 ( .A1(\mem[4][12] ), .A2(n383), .ZN(n104) );
  OAI21_X1 U321 ( .B1(n400), .B2(n384), .A(n107), .ZN(n239) );
  NAND2_X1 U322 ( .A1(\mem[4][15] ), .A2(n383), .ZN(n107) );
  MUX2_X1 U323 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n373), .Z(n3) );
  MUX2_X1 U324 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n370), .Z(n4) );
  MUX2_X1 U325 ( .A(n4), .B(n3), .S(n366), .Z(n5) );
  MUX2_X1 U326 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n369), .Z(n6) );
  MUX2_X1 U327 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n371), .Z(n7) );
  MUX2_X1 U328 ( .A(n7), .B(n6), .S(n366), .Z(n8) );
  MUX2_X1 U329 ( .A(n8), .B(n5), .S(N12), .Z(N28) );
  MUX2_X1 U330 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n369), .Z(n9) );
  MUX2_X1 U331 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n369), .Z(n10) );
  MUX2_X1 U332 ( .A(n10), .B(n9), .S(n366), .Z(n11) );
  MUX2_X1 U333 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n369), .Z(n12) );
  MUX2_X1 U334 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n369), .Z(n13) );
  MUX2_X1 U335 ( .A(n13), .B(n12), .S(n366), .Z(n14) );
  MUX2_X1 U336 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n369), .Z(n15) );
  MUX2_X1 U337 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n369), .Z(n16) );
  MUX2_X1 U338 ( .A(n16), .B(n15), .S(n366), .Z(n17) );
  MUX2_X1 U339 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n369), .Z(n18) );
  MUX2_X1 U340 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n369), .Z(n19) );
  MUX2_X1 U341 ( .A(n19), .B(n18), .S(n366), .Z(n20) );
  MUX2_X1 U342 ( .A(n20), .B(n17), .S(N12), .Z(N26) );
  MUX2_X1 U343 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n369), .Z(n288) );
  MUX2_X1 U344 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n369), .Z(n289) );
  MUX2_X1 U345 ( .A(n289), .B(n288), .S(n366), .Z(n290) );
  MUX2_X1 U346 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n369), .Z(n291) );
  MUX2_X1 U347 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n369), .Z(n292) );
  MUX2_X1 U348 ( .A(n292), .B(n291), .S(n366), .Z(n293) );
  MUX2_X1 U349 ( .A(n293), .B(n290), .S(N12), .Z(N25) );
  MUX2_X1 U350 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n370), .Z(n294) );
  MUX2_X1 U351 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n370), .Z(n295) );
  MUX2_X1 U352 ( .A(n295), .B(n294), .S(n367), .Z(n296) );
  MUX2_X1 U353 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n370), .Z(n297) );
  MUX2_X1 U354 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n370), .Z(n298) );
  MUX2_X1 U355 ( .A(n298), .B(n297), .S(n367), .Z(n299) );
  MUX2_X1 U356 ( .A(n299), .B(n296), .S(N12), .Z(N24) );
  MUX2_X1 U357 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n370), .Z(n300) );
  MUX2_X1 U358 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n370), .Z(n301) );
  MUX2_X1 U359 ( .A(n301), .B(n300), .S(n367), .Z(n302) );
  MUX2_X1 U360 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n370), .Z(n303) );
  MUX2_X1 U361 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n370), .Z(n304) );
  MUX2_X1 U362 ( .A(n304), .B(n303), .S(n367), .Z(n305) );
  MUX2_X1 U363 ( .A(n305), .B(n302), .S(N12), .Z(N23) );
  MUX2_X1 U364 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n370), .Z(n306) );
  MUX2_X1 U365 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n370), .Z(n307) );
  MUX2_X1 U366 ( .A(n307), .B(n306), .S(n367), .Z(n308) );
  MUX2_X1 U367 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n370), .Z(n309) );
  MUX2_X1 U368 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n370), .Z(n310) );
  MUX2_X1 U369 ( .A(n310), .B(n309), .S(n367), .Z(n311) );
  MUX2_X1 U370 ( .A(n311), .B(n308), .S(N12), .Z(N22) );
  MUX2_X1 U371 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n371), .Z(n312) );
  MUX2_X1 U372 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n371), .Z(n313) );
  MUX2_X1 U373 ( .A(n313), .B(n312), .S(n367), .Z(n314) );
  MUX2_X1 U374 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n371), .Z(n315) );
  MUX2_X1 U375 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n371), .Z(n316) );
  MUX2_X1 U376 ( .A(n316), .B(n315), .S(n367), .Z(n317) );
  MUX2_X1 U377 ( .A(n317), .B(n314), .S(N12), .Z(N21) );
  MUX2_X1 U378 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n371), .Z(n318) );
  MUX2_X1 U379 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n371), .Z(n319) );
  MUX2_X1 U380 ( .A(n319), .B(n318), .S(n367), .Z(n320) );
  MUX2_X1 U381 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n371), .Z(n321) );
  MUX2_X1 U382 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n371), .Z(n322) );
  MUX2_X1 U383 ( .A(n322), .B(n321), .S(n367), .Z(n323) );
  MUX2_X1 U384 ( .A(n323), .B(n320), .S(N12), .Z(N20) );
  MUX2_X1 U385 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n371), .Z(n324) );
  MUX2_X1 U386 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n371), .Z(n325) );
  MUX2_X1 U387 ( .A(n325), .B(n324), .S(n367), .Z(n326) );
  MUX2_X1 U388 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n371), .Z(n327) );
  MUX2_X1 U389 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n371), .Z(n328) );
  MUX2_X1 U390 ( .A(n328), .B(n327), .S(n367), .Z(n329) );
  MUX2_X1 U391 ( .A(n329), .B(n326), .S(N12), .Z(N19) );
  MUX2_X1 U392 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n372), .Z(n330) );
  MUX2_X1 U393 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n372), .Z(n331) );
  MUX2_X1 U394 ( .A(n331), .B(n330), .S(n368), .Z(n332) );
  MUX2_X1 U395 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n372), .Z(n333) );
  MUX2_X1 U396 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n372), .Z(n334) );
  MUX2_X1 U397 ( .A(n334), .B(n333), .S(n368), .Z(n335) );
  MUX2_X1 U398 ( .A(n335), .B(n332), .S(N12), .Z(N18) );
  MUX2_X1 U399 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n372), .Z(n336) );
  MUX2_X1 U400 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n372), .Z(n337) );
  MUX2_X1 U401 ( .A(n337), .B(n336), .S(n368), .Z(n338) );
  MUX2_X1 U402 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n372), .Z(n339) );
  MUX2_X1 U403 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n372), .Z(n340) );
  MUX2_X1 U404 ( .A(n340), .B(n339), .S(n368), .Z(n341) );
  MUX2_X1 U405 ( .A(n341), .B(n338), .S(N12), .Z(N17) );
  MUX2_X1 U406 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n372), .Z(n342) );
  MUX2_X1 U407 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n372), .Z(n343) );
  MUX2_X1 U408 ( .A(n343), .B(n342), .S(n368), .Z(n344) );
  MUX2_X1 U409 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n372), .Z(n345) );
  MUX2_X1 U410 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n372), .Z(n346) );
  MUX2_X1 U411 ( .A(n346), .B(n345), .S(n368), .Z(n347) );
  MUX2_X1 U412 ( .A(n347), .B(n344), .S(N12), .Z(N16) );
  MUX2_X1 U413 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n373), .Z(n348) );
  MUX2_X1 U414 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n373), .Z(n349) );
  MUX2_X1 U415 ( .A(n349), .B(n348), .S(n368), .Z(n350) );
  MUX2_X1 U416 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n373), .Z(n351) );
  MUX2_X1 U417 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n373), .Z(n352) );
  MUX2_X1 U418 ( .A(n352), .B(n351), .S(n368), .Z(n353) );
  MUX2_X1 U419 ( .A(n353), .B(n350), .S(N12), .Z(N15) );
  MUX2_X1 U420 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n373), .Z(n354) );
  MUX2_X1 U421 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n373), .Z(n355) );
  MUX2_X1 U422 ( .A(n355), .B(n354), .S(n368), .Z(n356) );
  MUX2_X1 U423 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n373), .Z(n357) );
  MUX2_X1 U424 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n373), .Z(n358) );
  MUX2_X1 U425 ( .A(n358), .B(n357), .S(n368), .Z(n359) );
  MUX2_X1 U426 ( .A(n359), .B(n356), .S(N12), .Z(N14) );
  MUX2_X1 U427 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n373), .Z(n360) );
  MUX2_X1 U428 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n373), .Z(n361) );
  MUX2_X1 U429 ( .A(n361), .B(n360), .S(n368), .Z(n362) );
  MUX2_X1 U430 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(n373), .Z(n363) );
  MUX2_X1 U431 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(n373), .Z(n364) );
  MUX2_X1 U432 ( .A(n364), .B(n363), .S(n368), .Z(n365) );
  MUX2_X1 U433 ( .A(n365), .B(n362), .S(N12), .Z(N13) );
endmodule


module layer2_12_8_12_16_W_rom_0 ( clk, addr, z );
  input [3:0] addr;
  output [15:0] z;
  input clk;
  wire   n11, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n12, n48, n49, n50, n51, n52, n53, n54, n55;

  DFF_X1 \z_reg[15]  ( .D(n47), .CK(clk), .Q(z[15]), .QN(n16) );
  DFF_X1 \z_reg[14]  ( .D(n46), .CK(clk), .Q(z[14]), .QN(n17) );
  DFF_X1 \z_reg[13]  ( .D(n45), .CK(clk), .Q(z[13]), .QN(n18) );
  DFF_X1 \z_reg[12]  ( .D(n44), .CK(clk), .Q(z[12]), .QN(n19) );
  DFF_X1 \z_reg[11]  ( .D(n43), .CK(clk), .Q(z[11]), .QN(n20) );
  DFF_X1 \z_reg[10]  ( .D(n42), .CK(clk), .Q(z[10]), .QN(n21) );
  DFF_X1 \z_reg[9]  ( .D(n41), .CK(clk), .Q(z[9]), .QN(n22) );
  DFF_X1 \z_reg[8]  ( .D(n40), .CK(clk), .Q(z[8]), .QN(n23) );
  DFF_X1 \z_reg[7]  ( .D(n39), .CK(clk), .Q(z[7]), .QN(n24) );
  DFF_X1 \z_reg[6]  ( .D(n38), .CK(clk), .Q(z[6]), .QN(n25) );
  DFF_X1 \z_reg[5]  ( .D(n37), .CK(clk), .Q(z[5]), .QN(n26) );
  DFF_X1 \z_reg[4]  ( .D(n36), .CK(clk), .Q(z[4]), .QN(n27) );
  DFF_X1 \z_reg[3]  ( .D(n35), .CK(clk), .Q(z[3]), .QN(n28) );
  DFF_X1 \z_reg[2]  ( .D(n34), .CK(clk), .Q(z[2]), .QN(n29) );
  DFF_X1 \z_reg[1]  ( .D(n33), .CK(clk), .Q(z[1]), .QN(n30) );
  DFF_X1 \z_reg[0]  ( .D(n32), .CK(clk), .Q(z[0]), .QN(n31) );
  OAI21_X1 U3 ( .B1(addr[2]), .B2(addr[0]), .A(n15), .ZN(n14) );
  OAI21_X1 U4 ( .B1(addr[0]), .B2(n55), .A(addr[2]), .ZN(n15) );
  INV_X1 U5 ( .A(addr[3]), .ZN(n54) );
  OAI21_X1 U6 ( .B1(n54), .B2(n19), .A(n13), .ZN(n44) );
  OAI21_X1 U7 ( .B1(n54), .B2(n18), .A(n13), .ZN(n45) );
  OAI21_X1 U8 ( .B1(n54), .B2(n17), .A(n13), .ZN(n46) );
  OAI21_X1 U9 ( .B1(n54), .B2(n16), .A(n13), .ZN(n47) );
  XNOR2_X1 U10 ( .A(addr[1]), .B(addr[2]), .ZN(n11) );
  INV_X1 U11 ( .A(addr[1]), .ZN(n55) );
  NAND2_X1 U12 ( .A1(n14), .A2(n54), .ZN(n13) );
  NAND2_X1 U13 ( .A1(addr[1]), .A2(n54), .ZN(n3) );
  INV_X1 U14 ( .A(n3), .ZN(n1) );
  INV_X1 U15 ( .A(addr[2]), .ZN(n8) );
  NAND2_X1 U16 ( .A1(n1), .A2(n8), .ZN(n52) );
  INV_X1 U17 ( .A(n52), .ZN(n2) );
  NAND2_X1 U18 ( .A1(addr[0]), .A2(n2), .ZN(n7) );
  INV_X1 U19 ( .A(addr[0]), .ZN(n5) );
  NAND3_X1 U20 ( .A1(n11), .A2(n54), .A3(n5), .ZN(n48) );
  OAI211_X1 U21 ( .C1(n31), .C2(n54), .A(n7), .B(n48), .ZN(n32) );
  NAND2_X1 U22 ( .A1(addr[2]), .A2(n54), .ZN(n49) );
  MUX2_X1 U23 ( .A(n3), .B(n49), .S(addr[0]), .Z(n4) );
  OAI21_X1 U24 ( .B1(n30), .B2(n54), .A(n4), .ZN(n33) );
  MUX2_X1 U25 ( .A(n5), .B(n29), .S(addr[3]), .Z(n6) );
  NAND2_X1 U26 ( .A1(n49), .A2(n6), .ZN(n34) );
  OAI221_X1 U27 ( .B1(addr[0]), .B2(n49), .C1(n28), .C2(n54), .A(n7), .ZN(n35)
         );
  MUX2_X1 U28 ( .A(n8), .B(n55), .S(addr[0]), .Z(n9) );
  AOI21_X1 U29 ( .B1(addr[2]), .B2(addr[1]), .A(n9), .ZN(n10) );
  MUX2_X1 U30 ( .A(n10), .B(n27), .S(addr[3]), .Z(n12) );
  INV_X1 U31 ( .A(n12), .ZN(n36) );
  OAI21_X1 U32 ( .B1(n26), .B2(n54), .A(n48), .ZN(n37) );
  INV_X1 U33 ( .A(n49), .ZN(n50) );
  NAND2_X1 U34 ( .A1(n50), .A2(n55), .ZN(n51) );
  MUX2_X1 U35 ( .A(n52), .B(n51), .S(addr[0]), .Z(n53) );
  OAI21_X1 U36 ( .B1(n25), .B2(n54), .A(n53), .ZN(n38) );
  OAI21_X1 U37 ( .B1(n24), .B2(n54), .A(n13), .ZN(n39) );
  OAI21_X1 U38 ( .B1(n23), .B2(n54), .A(n13), .ZN(n40) );
  OAI21_X1 U39 ( .B1(n22), .B2(n54), .A(n13), .ZN(n41) );
  OAI21_X1 U40 ( .B1(n21), .B2(n54), .A(n13), .ZN(n42) );
  OAI21_X1 U41 ( .B1(n20), .B2(n54), .A(n13), .ZN(n43) );
endmodule


module layer2_12_8_12_16_B_rom_0 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b1;
  assign z[14] = 1'b1;
  assign z[13] = 1'b1;
  assign z[12] = 1'b1;
  assign z[11] = 1'b1;
  assign z[10] = 1'b1;
  assign z[9] = 1'b1;
  assign z[8] = 1'b1;
  assign z[7] = 1'b1;
  assign z[6] = 1'b1;
  assign z[5] = 1'b0;
  assign z[4] = 1'b1;
  assign z[3] = 1'b0;
  assign z[2] = 1'b0;
  assign z[1] = 1'b1;
  assign z[0] = 1'b1;

endmodule


module layer2_12_8_12_16_W_rom_1 ( clk, addr, z );
  input [3:0] addr;
  output [15:0] z;
  input clk;
  wire   n4, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n1, n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n44, n45, n46, n47, n48;

  DFF_X1 \z_reg[15]  ( .D(n43), .CK(clk), .Q(z[15]), .QN(n14) );
  DFF_X1 \z_reg[14]  ( .D(n42), .CK(clk), .Q(z[14]), .QN(n15) );
  DFF_X1 \z_reg[13]  ( .D(n41), .CK(clk), .Q(z[13]), .QN(n16) );
  DFF_X1 \z_reg[12]  ( .D(n40), .CK(clk), .Q(z[12]), .QN(n17) );
  DFF_X1 \z_reg[11]  ( .D(n39), .CK(clk), .Q(z[11]), .QN(n18) );
  DFF_X1 \z_reg[10]  ( .D(n38), .CK(clk), .Q(z[10]), .QN(n19) );
  DFF_X1 \z_reg[9]  ( .D(n37), .CK(clk), .Q(z[9]), .QN(n20) );
  DFF_X1 \z_reg[8]  ( .D(n36), .CK(clk), .Q(z[8]), .QN(n21) );
  DFF_X1 \z_reg[7]  ( .D(n35), .CK(clk), .Q(z[7]), .QN(n22) );
  DFF_X1 \z_reg[6]  ( .D(n34), .CK(clk), .Q(z[6]), .QN(n1) );
  DFF_X1 \z_reg[5]  ( .D(n33), .CK(clk), .Q(z[5]), .QN(n23) );
  DFF_X1 \z_reg[4]  ( .D(n32), .CK(clk), .Q(z[4]), .QN(n24) );
  DFF_X1 \z_reg[3]  ( .D(n31), .CK(clk), .Q(z[3]), .QN(n25) );
  DFF_X1 \z_reg[2]  ( .D(n30), .CK(clk), .Q(z[2]), .QN(n26) );
  DFF_X1 \z_reg[1]  ( .D(n29), .CK(clk), .Q(z[1]) );
  DFF_X1 \z_reg[0]  ( .D(n28), .CK(clk), .Q(z[0]), .QN(n27) );
  INV_X1 U3 ( .A(addr[3]), .ZN(n48) );
  OAI21_X1 U4 ( .B1(n48), .B2(n17), .A(n4), .ZN(n40) );
  OAI21_X1 U5 ( .B1(n48), .B2(n16), .A(n4), .ZN(n41) );
  OAI21_X1 U6 ( .B1(n48), .B2(n15), .A(n4), .ZN(n42) );
  OAI21_X1 U7 ( .B1(n48), .B2(n14), .A(n4), .ZN(n43) );
  INV_X1 U8 ( .A(addr[2]), .ZN(n10) );
  NAND2_X1 U9 ( .A1(addr[1]), .A2(n10), .ZN(n9) );
  INV_X1 U10 ( .A(n9), .ZN(n47) );
  NAND2_X1 U11 ( .A1(n47), .A2(n48), .ZN(n4) );
  INV_X1 U12 ( .A(addr[0]), .ZN(n2) );
  NAND2_X1 U13 ( .A1(n48), .A2(n2), .ZN(n46) );
  INV_X1 U14 ( .A(n46), .ZN(n6) );
  NAND2_X1 U15 ( .A1(n6), .A2(addr[1]), .ZN(n11) );
  NAND3_X1 U16 ( .A1(addr[0]), .A2(addr[2]), .A3(n48), .ZN(n44) );
  OAI211_X1 U17 ( .C1(n27), .C2(n48), .A(n11), .B(n44), .ZN(n28) );
  INV_X1 U18 ( .A(addr[1]), .ZN(n7) );
  NAND3_X1 U19 ( .A1(addr[2]), .A2(n48), .A3(n7), .ZN(n45) );
  INV_X1 U20 ( .A(n44), .ZN(n3) );
  AOI21_X1 U21 ( .B1(z[1]), .B2(addr[3]), .A(n3), .ZN(n5) );
  NAND3_X1 U22 ( .A1(n45), .A2(n4), .A3(n5), .ZN(n29) );
  OAI21_X1 U23 ( .B1(n7), .B2(n10), .A(n6), .ZN(n8) );
  OAI21_X1 U24 ( .B1(n26), .B2(n48), .A(n8), .ZN(n30) );
  OAI21_X1 U25 ( .B1(addr[1]), .B2(n10), .A(n9), .ZN(n12) );
  OAI222_X1 U26 ( .A1(addr[1]), .A2(n44), .B1(n46), .B2(n12), .C1(n25), .C2(
        n48), .ZN(n31) );
  OAI211_X1 U27 ( .C1(n24), .C2(n48), .A(n11), .B(n45), .ZN(n32) );
  MUX2_X1 U28 ( .A(n12), .B(n23), .S(addr[3]), .Z(n13) );
  NAND2_X1 U29 ( .A1(n44), .A2(n13), .ZN(n33) );
  OAI221_X1 U30 ( .B1(n47), .B2(n46), .C1(n48), .C2(n1), .A(n45), .ZN(n34) );
  OAI21_X1 U31 ( .B1(n22), .B2(n48), .A(n4), .ZN(n35) );
  OAI21_X1 U32 ( .B1(n21), .B2(n48), .A(n4), .ZN(n36) );
  OAI21_X1 U33 ( .B1(n20), .B2(n48), .A(n4), .ZN(n37) );
  OAI21_X1 U34 ( .B1(n19), .B2(n48), .A(n4), .ZN(n38) );
  OAI21_X1 U35 ( .B1(n18), .B2(n48), .A(n4), .ZN(n39) );
endmodule


module layer2_12_8_12_16_B_rom_1 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b1;
  assign z[14] = 1'b1;
  assign z[13] = 1'b1;
  assign z[12] = 1'b1;
  assign z[11] = 1'b1;
  assign z[10] = 1'b1;
  assign z[9] = 1'b1;
  assign z[8] = 1'b1;
  assign z[7] = 1'b1;
  assign z[6] = 1'b0;
  assign z[5] = 1'b0;
  assign z[4] = 1'b1;
  assign z[3] = 1'b1;
  assign z[2] = 1'b0;
  assign z[1] = 1'b1;
  assign z[0] = 1'b1;

endmodule


module layer2_12_8_12_16_W_rom_2 ( clk, addr, z );
  input [3:0] addr;
  output [15:0] z;
  input clk;
  wire   n5, n10, n13, n14, n16, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n1, n2, n3, n4, n6,
         n7, n8, n9, n11, n12, n15, n17, n51, n52, n53, n54, n55, n56, n57,
         n58;

  DFF_X1 \z_reg[15]  ( .D(n50), .CK(clk), .Q(z[15]), .QN(n19) );
  DFF_X1 \z_reg[14]  ( .D(n49), .CK(clk), .Q(z[14]), .QN(n20) );
  DFF_X1 \z_reg[13]  ( .D(n48), .CK(clk), .Q(z[13]), .QN(n21) );
  DFF_X1 \z_reg[12]  ( .D(n47), .CK(clk), .Q(z[12]), .QN(n22) );
  DFF_X1 \z_reg[11]  ( .D(n46), .CK(clk), .Q(z[11]), .QN(n23) );
  DFF_X1 \z_reg[10]  ( .D(n45), .CK(clk), .Q(z[10]), .QN(n24) );
  DFF_X1 \z_reg[9]  ( .D(n44), .CK(clk), .Q(z[9]), .QN(n25) );
  DFF_X1 \z_reg[8]  ( .D(n43), .CK(clk), .Q(z[8]), .QN(n26) );
  DFF_X1 \z_reg[7]  ( .D(n42), .CK(clk), .Q(z[7]), .QN(n27) );
  DFF_X1 \z_reg[6]  ( .D(n41), .CK(clk), .Q(z[6]), .QN(n28) );
  DFF_X1 \z_reg[5]  ( .D(n40), .CK(clk), .Q(z[5]), .QN(n29) );
  DFF_X1 \z_reg[4]  ( .D(n39), .CK(clk), .Q(z[4]), .QN(n30) );
  DFF_X1 \z_reg[3]  ( .D(n38), .CK(clk), .Q(z[3]), .QN(n31) );
  DFF_X1 \z_reg[2]  ( .D(n37), .CK(clk), .Q(z[2]), .QN(n32) );
  DFF_X1 \z_reg[1]  ( .D(n36), .CK(clk), .Q(z[1]), .QN(n33) );
  DFF_X1 \z_reg[0]  ( .D(n35), .CK(clk), .Q(z[0]), .QN(n34) );
  AND2_X1 U3 ( .A1(addr[2]), .A2(addr[1]), .ZN(n1) );
  AND2_X1 U4 ( .A1(n1), .A2(n58), .ZN(n2) );
  NAND2_X1 U5 ( .A1(n56), .A2(n58), .ZN(n10) );
  NAND3_X1 U6 ( .A1(n14), .A2(addr[2]), .A3(n55), .ZN(n18) );
  OAI21_X1 U7 ( .B1(n55), .B2(n22), .A(n18), .ZN(n47) );
  OAI21_X1 U8 ( .B1(n55), .B2(n21), .A(n18), .ZN(n48) );
  OAI21_X1 U9 ( .B1(n55), .B2(n20), .A(n18), .ZN(n49) );
  OAI21_X1 U10 ( .B1(n55), .B2(n19), .A(n18), .ZN(n50) );
  NAND2_X1 U11 ( .A1(addr[0]), .A2(addr[1]), .ZN(n14) );
  XNOR2_X1 U12 ( .A(n14), .B(n56), .ZN(n13) );
  NAND2_X1 U13 ( .A1(n57), .A2(n58), .ZN(n5) );
  NOR3_X1 U14 ( .A1(n58), .A2(addr[2]), .A3(addr[1]), .ZN(n16) );
  INV_X1 U15 ( .A(addr[3]), .ZN(n55) );
  INV_X1 U16 ( .A(addr[2]), .ZN(n56) );
  INV_X1 U17 ( .A(addr[0]), .ZN(n58) );
  INV_X1 U18 ( .A(addr[1]), .ZN(n57) );
  NOR2_X1 U19 ( .A1(addr[0]), .A2(n1), .ZN(n3) );
  MUX2_X1 U20 ( .A(n3), .B(n34), .S(addr[3]), .Z(n4) );
  INV_X1 U21 ( .A(n4), .ZN(n35) );
  MUX2_X1 U22 ( .A(n2), .B(n33), .S(addr[3]), .Z(n6) );
  INV_X1 U23 ( .A(n6), .ZN(n36) );
  MUX2_X1 U24 ( .A(n5), .B(n58), .S(addr[2]), .Z(n8) );
  INV_X1 U25 ( .A(n32), .ZN(n7) );
  MUX2_X1 U26 ( .A(n8), .B(n7), .S(addr[3]), .Z(n37) );
  OAI22_X1 U27 ( .A1(n58), .A2(n56), .B1(n10), .B2(n57), .ZN(n52) );
  AOI21_X1 U28 ( .B1(n10), .B2(n57), .A(n52), .ZN(n9) );
  MUX2_X1 U29 ( .A(n9), .B(n31), .S(addr[3]), .Z(n11) );
  INV_X1 U30 ( .A(n11), .ZN(n38) );
  AOI21_X1 U31 ( .B1(n58), .B2(n57), .A(n13), .ZN(n12) );
  MUX2_X1 U32 ( .A(n12), .B(n30), .S(addr[3]), .Z(n15) );
  INV_X1 U33 ( .A(n15), .ZN(n39) );
  NOR2_X1 U34 ( .A1(n16), .A2(n2), .ZN(n17) );
  MUX2_X1 U35 ( .A(n17), .B(n29), .S(addr[3]), .Z(n51) );
  INV_X1 U36 ( .A(n51), .ZN(n40) );
  INV_X1 U37 ( .A(n52), .ZN(n53) );
  MUX2_X1 U38 ( .A(n53), .B(n28), .S(addr[3]), .Z(n54) );
  INV_X1 U39 ( .A(n54), .ZN(n41) );
  OAI21_X1 U40 ( .B1(n27), .B2(n55), .A(n18), .ZN(n42) );
  OAI21_X1 U41 ( .B1(n26), .B2(n55), .A(n18), .ZN(n43) );
  OAI21_X1 U42 ( .B1(n25), .B2(n55), .A(n18), .ZN(n44) );
  OAI21_X1 U43 ( .B1(n24), .B2(n55), .A(n18), .ZN(n45) );
  OAI21_X1 U44 ( .B1(n23), .B2(n55), .A(n18), .ZN(n46) );
endmodule


module layer2_12_8_12_16_B_rom_2 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b1;
  assign z[14] = 1'b1;
  assign z[13] = 1'b1;
  assign z[12] = 1'b1;
  assign z[11] = 1'b1;
  assign z[10] = 1'b1;
  assign z[9] = 1'b1;
  assign z[8] = 1'b1;
  assign z[7] = 1'b1;
  assign z[6] = 1'b0;
  assign z[5] = 1'b0;
  assign z[4] = 1'b0;
  assign z[3] = 1'b0;
  assign z[2] = 1'b0;
  assign z[1] = 1'b1;
  assign z[0] = 1'b0;

endmodule


module layer2_12_8_12_16_W_rom_3 ( clk, addr, z );
  input [3:0] addr;
  output [15:0] z;
  input clk;
  wire   n7, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n1, n2, n3, n4, n5, n6, n8, n41, n42, n43,
         n44, n45, n46;

  DFF_X1 \z_reg[15]  ( .D(n40), .CK(clk), .Q(z[15]), .QN(n9) );
  DFF_X1 \z_reg[14]  ( .D(n39), .CK(clk), .Q(z[14]), .QN(n10) );
  DFF_X1 \z_reg[13]  ( .D(n38), .CK(clk), .Q(z[13]), .QN(n11) );
  DFF_X1 \z_reg[12]  ( .D(n37), .CK(clk), .Q(z[12]), .QN(n12) );
  DFF_X1 \z_reg[11]  ( .D(n36), .CK(clk), .Q(z[11]), .QN(n13) );
  DFF_X1 \z_reg[10]  ( .D(n35), .CK(clk), .Q(z[10]), .QN(n14) );
  DFF_X1 \z_reg[9]  ( .D(n34), .CK(clk), .Q(z[9]), .QN(n15) );
  DFF_X1 \z_reg[8]  ( .D(n33), .CK(clk), .Q(z[8]), .QN(n16) );
  DFF_X1 \z_reg[7]  ( .D(n32), .CK(clk), .Q(z[7]), .QN(n17) );
  DFF_X1 \z_reg[6]  ( .D(n31), .CK(clk), .Q(z[6]), .QN(n18) );
  DFF_X1 \z_reg[5]  ( .D(n30), .CK(clk), .Q(z[5]), .QN(n19) );
  DFF_X1 \z_reg[4]  ( .D(n29), .CK(clk), .Q(z[4]), .QN(n20) );
  DFF_X1 \z_reg[3]  ( .D(n28), .CK(clk), .Q(z[3]), .QN(n21) );
  DFF_X1 \z_reg[2]  ( .D(n27), .CK(clk), .Q(z[2]), .QN(n22) );
  DFF_X1 \z_reg[1]  ( .D(n26), .CK(clk), .Q(z[1]), .QN(n23) );
  DFF_X1 \z_reg[0]  ( .D(n25), .CK(clk), .Q(z[0]), .QN(n24) );
  XNOR2_X1 U3 ( .A(n41), .B(addr[0]), .ZN(n1) );
  INV_X1 U4 ( .A(addr[3]), .ZN(n46) );
  OAI21_X1 U5 ( .B1(n46), .B2(n12), .A(n7), .ZN(n37) );
  OAI21_X1 U6 ( .B1(n46), .B2(n11), .A(n7), .ZN(n38) );
  OAI21_X1 U7 ( .B1(n46), .B2(n10), .A(n7), .ZN(n39) );
  OAI21_X1 U8 ( .B1(n46), .B2(n9), .A(n7), .ZN(n40) );
  INV_X1 U9 ( .A(addr[2]), .ZN(n41) );
  INV_X1 U10 ( .A(addr[1]), .ZN(n2) );
  NAND3_X1 U11 ( .A1(n46), .A2(n41), .A3(n2), .ZN(n7) );
  NAND2_X1 U12 ( .A1(addr[2]), .A2(n46), .ZN(n43) );
  INV_X1 U13 ( .A(n43), .ZN(n3) );
  NAND2_X1 U14 ( .A1(n3), .A2(n2), .ZN(n42) );
  MUX2_X1 U15 ( .A(addr[0]), .B(n24), .S(addr[3]), .Z(n4) );
  NAND2_X1 U16 ( .A1(n42), .A2(n4), .ZN(n25) );
  NAND2_X1 U17 ( .A1(addr[1]), .A2(n46), .ZN(n44) );
  INV_X1 U18 ( .A(n44), .ZN(n5) );
  NAND2_X1 U19 ( .A1(n5), .A2(n41), .ZN(n6) );
  MUX2_X1 U20 ( .A(n42), .B(n6), .S(addr[0]), .Z(n8) );
  OAI21_X1 U21 ( .B1(n23), .B2(n46), .A(n8), .ZN(n26) );
  OAI22_X1 U22 ( .A1(n1), .A2(n44), .B1(n22), .B2(n46), .ZN(n27) );
  OAI22_X1 U23 ( .A1(addr[0]), .A2(n7), .B1(n21), .B2(n46), .ZN(n28) );
  OAI221_X1 U24 ( .B1(addr[0]), .B2(n43), .C1(n20), .C2(n46), .A(n42), .ZN(n29) );
  OAI221_X1 U25 ( .B1(addr[0]), .B2(n44), .C1(n19), .C2(n46), .A(n43), .ZN(n30) );
  MUX2_X1 U26 ( .A(n1), .B(n18), .S(addr[3]), .Z(n45) );
  NAND2_X1 U27 ( .A1(n7), .A2(n45), .ZN(n31) );
  OAI21_X1 U28 ( .B1(n17), .B2(n46), .A(n7), .ZN(n32) );
  OAI21_X1 U29 ( .B1(n16), .B2(n46), .A(n7), .ZN(n33) );
  OAI21_X1 U30 ( .B1(n15), .B2(n46), .A(n7), .ZN(n34) );
  OAI21_X1 U31 ( .B1(n14), .B2(n46), .A(n7), .ZN(n35) );
  OAI21_X1 U32 ( .B1(n13), .B2(n46), .A(n7), .ZN(n36) );
endmodule


module layer2_12_8_12_16_B_rom_3 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b0;
  assign z[14] = 1'b0;
  assign z[13] = 1'b0;
  assign z[12] = 1'b0;
  assign z[11] = 1'b0;
  assign z[10] = 1'b0;
  assign z[9] = 1'b0;
  assign z[8] = 1'b0;
  assign z[7] = 1'b0;
  assign z[6] = 1'b1;
  assign z[5] = 1'b0;
  assign z[4] = 1'b0;
  assign z[3] = 1'b0;
  assign z[2] = 1'b1;
  assign z[1] = 1'b1;
  assign z[0] = 1'b0;

endmodule


module layer2_12_8_12_16_W_rom_4 ( clk, addr, z );
  input [3:0] addr;
  output [15:0] z;
  input clk;
  wire   n3, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n1, n2, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n52, n53;

  DFF_X1 \z_reg[15]  ( .D(n51), .CK(clk), .Q(z[15]), .QN(n20) );
  DFF_X1 \z_reg[14]  ( .D(n50), .CK(clk), .Q(z[14]), .QN(n21) );
  DFF_X1 \z_reg[13]  ( .D(n49), .CK(clk), .Q(z[13]), .QN(n22) );
  DFF_X1 \z_reg[12]  ( .D(n48), .CK(clk), .Q(z[12]), .QN(n23) );
  DFF_X1 \z_reg[11]  ( .D(n47), .CK(clk), .Q(z[11]), .QN(n24) );
  DFF_X1 \z_reg[10]  ( .D(n46), .CK(clk), .Q(z[10]), .QN(n25) );
  DFF_X1 \z_reg[9]  ( .D(n45), .CK(clk), .Q(z[9]), .QN(n26) );
  DFF_X1 \z_reg[8]  ( .D(n44), .CK(clk), .Q(z[8]), .QN(n27) );
  DFF_X1 \z_reg[7]  ( .D(n43), .CK(clk), .Q(z[7]), .QN(n28) );
  DFF_X1 \z_reg[6]  ( .D(n42), .CK(clk), .Q(z[6]), .QN(n29) );
  DFF_X1 \z_reg[5]  ( .D(n41), .CK(clk), .Q(z[5]), .QN(n30) );
  DFF_X1 \z_reg[4]  ( .D(n40), .CK(clk), .Q(z[4]), .QN(n31) );
  DFF_X1 \z_reg[3]  ( .D(n39), .CK(clk), .Q(z[3]), .QN(n32) );
  DFF_X1 \z_reg[2]  ( .D(n38), .CK(clk), .Q(z[2]), .QN(n33) );
  DFF_X1 \z_reg[1]  ( .D(n37), .CK(clk), .Q(z[1]), .QN(n34) );
  DFF_X1 \z_reg[0]  ( .D(n36), .CK(clk), .Q(z[0]), .QN(n35) );
  XOR2_X1 U34 ( .A(n3), .B(addr[0]), .Z(n19) );
  AND2_X1 U3 ( .A1(addr[2]), .A2(n52), .ZN(n1) );
  INV_X1 U4 ( .A(addr[3]), .ZN(n52) );
  OAI21_X1 U5 ( .B1(addr[1]), .B2(n53), .A(n19), .ZN(n18) );
  OAI21_X1 U6 ( .B1(n52), .B2(n23), .A(n17), .ZN(n48) );
  OAI21_X1 U7 ( .B1(n52), .B2(n22), .A(n17), .ZN(n49) );
  OAI21_X1 U8 ( .B1(n52), .B2(n21), .A(n17), .ZN(n50) );
  OAI21_X1 U9 ( .B1(n52), .B2(n20), .A(n17), .ZN(n51) );
  NAND2_X1 U10 ( .A1(addr[1]), .A2(n53), .ZN(n3) );
  INV_X1 U11 ( .A(addr[2]), .ZN(n53) );
  NAND2_X1 U12 ( .A1(n18), .A2(n52), .ZN(n17) );
  NOR2_X1 U13 ( .A1(n3), .A2(addr[0]), .ZN(n2) );
  MUX2_X1 U14 ( .A(n2), .B(n35), .S(addr[3]), .Z(n4) );
  INV_X1 U15 ( .A(n4), .ZN(n36) );
  INV_X1 U16 ( .A(addr[0]), .ZN(n6) );
  INV_X1 U17 ( .A(addr[1]), .ZN(n10) );
  NAND3_X1 U18 ( .A1(n53), .A2(n52), .A3(n10), .ZN(n5) );
  NAND3_X1 U19 ( .A1(addr[1]), .A2(n52), .A3(n6), .ZN(n11) );
  OAI221_X1 U20 ( .B1(n6), .B2(n5), .C1(n34), .C2(n52), .A(n11), .ZN(n37) );
  NAND2_X1 U21 ( .A1(addr[1]), .A2(n1), .ZN(n14) );
  OAI221_X1 U22 ( .B1(addr[0]), .B2(n5), .C1(n33), .C2(n52), .A(n14), .ZN(n38)
         );
  NAND3_X1 U23 ( .A1(n1), .A2(n10), .A3(n6), .ZN(n7) );
  OAI21_X1 U24 ( .B1(n32), .B2(n52), .A(n7), .ZN(n39) );
  OAI21_X1 U25 ( .B1(addr[1]), .B2(n53), .A(n3), .ZN(n13) );
  INV_X1 U26 ( .A(n13), .ZN(n8) );
  MUX2_X1 U27 ( .A(n8), .B(n31), .S(addr[3]), .Z(n9) );
  INV_X1 U28 ( .A(n9), .ZN(n40) );
  NAND3_X1 U29 ( .A1(addr[0]), .A2(n1), .A3(n10), .ZN(n12) );
  OAI211_X1 U30 ( .C1(n30), .C2(n52), .A(n12), .B(n11), .ZN(n41) );
  NAND2_X1 U31 ( .A1(n13), .A2(n52), .ZN(n15) );
  MUX2_X1 U32 ( .A(n15), .B(n14), .S(addr[0]), .Z(n16) );
  OAI21_X1 U33 ( .B1(n29), .B2(n52), .A(n16), .ZN(n42) );
  OAI21_X1 U35 ( .B1(n28), .B2(n52), .A(n17), .ZN(n43) );
  OAI21_X1 U36 ( .B1(n27), .B2(n52), .A(n17), .ZN(n44) );
  OAI21_X1 U37 ( .B1(n26), .B2(n52), .A(n17), .ZN(n45) );
  OAI21_X1 U38 ( .B1(n25), .B2(n52), .A(n17), .ZN(n46) );
  OAI21_X1 U39 ( .B1(n24), .B2(n52), .A(n17), .ZN(n47) );
endmodule


module layer2_12_8_12_16_B_rom_4 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b0;
  assign z[14] = 1'b0;
  assign z[13] = 1'b0;
  assign z[12] = 1'b0;
  assign z[11] = 1'b0;
  assign z[10] = 1'b0;
  assign z[9] = 1'b0;
  assign z[8] = 1'b0;
  assign z[7] = 1'b0;
  assign z[6] = 1'b0;
  assign z[5] = 1'b1;
  assign z[4] = 1'b0;
  assign z[3] = 1'b1;
  assign z[2] = 1'b0;
  assign z[1] = 1'b0;
  assign z[0] = 1'b1;

endmodule


module layer2_12_8_12_16_W_rom_5 ( clk, addr, z );
  input [3:0] addr;
  output [15:0] z;
  input clk;
  wire   n17, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n18, n50, n51, n52, n53, n54, n55;

  DFF_X1 \z_reg[15]  ( .D(n49), .CK(clk), .Q(z[15]), .QN(n19) );
  DFF_X1 \z_reg[14]  ( .D(n48), .CK(clk), .Q(z[14]), .QN(n20) );
  DFF_X1 \z_reg[13]  ( .D(n47), .CK(clk), .Q(z[13]), .QN(n21) );
  DFF_X1 \z_reg[12]  ( .D(n46), .CK(clk), .Q(z[12]), .QN(n22) );
  DFF_X1 \z_reg[11]  ( .D(n45), .CK(clk), .Q(z[11]), .QN(n23) );
  DFF_X1 \z_reg[10]  ( .D(n44), .CK(clk), .Q(z[10]), .QN(n24) );
  DFF_X1 \z_reg[9]  ( .D(n43), .CK(clk), .Q(z[9]), .QN(n25) );
  DFF_X1 \z_reg[8]  ( .D(n42), .CK(clk), .Q(z[8]), .QN(n26) );
  DFF_X1 \z_reg[7]  ( .D(n41), .CK(clk), .Q(z[7]), .QN(n27) );
  DFF_X1 \z_reg[6]  ( .D(n40), .CK(clk), .Q(z[6]), .QN(n28) );
  DFF_X1 \z_reg[5]  ( .D(n39), .CK(clk), .Q(z[5]), .QN(n29) );
  DFF_X1 \z_reg[4]  ( .D(n38), .CK(clk), .Q(z[4]), .QN(n30) );
  DFF_X1 \z_reg[3]  ( .D(n37), .CK(clk), .Q(z[3]), .QN(n31) );
  DFF_X1 \z_reg[2]  ( .D(n36), .CK(clk), .Q(z[2]), .QN(n32) );
  DFF_X1 \z_reg[1]  ( .D(n35), .CK(clk), .Q(z[1]) );
  DFF_X1 \z_reg[0]  ( .D(n34), .CK(clk), .Q(z[0]), .QN(n33) );
  AND2_X1 U3 ( .A1(addr[1]), .A2(n53), .ZN(n1) );
  AND2_X1 U4 ( .A1(n4), .A2(n11), .ZN(n2) );
  NOR2_X1 U5 ( .A1(n54), .A2(n55), .ZN(n17) );
  INV_X1 U6 ( .A(addr[3]), .ZN(n53) );
  INV_X1 U7 ( .A(n3), .ZN(n52) );
  OAI21_X1 U8 ( .B1(n53), .B2(n22), .A(n52), .ZN(n46) );
  OAI21_X1 U9 ( .B1(n53), .B2(n21), .A(n52), .ZN(n47) );
  OAI21_X1 U10 ( .B1(n53), .B2(n20), .A(n52), .ZN(n48) );
  OAI21_X1 U11 ( .B1(n53), .B2(n19), .A(n52), .ZN(n49) );
  INV_X1 U12 ( .A(addr[2]), .ZN(n54) );
  INV_X1 U13 ( .A(addr[0]), .ZN(n55) );
  INV_X1 U14 ( .A(n17), .ZN(n16) );
  NAND2_X1 U15 ( .A1(n1), .A2(n55), .ZN(n7) );
  OAI21_X1 U16 ( .B1(addr[3]), .B2(n16), .A(n7), .ZN(n3) );
  NAND3_X1 U17 ( .A1(n55), .A2(n53), .A3(n54), .ZN(n50) );
  OAI211_X1 U18 ( .C1(n33), .C2(n53), .A(n50), .B(n7), .ZN(n34) );
  NAND3_X1 U19 ( .A1(addr[2]), .A2(n53), .A3(n55), .ZN(n15) );
  NAND3_X1 U20 ( .A1(addr[0]), .A2(n53), .A3(n54), .ZN(n14) );
  INV_X1 U21 ( .A(n14), .ZN(n4) );
  INV_X1 U22 ( .A(addr[1]), .ZN(n11) );
  AOI21_X1 U23 ( .B1(z[1]), .B2(addr[3]), .A(n2), .ZN(n5) );
  NAND3_X1 U24 ( .A1(n15), .A2(n7), .A3(n5), .ZN(n35) );
  AOI21_X1 U25 ( .B1(n17), .B2(n1), .A(n2), .ZN(n6) );
  OAI221_X1 U26 ( .B1(addr[2]), .B2(n7), .C1(n32), .C2(n53), .A(n6), .ZN(n36)
         );
  NAND2_X1 U27 ( .A1(n1), .A2(addr[2]), .ZN(n51) );
  INV_X1 U28 ( .A(n51), .ZN(n9) );
  INV_X1 U29 ( .A(n15), .ZN(n8) );
  NOR2_X1 U30 ( .A1(n9), .A2(n8), .ZN(n10) );
  OAI211_X1 U31 ( .C1(n31), .C2(n53), .A(n14), .B(n10), .ZN(n37) );
  NAND2_X1 U32 ( .A1(n11), .A2(n16), .ZN(n12) );
  MUX2_X1 U33 ( .A(n12), .B(n30), .S(addr[3]), .Z(n13) );
  INV_X1 U34 ( .A(n13), .ZN(n38) );
  OAI221_X1 U35 ( .B1(addr[1]), .B2(n15), .C1(n29), .C2(n53), .A(n14), .ZN(n39) );
  MUX2_X1 U36 ( .A(n16), .B(n28), .S(addr[3]), .Z(n18) );
  NAND3_X1 U37 ( .A1(n51), .A2(n50), .A3(n18), .ZN(n40) );
  OAI21_X1 U38 ( .B1(n27), .B2(n53), .A(n52), .ZN(n41) );
  OAI21_X1 U39 ( .B1(n26), .B2(n53), .A(n52), .ZN(n42) );
  OAI21_X1 U40 ( .B1(n25), .B2(n53), .A(n52), .ZN(n43) );
  OAI21_X1 U41 ( .B1(n24), .B2(n53), .A(n52), .ZN(n44) );
  OAI21_X1 U42 ( .B1(n23), .B2(n53), .A(n52), .ZN(n45) );
endmodule


module layer2_12_8_12_16_B_rom_5 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b0;
  assign z[14] = 1'b0;
  assign z[13] = 1'b0;
  assign z[12] = 1'b0;
  assign z[11] = 1'b0;
  assign z[10] = 1'b0;
  assign z[9] = 1'b0;
  assign z[8] = 1'b0;
  assign z[7] = 1'b0;
  assign z[6] = 1'b0;
  assign z[5] = 1'b0;
  assign z[4] = 1'b1;
  assign z[3] = 1'b0;
  assign z[2] = 1'b1;
  assign z[1] = 1'b0;
  assign z[0] = 1'b1;

endmodule


module layer2_12_8_12_16_W_rom_6 ( clk, addr, z );
  input [3:0] addr;
  output [15:0] z;
  input clk;
  wire   n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n45, n46, n47, n48, n49, n50, n51, n52;

  DFF_X1 \z_reg[15]  ( .D(n44), .CK(clk), .Q(z[15]), .QN(n13) );
  DFF_X1 \z_reg[14]  ( .D(n43), .CK(clk), .Q(z[14]), .QN(n14) );
  DFF_X1 \z_reg[13]  ( .D(n42), .CK(clk), .Q(z[13]), .QN(n15) );
  DFF_X1 \z_reg[12]  ( .D(n41), .CK(clk), .Q(z[12]), .QN(n16) );
  DFF_X1 \z_reg[11]  ( .D(n40), .CK(clk), .Q(z[11]), .QN(n17) );
  DFF_X1 \z_reg[10]  ( .D(n39), .CK(clk), .Q(z[10]), .QN(n18) );
  DFF_X1 \z_reg[9]  ( .D(n38), .CK(clk), .Q(z[9]), .QN(n19) );
  DFF_X1 \z_reg[8]  ( .D(n37), .CK(clk), .Q(z[8]), .QN(n20) );
  DFF_X1 \z_reg[7]  ( .D(n36), .CK(clk), .Q(z[7]), .QN(n21) );
  DFF_X1 \z_reg[6]  ( .D(n35), .CK(clk), .Q(z[6]), .QN(n22) );
  DFF_X1 \z_reg[5]  ( .D(n34), .CK(clk), .Q(z[5]), .QN(n23) );
  DFF_X1 \z_reg[4]  ( .D(n33), .CK(clk), .Q(z[4]), .QN(n24) );
  DFF_X1 \z_reg[3]  ( .D(n32), .CK(clk), .Q(z[3]), .QN(n25) );
  DFF_X1 \z_reg[2]  ( .D(n31), .CK(clk), .Q(z[2]), .QN(n26) );
  DFF_X1 \z_reg[1]  ( .D(n30), .CK(clk), .Q(z[1]), .QN(n27) );
  DFF_X1 \z_reg[0]  ( .D(n29), .CK(clk), .Q(z[0]), .QN(n28) );
  OAI21_X1 U3 ( .B1(n52), .B2(n16), .A(n51), .ZN(n41) );
  OAI21_X1 U4 ( .B1(n52), .B2(n15), .A(n51), .ZN(n42) );
  OAI21_X1 U5 ( .B1(n52), .B2(n14), .A(n51), .ZN(n43) );
  OAI21_X1 U6 ( .B1(n52), .B2(n13), .A(n51), .ZN(n44) );
  INV_X1 U7 ( .A(addr[3]), .ZN(n52) );
  NAND2_X1 U8 ( .A1(addr[2]), .A2(n52), .ZN(n48) );
  INV_X1 U9 ( .A(n48), .ZN(n1) );
  INV_X1 U10 ( .A(addr[1]), .ZN(n7) );
  NAND2_X1 U11 ( .A1(n1), .A2(n7), .ZN(n50) );
  INV_X1 U12 ( .A(addr[2]), .ZN(n2) );
  NAND2_X1 U13 ( .A1(n52), .A2(n2), .ZN(n5) );
  MUX2_X1 U14 ( .A(n50), .B(n5), .S(addr[0]), .Z(n51) );
  XOR2_X1 U15 ( .A(n2), .B(addr[1]), .Z(n10) );
  INV_X1 U16 ( .A(n10), .ZN(n3) );
  MUX2_X1 U17 ( .A(n3), .B(n28), .S(addr[3]), .Z(n4) );
  OAI21_X1 U18 ( .B1(addr[0]), .B2(n5), .A(n4), .ZN(n29) );
  NAND2_X1 U19 ( .A1(addr[0]), .A2(n7), .ZN(n6) );
  INV_X1 U20 ( .A(n6), .ZN(n45) );
  OAI22_X1 U21 ( .A1(n45), .A2(n5), .B1(n27), .B2(n52), .ZN(n30) );
  OAI21_X1 U22 ( .B1(addr[0]), .B2(n7), .A(n6), .ZN(n8) );
  MUX2_X1 U23 ( .A(n8), .B(n26), .S(addr[3]), .Z(n9) );
  INV_X1 U24 ( .A(n9), .ZN(n31) );
  NOR2_X1 U25 ( .A1(addr[0]), .A2(n10), .ZN(n11) );
  MUX2_X1 U26 ( .A(n11), .B(n25), .S(addr[3]), .Z(n12) );
  INV_X1 U27 ( .A(n12), .ZN(n32) );
  MUX2_X1 U28 ( .A(n45), .B(n24), .S(addr[3]), .Z(n46) );
  NAND2_X1 U29 ( .A1(n48), .A2(n46), .ZN(n33) );
  MUX2_X1 U30 ( .A(addr[1]), .B(n23), .S(addr[3]), .Z(n47) );
  NAND2_X1 U31 ( .A1(n48), .A2(n47), .ZN(n34) );
  MUX2_X1 U32 ( .A(addr[0]), .B(n22), .S(addr[3]), .Z(n49) );
  NAND2_X1 U33 ( .A1(n50), .A2(n49), .ZN(n35) );
  OAI21_X1 U34 ( .B1(n21), .B2(n52), .A(n51), .ZN(n36) );
  OAI21_X1 U35 ( .B1(n20), .B2(n52), .A(n51), .ZN(n37) );
  OAI21_X1 U36 ( .B1(n19), .B2(n52), .A(n51), .ZN(n38) );
  OAI21_X1 U37 ( .B1(n18), .B2(n52), .A(n51), .ZN(n39) );
  OAI21_X1 U38 ( .B1(n17), .B2(n52), .A(n51), .ZN(n40) );
endmodule


module layer2_12_8_12_16_B_rom_6 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b1;
  assign z[14] = 1'b1;
  assign z[13] = 1'b1;
  assign z[12] = 1'b1;
  assign z[11] = 1'b1;
  assign z[10] = 1'b1;
  assign z[9] = 1'b1;
  assign z[8] = 1'b1;
  assign z[7] = 1'b1;
  assign z[6] = 1'b0;
  assign z[5] = 1'b0;
  assign z[4] = 1'b0;
  assign z[3] = 1'b1;
  assign z[2] = 1'b0;
  assign z[1] = 1'b1;
  assign z[0] = 1'b1;

endmodule


module layer2_12_8_12_16_W_rom_7 ( clk, addr, z );
  input [3:0] addr;
  output [15:0] z;
  input clk;
  wire   n7, n8, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n1, n2, n3, n4, n5, n6, n9,
         n10, n11, n12, n47, n48, n49, n50, n51, n52, n53;

  DFF_X1 \z_reg[14]  ( .D(n45), .CK(clk), .Q(z[14]), .QN(n16) );
  DFF_X1 \z_reg[13]  ( .D(n44), .CK(clk), .Q(z[13]), .QN(n17) );
  DFF_X1 \z_reg[12]  ( .D(n43), .CK(clk), .Q(z[12]), .QN(n18) );
  DFF_X1 \z_reg[11]  ( .D(n42), .CK(clk), .Q(z[11]), .QN(n19) );
  DFF_X1 \z_reg[10]  ( .D(n41), .CK(clk), .Q(z[10]), .QN(n20) );
  DFF_X1 \z_reg[9]  ( .D(n40), .CK(clk), .Q(z[9]), .QN(n21) );
  DFF_X1 \z_reg[8]  ( .D(n39), .CK(clk), .Q(z[8]), .QN(n22) );
  DFF_X1 \z_reg[7]  ( .D(n38), .CK(clk), .Q(z[7]), .QN(n23) );
  DFF_X1 \z_reg[6]  ( .D(n37), .CK(clk), .Q(z[6]), .QN(n24) );
  DFF_X1 \z_reg[5]  ( .D(n36), .CK(clk), .Q(z[5]), .QN(n25) );
  DFF_X1 \z_reg[4]  ( .D(n35), .CK(clk), .Q(z[4]), .QN(n26) );
  DFF_X1 \z_reg[3]  ( .D(n34), .CK(clk), .Q(z[3]), .QN(n27) );
  DFF_X1 \z_reg[2]  ( .D(n33), .CK(clk), .Q(z[2]), .QN(n28) );
  DFF_X1 \z_reg[1]  ( .D(n32), .CK(clk), .Q(z[1]), .QN(n29) );
  DFF_X1 \z_reg[0]  ( .D(n31), .CK(clk), .Q(z[0]), .QN(n30) );
  DFF_X1 \z_reg[15]  ( .D(n46), .CK(clk), .Q(z[15]), .QN(n15) );
  AND2_X1 U3 ( .A1(n53), .A2(n51), .ZN(n1) );
  NOR3_X1 U4 ( .A1(n52), .A2(n53), .A3(n51), .ZN(n7) );
  OAI21_X1 U5 ( .B1(n50), .B2(n18), .A(n14), .ZN(n43) );
  OAI21_X1 U6 ( .B1(n50), .B2(n17), .A(n14), .ZN(n44) );
  OAI21_X1 U7 ( .B1(n50), .B2(n16), .A(n14), .ZN(n45) );
  OAI21_X1 U8 ( .B1(n50), .B2(n15), .A(n14), .ZN(n46) );
  NOR2_X1 U9 ( .A1(addr[1]), .A2(n53), .ZN(n13) );
  NOR3_X1 U10 ( .A1(n53), .A2(addr[2]), .A3(addr[1]), .ZN(n8) );
  INV_X1 U11 ( .A(addr[1]), .ZN(n52) );
  INV_X1 U12 ( .A(addr[0]), .ZN(n53) );
  INV_X1 U13 ( .A(addr[2]), .ZN(n51) );
  INV_X1 U14 ( .A(addr[3]), .ZN(n50) );
  OAI21_X1 U15 ( .B1(n7), .B2(n1), .A(n50), .ZN(n14) );
  OAI211_X1 U16 ( .C1(addr[0]), .C2(addr[1]), .A(n51), .B(n50), .ZN(n3) );
  NAND2_X1 U17 ( .A1(addr[1]), .A2(addr[0]), .ZN(n9) );
  MUX2_X1 U18 ( .A(n9), .B(n30), .S(addr[3]), .Z(n2) );
  NAND2_X1 U19 ( .A1(n3), .A2(n2), .ZN(n31) );
  OAI21_X1 U20 ( .B1(n29), .B2(n50), .A(n3), .ZN(n32) );
  AOI211_X1 U21 ( .C1(n1), .C2(addr[1]), .A(n8), .B(n7), .ZN(n4) );
  MUX2_X1 U22 ( .A(n4), .B(n28), .S(addr[3]), .Z(n5) );
  INV_X1 U23 ( .A(n5), .ZN(n33) );
  MUX2_X1 U24 ( .A(addr[2]), .B(n27), .S(addr[3]), .Z(n6) );
  INV_X1 U25 ( .A(n6), .ZN(n34) );
  NOR2_X1 U26 ( .A1(addr[2]), .A2(n9), .ZN(n10) );
  MUX2_X1 U27 ( .A(n10), .B(n26), .S(addr[3]), .Z(n11) );
  INV_X1 U28 ( .A(n11), .ZN(n35) );
  MUX2_X1 U29 ( .A(addr[1]), .B(n13), .S(addr[2]), .Z(n12) );
  NOR2_X1 U30 ( .A1(n1), .A2(n12), .ZN(n47) );
  MUX2_X1 U31 ( .A(n47), .B(n25), .S(addr[3]), .Z(n48) );
  INV_X1 U32 ( .A(n48), .ZN(n36) );
  MUX2_X1 U33 ( .A(n1), .B(n24), .S(addr[3]), .Z(n49) );
  INV_X1 U34 ( .A(n49), .ZN(n37) );
  OAI21_X1 U35 ( .B1(n23), .B2(n50), .A(n14), .ZN(n38) );
  OAI21_X1 U36 ( .B1(n22), .B2(n50), .A(n14), .ZN(n39) );
  OAI21_X1 U37 ( .B1(n21), .B2(n50), .A(n14), .ZN(n40) );
  OAI21_X1 U38 ( .B1(n20), .B2(n50), .A(n14), .ZN(n41) );
  OAI21_X1 U39 ( .B1(n19), .B2(n50), .A(n14), .ZN(n42) );
endmodule


module layer2_12_8_12_16_B_rom_7 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b0;
  assign z[14] = 1'b0;
  assign z[13] = 1'b0;
  assign z[12] = 1'b0;
  assign z[11] = 1'b0;
  assign z[10] = 1'b0;
  assign z[9] = 1'b0;
  assign z[8] = 1'b0;
  assign z[7] = 1'b0;
  assign z[6] = 1'b1;
  assign z[5] = 1'b1;
  assign z[4] = 1'b1;
  assign z[3] = 1'b0;
  assign z[2] = 1'b1;
  assign z[1] = 1'b0;
  assign z[0] = 1'b1;

endmodule


module layer2_12_8_12_16_W_rom_8 ( clk, addr, z );
  input [3:0] addr;
  output [15:0] z;
  input clk;
  wire   n13, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n14, n47, n48, n49, n50, n51, n52;

  DFF_X1 \z_reg[15]  ( .D(n46), .CK(clk), .Q(z[15]), .QN(n16) );
  DFF_X1 \z_reg[14]  ( .D(n45), .CK(clk), .Q(z[14]), .QN(n17) );
  DFF_X1 \z_reg[13]  ( .D(n44), .CK(clk), .Q(z[13]), .QN(n18) );
  DFF_X1 \z_reg[12]  ( .D(n43), .CK(clk), .Q(z[12]), .QN(n19) );
  DFF_X1 \z_reg[11]  ( .D(n42), .CK(clk), .Q(z[11]), .QN(n20) );
  DFF_X1 \z_reg[10]  ( .D(n41), .CK(clk), .Q(z[10]), .QN(n21) );
  DFF_X1 \z_reg[9]  ( .D(n40), .CK(clk), .Q(z[9]), .QN(n22) );
  DFF_X1 \z_reg[8]  ( .D(n39), .CK(clk), .Q(z[8]), .QN(n23) );
  DFF_X1 \z_reg[7]  ( .D(n38), .CK(clk), .Q(z[7]), .QN(n24) );
  DFF_X1 \z_reg[6]  ( .D(n37), .CK(clk), .Q(z[6]), .QN(n25) );
  DFF_X1 \z_reg[5]  ( .D(n36), .CK(clk), .Q(z[5]), .QN(n26) );
  DFF_X1 \z_reg[4]  ( .D(n35), .CK(clk), .Q(z[4]), .QN(n27) );
  DFF_X1 \z_reg[3]  ( .D(n34), .CK(clk), .Q(z[3]), .QN(n28) );
  DFF_X1 \z_reg[2]  ( .D(n33), .CK(clk), .Q(z[2]), .QN(n29) );
  DFF_X1 \z_reg[1]  ( .D(n32), .CK(clk), .Q(z[1]), .QN(n30) );
  DFF_X1 \z_reg[0]  ( .D(n31), .CK(clk), .Q(z[0]) );
  NAND3_X1 U30 ( .A1(n52), .A2(n51), .A3(addr[2]), .ZN(n15) );
  INV_X1 U3 ( .A(addr[3]), .ZN(n50) );
  OAI21_X1 U4 ( .B1(n50), .B2(n19), .A(n13), .ZN(n43) );
  OAI21_X1 U5 ( .B1(n50), .B2(n18), .A(n13), .ZN(n44) );
  OAI21_X1 U6 ( .B1(n50), .B2(n17), .A(n13), .ZN(n45) );
  OAI21_X1 U7 ( .B1(n50), .B2(n16), .A(n13), .ZN(n46) );
  INV_X1 U8 ( .A(addr[2]), .ZN(n4) );
  OAI21_X1 U9 ( .B1(addr[1]), .B2(n4), .A(addr[0]), .ZN(n1) );
  AOI21_X1 U10 ( .B1(n15), .B2(n1), .A(addr[3]), .ZN(n2) );
  INV_X1 U11 ( .A(n2), .ZN(n13) );
  NAND2_X1 U12 ( .A1(addr[2]), .A2(n50), .ZN(n12) );
  INV_X1 U13 ( .A(n12), .ZN(n3) );
  INV_X1 U14 ( .A(addr[1]), .ZN(n51) );
  NAND2_X1 U15 ( .A1(n3), .A2(n51), .ZN(n11) );
  INV_X1 U16 ( .A(addr[0]), .ZN(n52) );
  NAND3_X1 U17 ( .A1(n51), .A2(n52), .A3(n50), .ZN(n48) );
  NAND2_X1 U18 ( .A1(addr[0]), .A2(addr[1]), .ZN(n14) );
  INV_X1 U19 ( .A(n14), .ZN(n6) );
  NAND2_X1 U20 ( .A1(n50), .A2(n4), .ZN(n49) );
  INV_X1 U21 ( .A(n49), .ZN(n5) );
  NAND2_X1 U22 ( .A1(n6), .A2(n5), .ZN(n10) );
  INV_X1 U23 ( .A(n10), .ZN(n7) );
  AOI21_X1 U24 ( .B1(z[0]), .B2(addr[3]), .A(n7), .ZN(n8) );
  NAND3_X1 U25 ( .A1(n11), .A2(n48), .A3(n8), .ZN(n31) );
  MUX2_X1 U26 ( .A(addr[0]), .B(n30), .S(addr[3]), .Z(n9) );
  OAI21_X1 U27 ( .B1(addr[1]), .B2(n49), .A(n9), .ZN(n32) );
  OAI222_X1 U28 ( .A1(n51), .A2(n49), .B1(n52), .B2(n12), .C1(n29), .C2(n50), 
        .ZN(n33) );
  OAI221_X1 U29 ( .B1(n52), .B2(n11), .C1(n28), .C2(n50), .A(n10), .ZN(n34) );
  OAI221_X1 U31 ( .B1(addr[0]), .B2(n12), .C1(n27), .C2(n50), .A(n48), .ZN(n35) );
  OAI221_X1 U32 ( .B1(addr[0]), .B2(n49), .C1(n26), .C2(n50), .A(n48), .ZN(n36) );
  MUX2_X1 U33 ( .A(n14), .B(n25), .S(addr[3]), .Z(n47) );
  NAND3_X1 U34 ( .A1(n49), .A2(n48), .A3(n47), .ZN(n37) );
  OAI21_X1 U35 ( .B1(n24), .B2(n50), .A(n13), .ZN(n38) );
  OAI21_X1 U36 ( .B1(n23), .B2(n50), .A(n13), .ZN(n39) );
  OAI21_X1 U37 ( .B1(n22), .B2(n50), .A(n13), .ZN(n40) );
  OAI21_X1 U38 ( .B1(n21), .B2(n50), .A(n13), .ZN(n41) );
  OAI21_X1 U39 ( .B1(n20), .B2(n50), .A(n13), .ZN(n42) );
endmodule


module layer2_12_8_12_16_B_rom_8 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b1;
  assign z[14] = 1'b1;
  assign z[13] = 1'b1;
  assign z[12] = 1'b1;
  assign z[11] = 1'b1;
  assign z[10] = 1'b1;
  assign z[9] = 1'b1;
  assign z[8] = 1'b1;
  assign z[7] = 1'b1;
  assign z[6] = 1'b1;
  assign z[5] = 1'b1;
  assign z[4] = 1'b0;
  assign z[3] = 1'b1;
  assign z[2] = 1'b1;
  assign z[1] = 1'b1;
  assign z[0] = 1'b1;

endmodule


module layer2_12_8_12_16_W_rom_9 ( clk, addr, z );
  input [3:0] addr;
  output [15:0] z;
  input clk;
  wire   n10, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n12, n13, n48, n49, n50, n51, n52, n53;

  DFF_X1 \z_reg[14]  ( .D(n46), .CK(clk), .Q(z[14]), .QN(n17) );
  DFF_X1 \z_reg[13]  ( .D(n45), .CK(clk), .Q(z[13]), .QN(n18) );
  DFF_X1 \z_reg[12]  ( .D(n44), .CK(clk), .Q(z[12]), .QN(n19) );
  DFF_X1 \z_reg[11]  ( .D(n43), .CK(clk), .Q(z[11]), .QN(n20) );
  DFF_X1 \z_reg[10]  ( .D(n42), .CK(clk), .Q(z[10]), .QN(n21) );
  DFF_X1 \z_reg[9]  ( .D(n41), .CK(clk), .Q(z[9]), .QN(n22) );
  DFF_X1 \z_reg[8]  ( .D(n40), .CK(clk), .Q(z[8]), .QN(n23) );
  DFF_X1 \z_reg[7]  ( .D(n39), .CK(clk), .Q(z[7]), .QN(n24) );
  DFF_X1 \z_reg[6]  ( .D(n38), .CK(clk), .Q(z[6]), .QN(n25) );
  DFF_X1 \z_reg[5]  ( .D(n37), .CK(clk), .Q(z[5]), .QN(n26) );
  DFF_X1 \z_reg[4]  ( .D(n36), .CK(clk), .Q(z[4]), .QN(n27) );
  DFF_X1 \z_reg[3]  ( .D(n35), .CK(clk), .Q(z[3]), .QN(n28) );
  DFF_X1 \z_reg[2]  ( .D(n34), .CK(clk), .Q(z[2]), .QN(n29) );
  DFF_X1 \z_reg[1]  ( .D(n33), .CK(clk), .Q(z[1]), .QN(n30) );
  DFF_X1 \z_reg[0]  ( .D(n32), .CK(clk), .Q(z[0]), .QN(n31) );
  XOR2_X1 U9 ( .A(n11), .B(addr[2]), .Z(n10) );
  XOR2_X1 U31 ( .A(n53), .B(addr[1]), .Z(n15) );
  DFF_X1 \z_reg[15]  ( .D(n47), .CK(clk), .Q(z[15]), .QN(n16) );
  AND2_X1 U3 ( .A1(addr[0]), .A2(n5), .ZN(n1) );
  INV_X1 U4 ( .A(addr[3]), .ZN(n52) );
  OAI21_X1 U5 ( .B1(n52), .B2(n19), .A(n14), .ZN(n44) );
  OAI21_X1 U6 ( .B1(n52), .B2(n18), .A(n14), .ZN(n45) );
  OAI21_X1 U7 ( .B1(n52), .B2(n17), .A(n14), .ZN(n46) );
  OAI21_X1 U8 ( .B1(n52), .B2(n16), .A(n14), .ZN(n47) );
  NAND2_X1 U10 ( .A1(addr[1]), .A2(addr[0]), .ZN(n11) );
  OAI21_X1 U11 ( .B1(n15), .B2(addr[2]), .A(n52), .ZN(n14) );
  INV_X1 U12 ( .A(addr[1]), .ZN(n5) );
  NAND3_X1 U13 ( .A1(addr[2]), .A2(n52), .A3(n1), .ZN(n13) );
  OAI21_X1 U14 ( .B1(n31), .B2(n52), .A(n13), .ZN(n32) );
  NOR2_X1 U15 ( .A1(addr[0]), .A2(addr[2]), .ZN(n2) );
  MUX2_X1 U16 ( .A(n2), .B(n30), .S(addr[3]), .Z(n3) );
  INV_X1 U17 ( .A(n3), .ZN(n33) );
  INV_X1 U18 ( .A(addr[2]), .ZN(n4) );
  NAND2_X1 U19 ( .A1(n52), .A2(n4), .ZN(n50) );
  OAI221_X1 U20 ( .B1(n1), .B2(n50), .C1(n29), .C2(n52), .A(n13), .ZN(n34) );
  INV_X1 U21 ( .A(addr[0]), .ZN(n53) );
  AOI21_X1 U22 ( .B1(n5), .B2(n53), .A(n10), .ZN(n6) );
  MUX2_X1 U23 ( .A(n6), .B(n28), .S(addr[3]), .Z(n7) );
  INV_X1 U24 ( .A(n7), .ZN(n35) );
  NOR2_X1 U25 ( .A1(addr[2]), .A2(n1), .ZN(n8) );
  MUX2_X1 U26 ( .A(n8), .B(n27), .S(addr[3]), .Z(n9) );
  INV_X1 U27 ( .A(n9), .ZN(n36) );
  INV_X1 U28 ( .A(n50), .ZN(n12) );
  NAND3_X1 U29 ( .A1(addr[1]), .A2(n53), .A3(n12), .ZN(n48) );
  OAI211_X1 U30 ( .C1(n26), .C2(n52), .A(n48), .B(n13), .ZN(n37) );
  NAND2_X1 U32 ( .A1(n52), .A2(n53), .ZN(n49) );
  MUX2_X1 U33 ( .A(n50), .B(n49), .S(addr[1]), .Z(n51) );
  OAI21_X1 U34 ( .B1(n25), .B2(n52), .A(n51), .ZN(n38) );
  OAI21_X1 U35 ( .B1(n24), .B2(n52), .A(n14), .ZN(n39) );
  OAI21_X1 U36 ( .B1(n23), .B2(n52), .A(n14), .ZN(n40) );
  OAI21_X1 U37 ( .B1(n22), .B2(n52), .A(n14), .ZN(n41) );
  OAI21_X1 U38 ( .B1(n21), .B2(n52), .A(n14), .ZN(n42) );
  OAI21_X1 U39 ( .B1(n20), .B2(n52), .A(n14), .ZN(n43) );
endmodule


module layer2_12_8_12_16_B_rom_9 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b0;
  assign z[14] = 1'b0;
  assign z[13] = 1'b0;
  assign z[12] = 1'b0;
  assign z[11] = 1'b0;
  assign z[10] = 1'b0;
  assign z[9] = 1'b0;
  assign z[8] = 1'b0;
  assign z[7] = 1'b0;
  assign z[6] = 1'b1;
  assign z[5] = 1'b1;
  assign z[4] = 1'b1;
  assign z[3] = 1'b0;
  assign z[2] = 1'b1;
  assign z[1] = 1'b1;
  assign z[0] = 1'b1;

endmodule


module layer2_12_8_12_16_W_rom_10 ( clk, addr, z );
  input [3:0] addr;
  output [15:0] z;
  input clk;
  wire   n8, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n1, n2, n3, n4, n5, n6, n7, n9, n10,
         n11, n45, n46, n47, n48;

  DFF_X1 \z_reg[15]  ( .D(n44), .CK(clk), .Q(z[15]), .QN(n14) );
  DFF_X1 \z_reg[14]  ( .D(n43), .CK(clk), .Q(z[14]), .QN(n15) );
  DFF_X1 \z_reg[13]  ( .D(n42), .CK(clk), .Q(z[13]), .QN(n16) );
  DFF_X1 \z_reg[12]  ( .D(n41), .CK(clk), .Q(z[12]), .QN(n17) );
  DFF_X1 \z_reg[11]  ( .D(n40), .CK(clk), .Q(z[11]), .QN(n18) );
  DFF_X1 \z_reg[10]  ( .D(n39), .CK(clk), .Q(z[10]), .QN(n19) );
  DFF_X1 \z_reg[9]  ( .D(n38), .CK(clk), .Q(z[9]), .QN(n20) );
  DFF_X1 \z_reg[8]  ( .D(n37), .CK(clk), .Q(z[8]), .QN(n21) );
  DFF_X1 \z_reg[7]  ( .D(n36), .CK(clk), .Q(z[7]), .QN(n22) );
  DFF_X1 \z_reg[6]  ( .D(n35), .CK(clk), .Q(z[6]), .QN(n23) );
  DFF_X1 \z_reg[5]  ( .D(n34), .CK(clk), .Q(z[5]), .QN(n24) );
  DFF_X1 \z_reg[4]  ( .D(n33), .CK(clk), .Q(z[4]), .QN(n25) );
  DFF_X1 \z_reg[3]  ( .D(n32), .CK(clk), .Q(z[3]), .QN(n26) );
  DFF_X1 \z_reg[2]  ( .D(n31), .CK(clk), .Q(z[2]), .QN(n1) );
  DFF_X1 \z_reg[1]  ( .D(n30), .CK(clk), .Q(z[1]), .QN(n27) );
  DFF_X1 \z_reg[0]  ( .D(n29), .CK(clk), .Q(z[0]), .QN(n28) );
  XOR2_X1 U29 ( .A(n48), .B(addr[2]), .Z(n13) );
  INV_X1 U3 ( .A(addr[3]), .ZN(n47) );
  NOR2_X1 U4 ( .A1(n48), .A2(addr[3]), .ZN(n8) );
  OAI21_X1 U5 ( .B1(n47), .B2(n17), .A(n12), .ZN(n41) );
  OAI21_X1 U6 ( .B1(n47), .B2(n16), .A(n12), .ZN(n42) );
  OAI21_X1 U7 ( .B1(n47), .B2(n15), .A(n12), .ZN(n43) );
  OAI21_X1 U8 ( .B1(n47), .B2(n14), .A(n12), .ZN(n44) );
  INV_X1 U9 ( .A(addr[1]), .ZN(n7) );
  OAI21_X1 U10 ( .B1(n13), .B2(n7), .A(n47), .ZN(n12) );
  INV_X1 U11 ( .A(addr[0]), .ZN(n48) );
  NAND2_X1 U12 ( .A1(addr[2]), .A2(n47), .ZN(n10) );
  INV_X1 U13 ( .A(n10), .ZN(n3) );
  OAI21_X1 U14 ( .B1(n8), .B2(n3), .A(n7), .ZN(n2) );
  OAI21_X1 U15 ( .B1(n28), .B2(n47), .A(n2), .ZN(n29) );
  OAI22_X1 U16 ( .A1(n7), .A2(n10), .B1(n27), .B2(n47), .ZN(n30) );
  INV_X1 U17 ( .A(addr[2]), .ZN(n5) );
  OAI21_X1 U18 ( .B1(addr[1]), .B2(n5), .A(n8), .ZN(n4) );
  NAND3_X1 U19 ( .A1(n3), .A2(n48), .A3(n7), .ZN(n6) );
  OAI211_X1 U20 ( .C1(n47), .C2(n1), .A(n4), .B(n6), .ZN(n31) );
  NAND3_X1 U21 ( .A1(n47), .A2(n48), .A3(n5), .ZN(n45) );
  OAI221_X1 U22 ( .B1(n7), .B2(n45), .C1(n26), .C2(n47), .A(n6), .ZN(n32) );
  MUX2_X1 U23 ( .A(n7), .B(n25), .S(addr[3]), .Z(n9) );
  NAND2_X1 U24 ( .A1(n10), .A2(n9), .ZN(n33) );
  INV_X1 U25 ( .A(n8), .ZN(n11) );
  OAI221_X1 U26 ( .B1(addr[1]), .B2(n11), .C1(n24), .C2(n47), .A(n45), .ZN(n34) );
  MUX2_X1 U27 ( .A(n45), .B(n11), .S(addr[1]), .Z(n46) );
  OAI21_X1 U28 ( .B1(n23), .B2(n47), .A(n46), .ZN(n35) );
  OAI21_X1 U30 ( .B1(n22), .B2(n47), .A(n12), .ZN(n36) );
  OAI21_X1 U31 ( .B1(n21), .B2(n47), .A(n12), .ZN(n37) );
  OAI21_X1 U32 ( .B1(n20), .B2(n47), .A(n12), .ZN(n38) );
  OAI21_X1 U33 ( .B1(n19), .B2(n47), .A(n12), .ZN(n39) );
  OAI21_X1 U34 ( .B1(n18), .B2(n47), .A(n12), .ZN(n40) );
endmodule


module layer2_12_8_12_16_B_rom_10 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b0;
  assign z[14] = 1'b0;
  assign z[13] = 1'b0;
  assign z[12] = 1'b0;
  assign z[11] = 1'b0;
  assign z[10] = 1'b0;
  assign z[9] = 1'b0;
  assign z[8] = 1'b0;
  assign z[7] = 1'b0;
  assign z[6] = 1'b1;
  assign z[5] = 1'b1;
  assign z[4] = 1'b1;
  assign z[3] = 1'b1;
  assign z[2] = 1'b0;
  assign z[1] = 1'b1;
  assign z[0] = 1'b1;

endmodule


module layer2_12_8_12_16_W_rom_11 ( clk, addr, z );
  input [3:0] addr;
  output [15:0] z;
  input clk;
  wire   n7, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n1, n2, n3, n4, n5, n6, n8, n9, n10,
         n11, n45, n46, n47, n48, n49, n50;
  assign z[3] = 1'b0;

  DFF_X1 \z_reg[15]  ( .D(n44), .CK(clk), .Q(z[15]), .QN(n16) );
  DFF_X1 \z_reg[14]  ( .D(n43), .CK(clk), .Q(z[14]), .QN(n17) );
  DFF_X1 \z_reg[13]  ( .D(n42), .CK(clk), .Q(z[13]), .QN(n18) );
  DFF_X1 \z_reg[12]  ( .D(n41), .CK(clk), .Q(z[12]), .QN(n19) );
  DFF_X1 \z_reg[11]  ( .D(n40), .CK(clk), .Q(z[11]), .QN(n20) );
  DFF_X1 \z_reg[10]  ( .D(n39), .CK(clk), .Q(z[10]), .QN(n21) );
  DFF_X1 \z_reg[9]  ( .D(n38), .CK(clk), .Q(z[9]), .QN(n22) );
  DFF_X1 \z_reg[8]  ( .D(n37), .CK(clk), .Q(z[8]), .QN(n23) );
  DFF_X1 \z_reg[7]  ( .D(n36), .CK(clk), .Q(z[7]), .QN(n24) );
  DFF_X1 \z_reg[6]  ( .D(n35), .CK(clk), .Q(z[6]), .QN(n25) );
  DFF_X1 \z_reg[5]  ( .D(n34), .CK(clk), .Q(z[5]), .QN(n26) );
  DFF_X1 \z_reg[4]  ( .D(n33), .CK(clk), .Q(z[4]), .QN(n1) );
  DFF_X1 \z_reg[2]  ( .D(n32), .CK(clk), .Q(z[2]), .QN(n27) );
  DFF_X1 \z_reg[1]  ( .D(n31), .CK(clk), .Q(z[1]), .QN(n28) );
  DFF_X1 \z_reg[0]  ( .D(n30), .CK(clk), .Q(z[0]), .QN(n29) );
  XOR2_X1 U29 ( .A(n15), .B(addr[0]), .Z(n14) );
  NAND2_X1 U3 ( .A1(addr[2]), .A2(n50), .ZN(n15) );
  INV_X1 U4 ( .A(addr[3]), .ZN(n48) );
  NOR2_X1 U5 ( .A1(addr[1]), .A2(addr[0]), .ZN(n12) );
  OAI21_X1 U6 ( .B1(n48), .B2(n19), .A(n13), .ZN(n41) );
  OAI21_X1 U7 ( .B1(n48), .B2(n18), .A(n13), .ZN(n42) );
  OAI21_X1 U8 ( .B1(n48), .B2(n17), .A(n13), .ZN(n43) );
  OAI21_X1 U9 ( .B1(n48), .B2(n16), .A(n13), .ZN(n44) );
  NOR2_X1 U10 ( .A1(n49), .A2(addr[3]), .ZN(n7) );
  INV_X1 U11 ( .A(addr[1]), .ZN(n50) );
  NAND2_X1 U12 ( .A1(n14), .A2(n48), .ZN(n13) );
  INV_X1 U13 ( .A(addr[2]), .ZN(n49) );
  NAND2_X1 U14 ( .A1(n7), .A2(addr[1]), .ZN(n11) );
  XOR2_X1 U15 ( .A(n50), .B(addr[0]), .Z(n2) );
  MUX2_X1 U16 ( .A(n2), .B(n29), .S(addr[3]), .Z(n3) );
  NAND2_X1 U17 ( .A1(n11), .A2(n3), .ZN(n30) );
  INV_X1 U18 ( .A(n7), .ZN(n45) );
  INV_X1 U19 ( .A(n12), .ZN(n4) );
  OAI22_X1 U20 ( .A1(n45), .A2(n4), .B1(n28), .B2(n48), .ZN(n31) );
  OAI21_X1 U21 ( .B1(n27), .B2(n48), .A(n11), .ZN(n32) );
  INV_X1 U22 ( .A(addr[0]), .ZN(n8) );
  NAND2_X1 U23 ( .A1(n50), .A2(n49), .ZN(n5) );
  MUX2_X1 U24 ( .A(n5), .B(n1), .S(addr[3]), .Z(n6) );
  OAI211_X1 U25 ( .C1(n45), .C2(n8), .A(n11), .B(n6), .ZN(n33) );
  NAND2_X1 U26 ( .A1(addr[0]), .A2(addr[1]), .ZN(n9) );
  MUX2_X1 U27 ( .A(n9), .B(n26), .S(addr[3]), .Z(n10) );
  NAND2_X1 U28 ( .A1(n11), .A2(n10), .ZN(n34) );
  NAND2_X1 U30 ( .A1(n48), .A2(n49), .ZN(n46) );
  MUX2_X1 U31 ( .A(n46), .B(n45), .S(n12), .Z(n47) );
  OAI21_X1 U32 ( .B1(n25), .B2(n48), .A(n47), .ZN(n35) );
  OAI21_X1 U34 ( .B1(n24), .B2(n48), .A(n13), .ZN(n36) );
  OAI21_X1 U35 ( .B1(n23), .B2(n48), .A(n13), .ZN(n37) );
  OAI21_X1 U36 ( .B1(n22), .B2(n48), .A(n13), .ZN(n38) );
  OAI21_X1 U37 ( .B1(n21), .B2(n48), .A(n13), .ZN(n39) );
  OAI21_X1 U38 ( .B1(n20), .B2(n48), .A(n13), .ZN(n40) );
endmodule


module layer2_12_8_12_16_B_rom_11 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b0;
  assign z[14] = 1'b0;
  assign z[13] = 1'b0;
  assign z[12] = 1'b0;
  assign z[11] = 1'b0;
  assign z[10] = 1'b0;
  assign z[9] = 1'b0;
  assign z[8] = 1'b0;
  assign z[7] = 1'b0;
  assign z[6] = 1'b0;
  assign z[5] = 1'b0;
  assign z[4] = 1'b0;
  assign z[3] = 1'b1;
  assign z[2] = 1'b0;
  assign z[1] = 1'b0;
  assign z[0] = 1'b1;

endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_0_DW_mult_tc_1 ( a, b, 
        product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n9, n12, n13, n16, n18, n19, n21, n23, n25, n27, n29, n31,
         n32, n34, n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n50,
         n52, n53, n55, n56, n57, n58, n59, n62, n63, n64, n65, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n93, n95, n96, n97, n98, n99, n101,
         n103, n104, n105, n106, n107, n111, n112, n113, n114, n115, n117,
         n119, n120, n122, n125, n131, n135, n139, n141, n142, n143, n144,
         n145, n146, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n245, n247, n249, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n418,
         n419, n420, n421, n422, n423, n424, n426, n427, n428, n429, n433,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U148 ( .A(n265), .B(n144), .Z(n145) );
  XOR2_X1 U152 ( .A(n301), .B(n148), .Z(n149) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U162 ( .A(n170), .B(n172), .CI(n179), .CO(n165), .S(n166) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n263), .CI(n291), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n317), .B(n252), .CO(n173), .S(n174) );
  FA_X1 U167 ( .A(n180), .B(n187), .CI(n178), .CO(n175), .S(n176) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U169 ( .A(n193), .B(n282), .CI(n191), .CO(n179), .S(n180) );
  FA_X1 U170 ( .A(n268), .B(n274), .CI(n292), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U172 ( .A(n197), .B(n190), .CI(n188), .CO(n185), .S(n186) );
  FA_X1 U173 ( .A(n199), .B(n201), .CI(n192), .CO(n187), .S(n188) );
  FA_X1 U174 ( .A(n275), .B(n293), .CI(n194), .CO(n189), .S(n190) );
  FA_X1 U175 ( .A(n253), .B(n283), .CI(n305), .CO(n191), .S(n192) );
  HA_X1 U176 ( .A(n269), .B(n319), .CO(n193), .S(n194) );
  FA_X1 U177 ( .A(n205), .B(n200), .CI(n198), .CO(n195), .S(n196) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U179 ( .A(n276), .B(n284), .CI(n294), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n320), .B(n270), .CI(n306), .CO(n201), .S(n202) );
  FA_X1 U181 ( .A(n208), .B(n213), .CI(n206), .CO(n203), .S(n204) );
  FA_X1 U182 ( .A(n215), .B(n307), .CI(n210), .CO(n205), .S(n206) );
  FA_X1 U183 ( .A(n254), .B(n285), .CI(n295), .CO(n207), .S(n208) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U185 ( .A(n216), .B(n219), .CI(n214), .CO(n211), .S(n212) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n322), .B(n278), .CI(n308), .CO(n215), .S(n216) );
  FA_X1 U188 ( .A(n225), .B(n222), .CI(n220), .CO(n217), .S(n218) );
  FA_X1 U189 ( .A(n255), .B(n309), .CI(n297), .CO(n219), .S(n220) );
  HA_X1 U190 ( .A(n287), .B(n323), .CO(n221), .S(n222) );
  FA_X1 U192 ( .A(n324), .B(n288), .CI(n310), .CO(n225), .S(n226) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  HA_X1 U194 ( .A(n311), .B(n325), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n326), .B(n312), .CI(n300), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  CLKBUF_X1 U414 ( .A(n1), .Z(n490) );
  NAND2_X1 U415 ( .A1(n556), .A2(n9), .ZN(n491) );
  XNOR2_X1 U416 ( .A(n518), .B(n492), .ZN(product[7]) );
  AND2_X1 U417 ( .A1(n131), .A2(n98), .ZN(n492) );
  AOI21_X1 U418 ( .B1(n96), .B2(n558), .A(n93), .ZN(n493) );
  NOR2_X1 U419 ( .A1(n164), .A2(n175), .ZN(n75) );
  OR2_X1 U420 ( .A1(n186), .A2(n195), .ZN(n494) );
  OR2_X1 U421 ( .A1(n329), .A2(n258), .ZN(n495) );
  OR2_X1 U422 ( .A1(n232), .A2(n233), .ZN(n496) );
  OR2_X1 U423 ( .A1(n228), .A2(n231), .ZN(n497) );
  AND2_X1 U424 ( .A1(n232), .A2(n233), .ZN(n498) );
  BUF_X1 U425 ( .A(n546), .Z(n518) );
  AND2_X1 U426 ( .A1(n552), .A2(n553), .ZN(n499) );
  AND2_X1 U427 ( .A1(n553), .A2(n552), .ZN(n45) );
  NAND2_X1 U428 ( .A1(n555), .A2(n516), .ZN(n500) );
  NAND2_X1 U429 ( .A1(n555), .A2(n516), .ZN(n501) );
  NAND2_X1 U430 ( .A1(n555), .A2(n516), .ZN(n18) );
  NOR2_X1 U431 ( .A1(n186), .A2(n195), .ZN(n502) );
  NOR2_X1 U432 ( .A1(n186), .A2(n195), .ZN(n82) );
  CLKBUF_X1 U433 ( .A(n29), .Z(n503) );
  BUF_X1 U434 ( .A(n12), .Z(n531) );
  NAND2_X1 U435 ( .A1(n429), .A2(n27), .ZN(n29) );
  INV_X1 U436 ( .A(n32), .ZN(n504) );
  XNOR2_X1 U437 ( .A(n571), .B(n249), .ZN(n505) );
  XOR2_X1 U438 ( .A(n578), .B(a[6]), .Z(n526) );
  XNOR2_X1 U439 ( .A(n149), .B(n506), .ZN(n144) );
  XNOR2_X1 U440 ( .A(n271), .B(n146), .ZN(n506) );
  BUF_X2 U441 ( .A(n12), .Z(n532) );
  XNOR2_X1 U442 ( .A(n166), .B(n507), .ZN(n164) );
  XNOR2_X1 U443 ( .A(n177), .B(n168), .ZN(n507) );
  INV_X1 U444 ( .A(n515), .ZN(n37) );
  BUF_X1 U445 ( .A(n23), .Z(n512) );
  XNOR2_X1 U446 ( .A(n88), .B(n508), .ZN(product[10]) );
  NAND2_X1 U447 ( .A1(n530), .A2(n86), .ZN(n508) );
  CLKBUF_X1 U448 ( .A(n21), .Z(n509) );
  CLKBUF_X1 U449 ( .A(n1), .Z(n510) );
  BUF_X4 U450 ( .A(n9), .Z(n566) );
  CLKBUF_X1 U451 ( .A(n580), .Z(n511) );
  INV_X1 U452 ( .A(n574), .ZN(n573) );
  INV_X2 U453 ( .A(n574), .ZN(n572) );
  XOR2_X1 U454 ( .A(n511), .B(n424), .Z(n351) );
  XOR2_X1 U455 ( .A(n25), .B(a[10]), .Z(n529) );
  XNOR2_X1 U456 ( .A(n517), .B(a[4]), .ZN(n555) );
  INV_X1 U457 ( .A(n577), .ZN(n575) );
  INV_X1 U458 ( .A(n510), .ZN(n513) );
  INV_X1 U459 ( .A(n529), .ZN(n514) );
  XNOR2_X1 U460 ( .A(n582), .B(a[12]), .ZN(n515) );
  BUF_X1 U461 ( .A(n16), .Z(n516) );
  INV_X1 U462 ( .A(n13), .ZN(n517) );
  XNOR2_X1 U463 ( .A(n580), .B(a[8]), .ZN(n429) );
  OR2_X1 U464 ( .A1(n204), .A2(n211), .ZN(n519) );
  INV_X1 U465 ( .A(n529), .ZN(n32) );
  XOR2_X1 U466 ( .A(n578), .B(a[8]), .Z(n27) );
  XNOR2_X1 U467 ( .A(n582), .B(a[10]), .ZN(n428) );
  INV_X1 U468 ( .A(n582), .ZN(n581) );
  OAI21_X1 U469 ( .B1(n89), .B2(n91), .A(n90), .ZN(n520) );
  OR2_X1 U470 ( .A1(n176), .A2(n185), .ZN(n521) );
  BUF_X1 U471 ( .A(n97), .Z(n524) );
  INV_X1 U472 ( .A(n572), .ZN(n522) );
  CLKBUF_X1 U473 ( .A(n107), .Z(n523) );
  INV_X1 U474 ( .A(n571), .ZN(n525) );
  OR2_X2 U475 ( .A1(n526), .A2(n554), .ZN(n23) );
  CLKBUF_X3 U476 ( .A(n19), .Z(n544) );
  XNOR2_X1 U477 ( .A(n226), .B(n527), .ZN(n224) );
  XNOR2_X1 U478 ( .A(n229), .B(n298), .ZN(n527) );
  NAND2_X1 U479 ( .A1(n428), .A2(n32), .ZN(n528) );
  OR2_X1 U480 ( .A1(n196), .A2(n203), .ZN(n530) );
  NAND2_X1 U481 ( .A1(n556), .A2(n9), .ZN(n12) );
  NOR2_X1 U482 ( .A1(n196), .A2(n203), .ZN(n85) );
  BUF_X2 U483 ( .A(n27), .Z(n533) );
  XOR2_X1 U484 ( .A(n544), .B(a[8]), .Z(n534) );
  BUF_X1 U485 ( .A(n104), .Z(n535) );
  INV_X1 U486 ( .A(n554), .ZN(n21) );
  NAND2_X1 U487 ( .A1(n226), .A2(n229), .ZN(n536) );
  NAND2_X1 U488 ( .A1(n226), .A2(n298), .ZN(n537) );
  NAND2_X1 U489 ( .A1(n229), .A2(n298), .ZN(n538) );
  NAND3_X1 U490 ( .A1(n536), .A2(n537), .A3(n538), .ZN(n223) );
  XNOR2_X1 U491 ( .A(n45), .B(n539), .ZN(product[12]) );
  AND2_X1 U492 ( .A1(n521), .A2(n79), .ZN(n539) );
  NAND2_X1 U493 ( .A1(n166), .A2(n177), .ZN(n540) );
  NAND2_X1 U494 ( .A1(n166), .A2(n168), .ZN(n541) );
  NAND2_X1 U495 ( .A1(n177), .A2(n168), .ZN(n542) );
  NAND3_X1 U496 ( .A1(n540), .A2(n541), .A3(n542), .ZN(n163) );
  BUF_X2 U497 ( .A(n570), .Z(n543) );
  INV_X1 U498 ( .A(n249), .ZN(n570) );
  XNOR2_X1 U499 ( .A(n571), .B(n249), .ZN(n433) );
  OAI21_X1 U500 ( .B1(n546), .B2(n524), .A(n98), .ZN(n545) );
  AOI21_X1 U501 ( .B1(n535), .B2(n567), .A(n101), .ZN(n546) );
  CLKBUF_X1 U502 ( .A(n91), .Z(n547) );
  OR2_X1 U503 ( .A1(n550), .A2(n403), .ZN(n548) );
  OR2_X1 U504 ( .A1(n402), .A2(n570), .ZN(n549) );
  NAND2_X1 U505 ( .A1(n548), .A2(n549), .ZN(n324) );
  XOR2_X1 U506 ( .A(n574), .B(a[4]), .Z(n16) );
  XNOR2_X1 U507 ( .A(n574), .B(a[2]), .ZN(n556) );
  INV_X2 U508 ( .A(n580), .ZN(n579) );
  CLKBUF_X3 U509 ( .A(n16), .Z(n565) );
  NAND2_X1 U510 ( .A1(n433), .A2(n570), .ZN(n550) );
  NAND2_X1 U511 ( .A1(n505), .A2(n570), .ZN(n551) );
  NAND2_X1 U512 ( .A1(n520), .A2(n80), .ZN(n552) );
  INV_X1 U513 ( .A(n81), .ZN(n553) );
  XNOR2_X1 U514 ( .A(n577), .B(a[6]), .ZN(n554) );
  BUF_X1 U515 ( .A(n43), .Z(n568) );
  NAND2_X1 U516 ( .A1(n557), .A2(n69), .ZN(n47) );
  INV_X1 U517 ( .A(n73), .ZN(n71) );
  AOI21_X1 U518 ( .B1(n74), .B2(n557), .A(n67), .ZN(n65) );
  INV_X1 U519 ( .A(n69), .ZN(n67) );
  NAND2_X1 U520 ( .A1(n73), .A2(n557), .ZN(n64) );
  INV_X1 U521 ( .A(n74), .ZN(n72) );
  INV_X1 U522 ( .A(n95), .ZN(n93) );
  NAND2_X1 U523 ( .A1(n519), .A2(n90), .ZN(n52) );
  NAND2_X1 U524 ( .A1(n125), .A2(n76), .ZN(n48) );
  INV_X1 U525 ( .A(n75), .ZN(n125) );
  OR2_X1 U526 ( .A1(n152), .A2(n163), .ZN(n557) );
  OAI21_X1 U527 ( .B1(n75), .B2(n79), .A(n76), .ZN(n74) );
  NAND2_X1 U528 ( .A1(n494), .A2(n83), .ZN(n50) );
  NOR2_X1 U529 ( .A1(n75), .A2(n78), .ZN(n73) );
  NAND2_X1 U530 ( .A1(n152), .A2(n163), .ZN(n69) );
  NAND2_X1 U531 ( .A1(n558), .A2(n95), .ZN(n53) );
  INV_X1 U532 ( .A(n119), .ZN(n117) );
  AOI21_X1 U533 ( .B1(n104), .B2(n567), .A(n101), .ZN(n99) );
  OAI21_X1 U534 ( .B1(n113), .B2(n115), .A(n114), .ZN(n112) );
  NAND2_X1 U535 ( .A1(n497), .A2(n106), .ZN(n56) );
  NOR2_X1 U536 ( .A1(n176), .A2(n185), .ZN(n78) );
  XOR2_X1 U537 ( .A(n58), .B(n115), .Z(product[3]) );
  NAND2_X1 U538 ( .A1(n135), .A2(n114), .ZN(n58) );
  OAI21_X1 U539 ( .B1(n99), .B2(n97), .A(n98), .ZN(n96) );
  INV_X1 U540 ( .A(n524), .ZN(n131) );
  XNOR2_X1 U541 ( .A(n57), .B(n112), .ZN(product[4]) );
  NAND2_X1 U542 ( .A1(n496), .A2(n111), .ZN(n57) );
  NAND2_X1 U543 ( .A1(n176), .A2(n185), .ZN(n79) );
  NAND2_X1 U544 ( .A1(n164), .A2(n175), .ZN(n76) );
  NAND2_X1 U545 ( .A1(n196), .A2(n203), .ZN(n86) );
  NAND2_X1 U546 ( .A1(n212), .A2(n217), .ZN(n95) );
  OR2_X1 U547 ( .A1(n212), .A2(n217), .ZN(n558) );
  XNOR2_X1 U548 ( .A(n59), .B(n120), .ZN(product[2]) );
  NAND2_X1 U549 ( .A1(n560), .A2(n119), .ZN(n59) );
  OR2_X1 U550 ( .A1(n139), .A2(n151), .ZN(n559) );
  NOR2_X1 U551 ( .A1(n218), .A2(n223), .ZN(n97) );
  XNOR2_X1 U552 ( .A(n63), .B(n46), .ZN(product[15]) );
  NAND2_X1 U553 ( .A1(n559), .A2(n62), .ZN(n46) );
  NAND2_X1 U554 ( .A1(n328), .A2(n314), .ZN(n119) );
  NOR2_X1 U555 ( .A1(n228), .A2(n231), .ZN(n105) );
  NAND2_X1 U556 ( .A1(n218), .A2(n223), .ZN(n98) );
  NAND2_X1 U557 ( .A1(n228), .A2(n231), .ZN(n106) );
  OR2_X1 U558 ( .A1(n328), .A2(n314), .ZN(n560) );
  OR2_X1 U559 ( .A1(n232), .A2(n233), .ZN(n561) );
  NAND2_X1 U560 ( .A1(n232), .A2(n233), .ZN(n111) );
  INV_X1 U561 ( .A(n41), .ZN(n235) );
  OR2_X1 U562 ( .A1(n224), .A2(n227), .ZN(n567) );
  AND2_X1 U563 ( .A1(n495), .A2(n122), .ZN(product[1]) );
  NAND2_X1 U564 ( .A1(n505), .A2(n570), .ZN(n6) );
  OAI22_X1 U565 ( .A1(n550), .A2(n407), .B1(n406), .B2(n543), .ZN(n328) );
  XNOR2_X1 U566 ( .A(n583), .B(a[14]), .ZN(n41) );
  OR2_X1 U567 ( .A1(n568), .A2(n522), .ZN(n392) );
  OR2_X1 U568 ( .A1(n568), .A2(n517), .ZN(n377) );
  OAI22_X1 U569 ( .A1(n6), .A2(n400), .B1(n399), .B2(n543), .ZN(n321) );
  XNOR2_X1 U570 ( .A(n579), .B(n568), .ZN(n352) );
  OAI22_X1 U571 ( .A1(n6), .A2(n406), .B1(n405), .B2(n543), .ZN(n327) );
  AND2_X1 U572 ( .A1(n569), .A2(n515), .ZN(n264) );
  OAI22_X1 U573 ( .A1(n6), .A2(n397), .B1(n396), .B2(n543), .ZN(n318) );
  OAI22_X1 U574 ( .A1(n550), .A2(n408), .B1(n407), .B2(n543), .ZN(n329) );
  XNOR2_X1 U575 ( .A(n155), .B(n563), .ZN(n139) );
  XNOR2_X1 U576 ( .A(n153), .B(n141), .ZN(n563) );
  XNOR2_X1 U577 ( .A(n157), .B(n564), .ZN(n141) );
  XNOR2_X1 U578 ( .A(n145), .B(n143), .ZN(n564) );
  OAI22_X1 U579 ( .A1(n39), .A2(n336), .B1(n37), .B2(n335), .ZN(n263) );
  OAI22_X1 U580 ( .A1(n34), .A2(n342), .B1(n341), .B2(n514), .ZN(n268) );
  OAI22_X1 U581 ( .A1(n528), .A2(n341), .B1(n340), .B2(n514), .ZN(n267) );
  OAI22_X1 U582 ( .A1(n550), .A2(n396), .B1(n395), .B2(n543), .ZN(n317) );
  OAI22_X1 U583 ( .A1(n39), .A2(n584), .B1(n337), .B2(n37), .ZN(n252) );
  OR2_X1 U584 ( .A1(n568), .A2(n584), .ZN(n337) );
  OAI22_X1 U585 ( .A1(n551), .A2(n398), .B1(n397), .B2(n543), .ZN(n319) );
  OAI22_X1 U586 ( .A1(n528), .A2(n343), .B1(n342), .B2(n514), .ZN(n269) );
  XNOR2_X1 U587 ( .A(n581), .B(n568), .ZN(n343) );
  OAI22_X1 U588 ( .A1(n42), .A2(n586), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U589 ( .A1(n568), .A2(n586), .ZN(n332) );
  OAI22_X1 U590 ( .A1(n551), .A2(n404), .B1(n403), .B2(n570), .ZN(n325) );
  XOR2_X1 U591 ( .A(n315), .B(n261), .Z(n150) );
  OAI22_X1 U592 ( .A1(n6), .A2(n394), .B1(n393), .B2(n543), .ZN(n315) );
  AND2_X1 U593 ( .A1(n569), .A2(n245), .ZN(n300) );
  OAI22_X1 U594 ( .A1(n550), .A2(n405), .B1(n404), .B2(n570), .ZN(n326) );
  XNOR2_X1 U595 ( .A(n583), .B(n568), .ZN(n336) );
  NAND2_X1 U596 ( .A1(n428), .A2(n32), .ZN(n34) );
  NAND2_X1 U597 ( .A1(n427), .A2(n37), .ZN(n39) );
  XOR2_X1 U598 ( .A(n583), .B(a[12]), .Z(n427) );
  XNOR2_X1 U599 ( .A(n576), .B(n568), .ZN(n376) );
  AND2_X1 U600 ( .A1(n569), .A2(n534), .ZN(n278) );
  OAI22_X1 U601 ( .A1(n550), .A2(n401), .B1(n400), .B2(n543), .ZN(n322) );
  AND2_X1 U602 ( .A1(n569), .A2(n554), .ZN(n288) );
  AND2_X1 U603 ( .A1(n569), .A2(n504), .ZN(n270) );
  OAI22_X1 U604 ( .A1(n399), .A2(n551), .B1(n398), .B2(n543), .ZN(n320) );
  AND2_X1 U605 ( .A1(n569), .A2(n235), .ZN(n260) );
  OAI22_X1 U606 ( .A1(n551), .A2(n395), .B1(n394), .B2(n543), .ZN(n316) );
  OAI22_X1 U607 ( .A1(n39), .A2(n335), .B1(n37), .B2(n334), .ZN(n262) );
  INV_X1 U608 ( .A(n25), .ZN(n580) );
  OAI22_X1 U609 ( .A1(n34), .A2(n582), .B1(n344), .B2(n514), .ZN(n253) );
  OAI22_X1 U610 ( .A1(n34), .A2(n340), .B1(n339), .B2(n514), .ZN(n266) );
  NAND2_X1 U611 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U612 ( .A(n585), .B(a[14]), .Z(n426) );
  INV_X1 U613 ( .A(n13), .ZN(n577) );
  INV_X1 U614 ( .A(n7), .ZN(n574) );
  OAI22_X1 U615 ( .A1(n6), .A2(n402), .B1(n401), .B2(n543), .ZN(n323) );
  XNOR2_X1 U616 ( .A(n544), .B(n568), .ZN(n363) );
  AND2_X1 U617 ( .A1(n569), .A2(n247), .ZN(n314) );
  OR2_X1 U618 ( .A1(n568), .A2(n582), .ZN(n344) );
  AND2_X1 U619 ( .A1(n569), .A2(n249), .ZN(product[0]) );
  OR2_X1 U620 ( .A1(n568), .A2(n511), .ZN(n353) );
  OR2_X1 U621 ( .A1(n568), .A2(n578), .ZN(n364) );
  XNOR2_X1 U622 ( .A(n544), .B(b[9]), .ZN(n354) );
  OAI22_X1 U623 ( .A1(n39), .A2(n334), .B1(n37), .B2(n333), .ZN(n261) );
  XNOR2_X1 U624 ( .A(n583), .B(n422), .ZN(n333) );
  XNOR2_X1 U625 ( .A(n576), .B(b[11]), .ZN(n365) );
  XNOR2_X1 U626 ( .A(n581), .B(n424), .ZN(n342) );
  XNOR2_X1 U627 ( .A(n581), .B(n423), .ZN(n341) );
  XNOR2_X1 U628 ( .A(n581), .B(n422), .ZN(n340) );
  XNOR2_X1 U629 ( .A(n581), .B(n421), .ZN(n339) );
  XNOR2_X1 U630 ( .A(n583), .B(n423), .ZN(n334) );
  XNOR2_X1 U631 ( .A(n583), .B(n424), .ZN(n335) );
  OAI22_X1 U632 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U633 ( .A(n585), .B(n424), .ZN(n330) );
  XNOR2_X1 U634 ( .A(n585), .B(n568), .ZN(n331) );
  XNOR2_X1 U635 ( .A(n525), .B(b[11]), .ZN(n397) );
  XNOR2_X1 U636 ( .A(n525), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U637 ( .A(n490), .B(b[13]), .ZN(n395) );
  XNOR2_X1 U638 ( .A(n525), .B(b[14]), .ZN(n394) );
  XNOR2_X1 U639 ( .A(n579), .B(n418), .ZN(n345) );
  OAI22_X1 U640 ( .A1(n528), .A2(n339), .B1(n338), .B2(n514), .ZN(n265) );
  XNOR2_X1 U641 ( .A(n581), .B(n420), .ZN(n338) );
  XNOR2_X1 U642 ( .A(n572), .B(b[13]), .ZN(n378) );
  XNOR2_X1 U643 ( .A(n544), .B(n424), .ZN(n362) );
  XNOR2_X1 U644 ( .A(n573), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U645 ( .A(n573), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U646 ( .A(n573), .B(n418), .ZN(n384) );
  XNOR2_X1 U647 ( .A(n572), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U648 ( .A(n572), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U649 ( .A(n572), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U650 ( .A(n572), .B(n419), .ZN(n385) );
  XNOR2_X1 U651 ( .A(n576), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U652 ( .A(n576), .B(n418), .ZN(n369) );
  XNOR2_X1 U653 ( .A(n576), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U654 ( .A(n576), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U655 ( .A(n544), .B(n423), .ZN(n361) );
  XNOR2_X1 U656 ( .A(n544), .B(n422), .ZN(n360) );
  XNOR2_X1 U657 ( .A(n579), .B(n422), .ZN(n349) );
  XNOR2_X1 U658 ( .A(n579), .B(n423), .ZN(n350) );
  XNOR2_X1 U659 ( .A(n544), .B(n421), .ZN(n359) );
  XNOR2_X1 U660 ( .A(n544), .B(n420), .ZN(n358) );
  XNOR2_X1 U661 ( .A(n579), .B(n421), .ZN(n348) );
  XNOR2_X1 U662 ( .A(n579), .B(n420), .ZN(n347) );
  XNOR2_X1 U663 ( .A(n544), .B(n418), .ZN(n356) );
  XNOR2_X1 U664 ( .A(n579), .B(n419), .ZN(n346) );
  XNOR2_X1 U665 ( .A(n544), .B(n419), .ZN(n357) );
  XNOR2_X1 U666 ( .A(n544), .B(b[8]), .ZN(n355) );
  XNOR2_X1 U667 ( .A(n490), .B(b[15]), .ZN(n393) );
  BUF_X1 U668 ( .A(n43), .Z(n569) );
  XNOR2_X1 U669 ( .A(n1), .B(a[2]), .ZN(n9) );
  XNOR2_X1 U670 ( .A(n84), .B(n50), .ZN(product[11]) );
  NAND2_X1 U671 ( .A1(n329), .A2(n258), .ZN(n122) );
  NOR2_X1 U672 ( .A1(n82), .A2(n85), .ZN(n80) );
  OAI21_X1 U673 ( .B1(n502), .B2(n86), .A(n83), .ZN(n81) );
  NAND2_X1 U674 ( .A1(n186), .A2(n195), .ZN(n83) );
  NOR2_X1 U675 ( .A1(n234), .A2(n257), .ZN(n113) );
  NAND2_X1 U676 ( .A1(n567), .A2(n103), .ZN(n55) );
  INV_X1 U677 ( .A(n103), .ZN(n101) );
  NAND2_X1 U678 ( .A1(n224), .A2(n227), .ZN(n103) );
  INV_X1 U679 ( .A(n19), .ZN(n578) );
  NAND2_X1 U680 ( .A1(n204), .A2(n211), .ZN(n90) );
  NOR2_X1 U681 ( .A1(n204), .A2(n211), .ZN(n89) );
  OAI22_X1 U682 ( .A1(n29), .A2(n350), .B1(n349), .B2(n533), .ZN(n275) );
  OAI22_X1 U683 ( .A1(n503), .A2(n346), .B1(n345), .B2(n533), .ZN(n271) );
  OAI22_X1 U684 ( .A1(n503), .A2(n347), .B1(n346), .B2(n533), .ZN(n272) );
  OAI22_X1 U685 ( .A1(n29), .A2(n348), .B1(n347), .B2(n533), .ZN(n273) );
  OAI22_X1 U686 ( .A1(n29), .A2(n349), .B1(n348), .B2(n533), .ZN(n274) );
  OAI22_X1 U687 ( .A1(n29), .A2(n511), .B1(n353), .B2(n533), .ZN(n254) );
  OAI22_X1 U688 ( .A1(n29), .A2(n351), .B1(n350), .B2(n533), .ZN(n276) );
  OAI22_X1 U689 ( .A1(n29), .A2(n352), .B1(n351), .B2(n533), .ZN(n277) );
  NAND2_X1 U690 ( .A1(n151), .A2(n139), .ZN(n62) );
  INV_X1 U691 ( .A(n113), .ZN(n135) );
  XNOR2_X1 U692 ( .A(n77), .B(n48), .ZN(product[13]) );
  XNOR2_X1 U693 ( .A(n535), .B(n55), .ZN(product[6]) );
  OAI21_X1 U694 ( .B1(n87), .B2(n85), .A(n86), .ZN(n84) );
  INV_X1 U695 ( .A(n1), .ZN(n571) );
  OR2_X1 U696 ( .A1(n568), .A2(n513), .ZN(n409) );
  XNOR2_X1 U697 ( .A(n70), .B(n47), .ZN(product[14]) );
  OAI22_X1 U698 ( .A1(n512), .A2(n358), .B1(n357), .B2(n509), .ZN(n282) );
  OAI22_X1 U699 ( .A1(n512), .A2(n356), .B1(n355), .B2(n509), .ZN(n280) );
  OAI22_X1 U700 ( .A1(n23), .A2(n362), .B1(n361), .B2(n21), .ZN(n286) );
  OAI22_X1 U701 ( .A1(n512), .A2(n357), .B1(n356), .B2(n509), .ZN(n281) );
  OAI22_X1 U702 ( .A1(n23), .A2(n360), .B1(n359), .B2(n21), .ZN(n284) );
  OAI22_X1 U703 ( .A1(n23), .A2(n578), .B1(n364), .B2(n21), .ZN(n255) );
  OAI22_X1 U704 ( .A1(n23), .A2(n361), .B1(n360), .B2(n21), .ZN(n285) );
  OAI22_X1 U705 ( .A1(n512), .A2(n355), .B1(n354), .B2(n509), .ZN(n279) );
  OAI22_X1 U706 ( .A1(n23), .A2(n363), .B1(n362), .B2(n21), .ZN(n287) );
  OAI22_X1 U707 ( .A1(n23), .A2(n359), .B1(n358), .B2(n21), .ZN(n283) );
  XNOR2_X1 U708 ( .A(n575), .B(n421), .ZN(n372) );
  XNOR2_X1 U709 ( .A(n575), .B(n423), .ZN(n374) );
  XNOR2_X1 U710 ( .A(n575), .B(n424), .ZN(n375) );
  XNOR2_X1 U711 ( .A(n575), .B(n422), .ZN(n373) );
  XNOR2_X1 U712 ( .A(n575), .B(n419), .ZN(n370) );
  XNOR2_X1 U713 ( .A(n575), .B(n420), .ZN(n371) );
  XOR2_X1 U714 ( .A(n547), .B(n52), .Z(product[9]) );
  XNOR2_X1 U715 ( .A(n545), .B(n53), .ZN(product[8]) );
  OAI21_X1 U716 ( .B1(n493), .B2(n89), .A(n90), .ZN(n88) );
  AOI21_X1 U717 ( .B1(n96), .B2(n558), .A(n93), .ZN(n91) );
  OAI22_X1 U718 ( .A1(n18), .A2(n370), .B1(n369), .B2(n565), .ZN(n293) );
  OAI22_X1 U719 ( .A1(n500), .A2(n367), .B1(n366), .B2(n565), .ZN(n290) );
  OAI22_X1 U720 ( .A1(n500), .A2(n375), .B1(n374), .B2(n565), .ZN(n298) );
  OAI22_X1 U721 ( .A1(n18), .A2(n368), .B1(n367), .B2(n565), .ZN(n291) );
  OAI22_X1 U722 ( .A1(n501), .A2(n373), .B1(n372), .B2(n565), .ZN(n296) );
  OAI22_X1 U723 ( .A1(n500), .A2(n371), .B1(n370), .B2(n565), .ZN(n294) );
  OAI22_X1 U724 ( .A1(n500), .A2(n369), .B1(n368), .B2(n565), .ZN(n292) );
  OAI22_X1 U725 ( .A1(n501), .A2(n372), .B1(n371), .B2(n565), .ZN(n295) );
  OAI22_X1 U726 ( .A1(n500), .A2(n517), .B1(n377), .B2(n565), .ZN(n256) );
  OAI22_X1 U727 ( .A1(n501), .A2(n376), .B1(n375), .B2(n565), .ZN(n299) );
  OAI22_X1 U728 ( .A1(n18), .A2(n374), .B1(n565), .B2(n373), .ZN(n297) );
  OAI22_X1 U729 ( .A1(n501), .A2(n366), .B1(n365), .B2(n565), .ZN(n289) );
  XNOR2_X1 U730 ( .A(n572), .B(n420), .ZN(n386) );
  INV_X1 U731 ( .A(n565), .ZN(n245) );
  XNOR2_X1 U732 ( .A(n572), .B(n568), .ZN(n391) );
  XNOR2_X1 U733 ( .A(n573), .B(n423), .ZN(n389) );
  XNOR2_X1 U734 ( .A(n572), .B(n424), .ZN(n390) );
  XNOR2_X1 U735 ( .A(n573), .B(n422), .ZN(n388) );
  XNOR2_X1 U736 ( .A(n572), .B(n421), .ZN(n387) );
  INV_X1 U737 ( .A(n88), .ZN(n87) );
  XNOR2_X1 U738 ( .A(n525), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U739 ( .A(n490), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U740 ( .A(n490), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U741 ( .A(n510), .B(n418), .ZN(n401) );
  XNOR2_X1 U742 ( .A(n490), .B(n568), .ZN(n408) );
  XNOR2_X1 U743 ( .A(n510), .B(n422), .ZN(n405) );
  XNOR2_X1 U744 ( .A(n490), .B(n423), .ZN(n406) );
  XNOR2_X1 U745 ( .A(n510), .B(n421), .ZN(n404) );
  XNOR2_X1 U746 ( .A(n525), .B(n424), .ZN(n407) );
  XNOR2_X1 U747 ( .A(n525), .B(n419), .ZN(n402) );
  XNOR2_X1 U748 ( .A(n510), .B(n420), .ZN(n403) );
  OAI21_X1 U749 ( .B1(n107), .B2(n105), .A(n106), .ZN(n104) );
  OAI21_X1 U750 ( .B1(n64), .B2(n499), .A(n65), .ZN(n63) );
  OAI21_X1 U751 ( .B1(n45), .B2(n78), .A(n79), .ZN(n77) );
  OAI21_X1 U752 ( .B1(n499), .B2(n71), .A(n72), .ZN(n70) );
  XOR2_X1 U753 ( .A(n56), .B(n523), .Z(product[5]) );
  AOI21_X1 U754 ( .B1(n560), .B2(n120), .A(n117), .ZN(n115) );
  INV_X1 U755 ( .A(n122), .ZN(n120) );
  AOI21_X1 U756 ( .B1(n561), .B2(n112), .A(n498), .ZN(n107) );
  OAI22_X1 U757 ( .A1(n551), .A2(n513), .B1(n409), .B2(n543), .ZN(n258) );
  OAI22_X1 U758 ( .A1(n491), .A2(n379), .B1(n378), .B2(n566), .ZN(n301) );
  OAI22_X1 U759 ( .A1(n532), .A2(n380), .B1(n566), .B2(n379), .ZN(n302) );
  OAI22_X1 U760 ( .A1(n532), .A2(n385), .B1(n384), .B2(n566), .ZN(n307) );
  OAI22_X1 U761 ( .A1(n491), .A2(n382), .B1(n381), .B2(n566), .ZN(n304) );
  OAI22_X1 U762 ( .A1(n491), .A2(n381), .B1(n380), .B2(n566), .ZN(n303) );
  NAND2_X1 U763 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U764 ( .A1(n491), .A2(n383), .B1(n382), .B2(n566), .ZN(n305) );
  OAI22_X1 U765 ( .A1(n531), .A2(n384), .B1(n383), .B2(n566), .ZN(n306) );
  OAI22_X1 U766 ( .A1(n532), .A2(n386), .B1(n385), .B2(n566), .ZN(n308) );
  OAI22_X1 U767 ( .A1(n532), .A2(n387), .B1(n386), .B2(n566), .ZN(n309) );
  OAI22_X1 U768 ( .A1(n491), .A2(n522), .B1(n392), .B2(n566), .ZN(n257) );
  OAI22_X1 U769 ( .A1(n531), .A2(n389), .B1(n566), .B2(n388), .ZN(n311) );
  OAI22_X1 U770 ( .A1(n532), .A2(n388), .B1(n387), .B2(n566), .ZN(n310) );
  OAI22_X1 U771 ( .A1(n532), .A2(n390), .B1(n389), .B2(n566), .ZN(n312) );
  INV_X1 U772 ( .A(n566), .ZN(n247) );
  OAI22_X1 U773 ( .A1(n491), .A2(n391), .B1(n390), .B2(n566), .ZN(n313) );
  INV_X1 U774 ( .A(n517), .ZN(n576) );
  INV_X1 U775 ( .A(n31), .ZN(n582) );
  INV_X1 U776 ( .A(n584), .ZN(n583) );
  INV_X1 U777 ( .A(n36), .ZN(n584) );
  INV_X1 U778 ( .A(n586), .ZN(n585) );
  INV_X1 U779 ( .A(n40), .ZN(n586) );
  XOR2_X1 U780 ( .A(n259), .B(n251), .Z(n148) );
  XOR2_X1 U781 ( .A(n279), .B(n289), .Z(n146) );
  XOR2_X1 U782 ( .A(n159), .B(n150), .Z(n142) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_0_DW01_add_2 ( A, B, CI, SUM, 
        CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n18,
         n19, n20, n21, n25, n26, n27, n28, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n48, n49, n51, n53, n54, n55, n56, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n69, n71, n72, n73, n74, n75,
         n77, n79, n80, n81, n82, n83, n85, n87, n88, n90, n95, n98, n99, n100,
         n102, n104, n161, n162, n163, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187;

  NOR2_X1 U126 ( .A1(A[8]), .A2(B[8]), .ZN(n161) );
  INV_X1 U127 ( .A(n169), .ZN(n162) );
  NOR2_X1 U128 ( .A1(A[8]), .A2(B[8]), .ZN(n58) );
  OR2_X1 U129 ( .A1(A[15]), .A2(B[15]), .ZN(n163) );
  AND2_X1 U130 ( .A1(n177), .A2(n90), .ZN(SUM[0]) );
  INV_X1 U131 ( .A(n53), .ZN(n165) );
  INV_X1 U132 ( .A(n42), .ZN(n166) );
  OAI21_X1 U133 ( .B1(n58), .B2(n62), .A(n59), .ZN(n167) );
  AOI21_X1 U134 ( .B1(n186), .B2(n51), .A(n187), .ZN(n168) );
  AOI21_X1 U135 ( .B1(n56), .B2(n64), .A(n167), .ZN(n169) );
  OAI21_X1 U136 ( .B1(n43), .B2(n55), .A(n168), .ZN(n170) );
  BUF_X1 U137 ( .A(n37), .Z(n171) );
  AND2_X1 U138 ( .A1(A[13]), .A2(B[13]), .ZN(n172) );
  OR2_X1 U139 ( .A1(A[10]), .A2(B[10]), .ZN(n173) );
  CLKBUF_X1 U140 ( .A(A[12]), .Z(n174) );
  NOR2_X1 U141 ( .A1(B[12]), .A2(A[12]), .ZN(n175) );
  AOI21_X1 U142 ( .B1(n170), .B2(n34), .A(n35), .ZN(n176) );
  OR2_X1 U143 ( .A1(A[0]), .A2(B[0]), .ZN(n177) );
  INV_X1 U144 ( .A(n55), .ZN(n54) );
  INV_X1 U145 ( .A(n64), .ZN(n63) );
  INV_X1 U146 ( .A(n42), .ZN(n41) );
  OAI21_X1 U147 ( .B1(n83), .B2(n81), .A(n82), .ZN(n80) );
  AOI21_X1 U148 ( .B1(n181), .B2(n80), .A(n77), .ZN(n75) );
  AOI21_X1 U149 ( .B1(n56), .B2(n64), .A(n167), .ZN(n55) );
  AOI21_X1 U150 ( .B1(n162), .B2(n178), .A(n51), .ZN(n49) );
  INV_X1 U151 ( .A(n90), .ZN(n88) );
  INV_X1 U152 ( .A(n53), .ZN(n51) );
  AOI21_X1 U153 ( .B1(n179), .B2(n88), .A(n85), .ZN(n83) );
  INV_X1 U154 ( .A(n87), .ZN(n85) );
  INV_X1 U155 ( .A(n39), .ZN(n95) );
  NAND2_X1 U156 ( .A1(n98), .A2(n59), .ZN(n8) );
  INV_X1 U157 ( .A(n161), .ZN(n98) );
  NAND2_X1 U158 ( .A1(n178), .A2(n53), .ZN(n7) );
  NAND2_X1 U159 ( .A1(n104), .A2(n82), .ZN(n14) );
  INV_X1 U160 ( .A(n81), .ZN(n104) );
  NAND2_X1 U161 ( .A1(n102), .A2(n74), .ZN(n12) );
  INV_X1 U162 ( .A(n73), .ZN(n102) );
  NAND2_X1 U163 ( .A1(n179), .A2(n87), .ZN(n15) );
  NAND2_X1 U164 ( .A1(n99), .A2(n62), .ZN(n9) );
  NAND2_X1 U165 ( .A1(n181), .A2(n79), .ZN(n13) );
  NAND2_X1 U166 ( .A1(n182), .A2(n71), .ZN(n11) );
  NAND2_X1 U167 ( .A1(n100), .A2(n66), .ZN(n10) );
  INV_X1 U168 ( .A(n65), .ZN(n100) );
  INV_X1 U169 ( .A(n71), .ZN(n69) );
  XOR2_X1 U170 ( .A(n41), .B(n5), .Z(SUM[11]) );
  NAND2_X1 U171 ( .A1(n95), .A2(n40), .ZN(n5) );
  XNOR2_X1 U172 ( .A(n60), .B(n8), .ZN(SUM[8]) );
  XOR2_X1 U173 ( .A(n63), .B(n9), .Z(SUM[7]) );
  XOR2_X1 U174 ( .A(n12), .B(n75), .Z(SUM[4]) );
  XNOR2_X1 U175 ( .A(n15), .B(n88), .ZN(SUM[1]) );
  AOI21_X1 U176 ( .B1(n170), .B2(n34), .A(n35), .ZN(n33) );
  NOR2_X1 U177 ( .A1(A[11]), .A2(B[11]), .ZN(n39) );
  OR2_X1 U178 ( .A1(A[9]), .A2(B[9]), .ZN(n178) );
  NAND2_X1 U179 ( .A1(n183), .A2(n171), .ZN(n4) );
  XOR2_X1 U180 ( .A(n49), .B(n6), .Z(SUM[10]) );
  NAND2_X1 U181 ( .A1(A[11]), .A2(B[11]), .ZN(n40) );
  OR2_X1 U182 ( .A1(A[1]), .A2(B[1]), .ZN(n179) );
  OR2_X1 U183 ( .A1(A[14]), .A2(B[14]), .ZN(n180) );
  NOR2_X1 U184 ( .A1(A[2]), .A2(B[2]), .ZN(n81) );
  XNOR2_X1 U185 ( .A(n54), .B(n7), .ZN(SUM[9]) );
  NOR2_X1 U186 ( .A1(A[4]), .A2(B[4]), .ZN(n73) );
  NOR2_X1 U187 ( .A1(A[6]), .A2(B[6]), .ZN(n65) );
  OR2_X1 U188 ( .A1(A[3]), .A2(B[3]), .ZN(n181) );
  NAND2_X1 U189 ( .A1(A[5]), .A2(B[5]), .ZN(n71) );
  NAND2_X1 U190 ( .A1(A[1]), .A2(B[1]), .ZN(n87) );
  NAND2_X1 U191 ( .A1(A[0]), .A2(B[0]), .ZN(n90) );
  NAND2_X1 U192 ( .A1(A[2]), .A2(B[2]), .ZN(n82) );
  OR2_X1 U193 ( .A1(A[5]), .A2(B[5]), .ZN(n182) );
  NAND2_X1 U194 ( .A1(A[8]), .A2(B[8]), .ZN(n59) );
  NAND2_X1 U195 ( .A1(A[4]), .A2(B[4]), .ZN(n74) );
  NAND2_X1 U196 ( .A1(A[6]), .A2(B[6]), .ZN(n66) );
  NAND2_X1 U197 ( .A1(A[7]), .A2(B[7]), .ZN(n62) );
  NAND2_X1 U198 ( .A1(A[3]), .A2(B[3]), .ZN(n79) );
  XNOR2_X1 U199 ( .A(n13), .B(n80), .ZN(SUM[3]) );
  XOR2_X1 U200 ( .A(n14), .B(n83), .Z(SUM[2]) );
  OR2_X1 U201 ( .A1(A[10]), .A2(B[10]), .ZN(n186) );
  OR2_X1 U202 ( .A1(A[13]), .A2(B[13]), .ZN(n185) );
  NAND2_X1 U203 ( .A1(n163), .A2(n18), .ZN(n1) );
  OR2_X1 U204 ( .A1(n174), .A2(B[12]), .ZN(n183) );
  NAND2_X1 U205 ( .A1(n185), .A2(n28), .ZN(n3) );
  NAND2_X1 U206 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  NOR2_X1 U207 ( .A1(n161), .A2(n61), .ZN(n56) );
  OAI21_X1 U208 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  INV_X1 U209 ( .A(n61), .ZN(n99) );
  NOR2_X1 U210 ( .A1(A[7]), .A2(B[7]), .ZN(n61) );
  AND2_X1 U211 ( .A1(A[14]), .A2(B[14]), .ZN(n184) );
  INV_X1 U212 ( .A(n187), .ZN(n48) );
  NAND2_X1 U213 ( .A1(n173), .A2(n48), .ZN(n6) );
  NAND2_X1 U214 ( .A1(A[9]), .A2(B[9]), .ZN(n53) );
  AND2_X1 U215 ( .A1(A[10]), .A2(B[10]), .ZN(n187) );
  NAND2_X1 U216 ( .A1(n180), .A2(n25), .ZN(n2) );
  NAND2_X1 U217 ( .A1(n180), .A2(n185), .ZN(n20) );
  AOI21_X1 U218 ( .B1(n180), .B2(n172), .A(n184), .ZN(n21) );
  XNOR2_X1 U219 ( .A(n11), .B(n72), .ZN(SUM[5]) );
  XOR2_X1 U220 ( .A(n10), .B(n67), .Z(SUM[6]) );
  OAI21_X1 U221 ( .B1(n67), .B2(n65), .A(n66), .ZN(n64) );
  AOI21_X1 U222 ( .B1(n182), .B2(n72), .A(n69), .ZN(n67) );
  OAI21_X1 U223 ( .B1(n36), .B2(n40), .A(n37), .ZN(n35) );
  NOR2_X1 U224 ( .A1(n175), .A2(n39), .ZN(n34) );
  NOR2_X1 U225 ( .A1(A[12]), .A2(B[12]), .ZN(n36) );
  NAND2_X1 U226 ( .A1(A[12]), .A2(B[12]), .ZN(n37) );
  NOR2_X1 U227 ( .A1(A[13]), .A2(B[13]), .ZN(n27) );
  XNOR2_X1 U228 ( .A(n26), .B(n2), .ZN(SUM[14]) );
  OAI21_X1 U229 ( .B1(n166), .B2(n39), .A(n40), .ZN(n38) );
  INV_X1 U230 ( .A(n79), .ZN(n77) );
  OAI21_X1 U231 ( .B1(n75), .B2(n73), .A(n74), .ZN(n72) );
  NAND2_X1 U232 ( .A1(A[14]), .A2(B[14]), .ZN(n25) );
  NAND2_X1 U233 ( .A1(A[15]), .A2(B[15]), .ZN(n18) );
  NAND2_X1 U234 ( .A1(n173), .A2(n178), .ZN(n43) );
  AOI21_X1 U235 ( .B1(n186), .B2(n165), .A(n187), .ZN(n44) );
  XNOR2_X1 U236 ( .A(n38), .B(n4), .ZN(SUM[12]) );
  XNOR2_X1 U237 ( .A(n19), .B(n1), .ZN(SUM[15]) );
  XOR2_X1 U238 ( .A(n33), .B(n3), .Z(SUM[13]) );
  OAI21_X1 U239 ( .B1(n33), .B2(n20), .A(n21), .ZN(n19) );
  OAI21_X1 U240 ( .B1(n176), .B2(n27), .A(n28), .ZN(n26) );
  OAI21_X1 U241 ( .B1(n169), .B2(n43), .A(n44), .ZN(n42) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_0 ( clk, clear_acc, 
        data_out_x, data_out, data_out_w, data_out_b, wr_en_y, m_valid, 
        m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [3:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N27, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, n30, n31, n86, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n105,
         n106, n107, n108, n109, n110, n111, n112, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n13), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n103), .CK(clk), .Q(n17) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n102), .CK(clk), .Q(n18) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n101), .CK(clk), .Q(n19) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n100), .CK(clk), .Q(n20) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n96), .CK(clk), .Q(n24) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n95), .CK(clk), .Q(n25) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n94), .CK(clk), .Q(n26) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n93), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n92), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n91), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n90), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n89), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n88), .CK(clk), .Q(n34) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_0_DW_mult_tc_1 mult_960 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_0_DW01_add_2 add_961 ( .A({n129, 
        n130, n131, n132, n133, n134, n120, n121, n122, n123, n124, n125, n126, 
        n127, n128, n135}), .B({f[15], n38, n39, n41, n43, n45, f[9:3], n53, 
        n55, n57}), .CI(1'b0), .SUM(adder) );
  DFF_X1 delay_reg ( .D(N27), .CK(clk), .Q(n2), .QN(n86) );
  DFF_X1 \data_out_reg[15]  ( .D(n167), .CK(clk), .Q(data_out[15]), .QN(n136)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n166), .CK(clk), .Q(data_out[14]), .QN(n137)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n165), .CK(clk), .Q(data_out[13]), .QN(n138)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n164), .CK(clk), .Q(data_out[12]), .QN(n139)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n163), .CK(clk), .Q(data_out[11]), .QN(n140)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n162), .CK(clk), .Q(data_out[10]), .QN(n141)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n161), .CK(clk), .Q(data_out[9]), .QN(n142) );
  DFF_X1 \data_out_reg[8]  ( .D(n160), .CK(clk), .Q(data_out[8]), .QN(n143) );
  DFF_X1 \data_out_reg[7]  ( .D(n159), .CK(clk), .Q(data_out[7]), .QN(n144) );
  DFF_X1 \data_out_reg[6]  ( .D(n158), .CK(clk), .Q(data_out[6]), .QN(n145) );
  DFF_X1 \data_out_reg[5]  ( .D(n157), .CK(clk), .Q(data_out[5]), .QN(n146) );
  DFF_X1 \data_out_reg[4]  ( .D(n156), .CK(clk), .Q(data_out[4]), .QN(n147) );
  DFF_X1 \data_out_reg[3]  ( .D(n155), .CK(clk), .Q(data_out[3]), .QN(n148) );
  DFF_X1 \data_out_reg[2]  ( .D(n154), .CK(clk), .Q(data_out[2]), .QN(n149) );
  DFF_X1 \data_out_reg[1]  ( .D(n153), .CK(clk), .Q(data_out[1]), .QN(n150) );
  DFF_X1 \data_out_reg[0]  ( .D(n152), .CK(clk), .Q(data_out[0]), .QN(n151) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n97), .CK(clk), .Q(n23) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n98), .CK(clk), .Q(n22) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n99), .CK(clk), .Q(n21) );
  DFF_X1 \f_reg[3]  ( .D(n82), .CK(clk), .Q(f[3]), .QN(n61) );
  DFF_X1 \f_reg[2]  ( .D(n83), .CK(clk), .Q(n53), .QN(n117) );
  DFF_X1 \f_reg[4]  ( .D(n81), .CK(clk), .Q(f[4]), .QN(n62) );
  DFF_X1 \f_reg[1]  ( .D(n84), .CK(clk), .Q(n55), .QN(n118) );
  DFF_X1 \f_reg[0]  ( .D(n85), .CK(clk), .Q(n57), .QN(n119) );
  DFF_X1 \f_reg[5]  ( .D(n80), .CK(clk), .Q(f[5]), .QN(n63) );
  DFF_X1 \f_reg[6]  ( .D(n79), .CK(clk), .Q(f[6]), .QN(n64) );
  DFF_X1 \f_reg[7]  ( .D(n78), .CK(clk), .Q(f[7]), .QN(n112) );
  DFF_X1 \f_reg[8]  ( .D(n77), .CK(clk), .Q(f[8]), .QN(n111) );
  DFF_X1 \f_reg[9]  ( .D(n76), .CK(clk), .Q(f[9]), .QN(n110) );
  DFF_X1 \f_reg[10]  ( .D(n75), .CK(clk), .Q(n45), .QN(n109) );
  DFF_X1 \f_reg[11]  ( .D(n74), .CK(clk), .Q(n43), .QN(n108) );
  DFF_X1 \f_reg[14]  ( .D(n71), .CK(clk), .Q(n38), .QN(n105) );
  DFF_X1 \f_reg[13]  ( .D(n72), .CK(clk), .Q(n39), .QN(n106) );
  DFF_X1 \f_reg[15]  ( .D(n7), .CK(clk), .Q(f[15]), .QN(n69) );
  DFF_X1 \f_reg[12]  ( .D(n73), .CK(clk), .Q(n41), .QN(n107) );
  AND2_X2 U3 ( .A1(n37), .A2(n14), .ZN(n11) );
  AND2_X1 U4 ( .A1(clear_acc_delay), .A2(n86), .ZN(n1) );
  INV_X1 U5 ( .A(clear_acc), .ZN(n14) );
  MUX2_X2 U6 ( .A(n24), .B(N37), .S(n86), .Z(n121) );
  MUX2_X2 U8 ( .A(n22), .B(N39), .S(n86), .Z(n134) );
  OAI222_X1 U9 ( .A1(n4), .A2(n14), .B1(n5), .B2(n6), .C1(n105), .C2(n37), 
        .ZN(n71) );
  INV_X1 U10 ( .A(data_out_b[14]), .ZN(n4) );
  INV_X1 U11 ( .A(adder[14]), .ZN(n5) );
  INV_X1 U12 ( .A(n11), .ZN(n6) );
  NAND3_X1 U13 ( .A1(n9), .A2(n8), .A3(n10), .ZN(n7) );
  MUX2_X1 U14 ( .A(n19), .B(N42), .S(n86), .Z(n131) );
  NAND2_X1 U15 ( .A1(data_out_b[15]), .A2(n13), .ZN(n8) );
  NAND2_X1 U16 ( .A1(adder[15]), .A2(n11), .ZN(n9) );
  NAND2_X1 U17 ( .A1(n59), .A2(f[15]), .ZN(n10) );
  INV_X2 U18 ( .A(n37), .ZN(n59) );
  MUX2_X2 U19 ( .A(n20), .B(N41), .S(n86), .Z(n132) );
  NAND2_X1 U20 ( .A1(n12), .A2(N27), .ZN(n30) );
  OAI22_X1 U21 ( .A1(n148), .A2(n30), .B1(n61), .B2(n31), .ZN(n155) );
  OAI22_X1 U22 ( .A1(n147), .A2(n30), .B1(n62), .B2(n31), .ZN(n156) );
  OAI22_X1 U23 ( .A1(n146), .A2(n30), .B1(n63), .B2(n31), .ZN(n157) );
  OAI22_X1 U24 ( .A1(n145), .A2(n30), .B1(n64), .B2(n31), .ZN(n158) );
  OAI22_X1 U25 ( .A1(n144), .A2(n30), .B1(n112), .B2(n31), .ZN(n159) );
  OAI22_X1 U26 ( .A1(n143), .A2(n30), .B1(n111), .B2(n31), .ZN(n160) );
  OAI22_X1 U27 ( .A1(n142), .A2(n30), .B1(n110), .B2(n31), .ZN(n161) );
  MUX2_X1 U28 ( .A(n29), .B(N32), .S(n86), .Z(n126) );
  MUX2_X1 U29 ( .A(n18), .B(N43), .S(n86), .Z(n130) );
  INV_X1 U30 ( .A(wr_en_y), .ZN(n12) );
  INV_X1 U31 ( .A(n14), .ZN(n13) );
  AND2_X1 U32 ( .A1(sel[0]), .A2(sel[1]), .ZN(n16) );
  INV_X1 U33 ( .A(m_ready), .ZN(n15) );
  NAND2_X1 U34 ( .A1(m_valid), .A2(n15), .ZN(n35) );
  OAI211_X1 U35 ( .C1(sel[2]), .C2(n16), .A(sel[3]), .B(n35), .ZN(N27) );
  MUX2_X1 U36 ( .A(n17), .B(N44), .S(n1), .Z(n103) );
  MUX2_X1 U37 ( .A(n17), .B(N44), .S(n86), .Z(n129) );
  MUX2_X1 U38 ( .A(n18), .B(N43), .S(n1), .Z(n102) );
  MUX2_X1 U39 ( .A(n19), .B(N42), .S(n1), .Z(n101) );
  MUX2_X1 U40 ( .A(n20), .B(N41), .S(n1), .Z(n100) );
  MUX2_X1 U41 ( .A(n21), .B(N40), .S(n1), .Z(n99) );
  MUX2_X1 U42 ( .A(n21), .B(N40), .S(n86), .Z(n133) );
  MUX2_X1 U43 ( .A(n22), .B(N39), .S(n1), .Z(n98) );
  MUX2_X1 U44 ( .A(n23), .B(N38), .S(n1), .Z(n97) );
  MUX2_X1 U45 ( .A(n23), .B(N38), .S(n86), .Z(n120) );
  MUX2_X1 U46 ( .A(n24), .B(N37), .S(n1), .Z(n96) );
  MUX2_X1 U47 ( .A(n25), .B(N36), .S(n1), .Z(n95) );
  MUX2_X1 U48 ( .A(n25), .B(N36), .S(n86), .Z(n122) );
  MUX2_X1 U49 ( .A(n26), .B(N35), .S(n1), .Z(n94) );
  MUX2_X1 U50 ( .A(n26), .B(N35), .S(n86), .Z(n123) );
  MUX2_X1 U51 ( .A(n27), .B(N34), .S(n1), .Z(n93) );
  MUX2_X1 U52 ( .A(n27), .B(N34), .S(n86), .Z(n124) );
  MUX2_X1 U53 ( .A(n28), .B(N33), .S(n1), .Z(n92) );
  MUX2_X1 U54 ( .A(n28), .B(N33), .S(n86), .Z(n125) );
  MUX2_X1 U55 ( .A(n29), .B(N32), .S(n1), .Z(n91) );
  MUX2_X1 U56 ( .A(n32), .B(N31), .S(n1), .Z(n90) );
  MUX2_X1 U57 ( .A(n32), .B(N31), .S(n86), .Z(n127) );
  MUX2_X1 U58 ( .A(n33), .B(N30), .S(n1), .Z(n89) );
  MUX2_X1 U59 ( .A(n33), .B(N30), .S(n86), .Z(n128) );
  MUX2_X1 U60 ( .A(n34), .B(N29), .S(n1), .Z(n88) );
  MUX2_X1 U61 ( .A(n34), .B(N29), .S(n86), .Z(n135) );
  INV_X1 U62 ( .A(n35), .ZN(n36) );
  OAI21_X1 U63 ( .B1(n36), .B2(n2), .A(n14), .ZN(n37) );
  AOI222_X1 U64 ( .A1(data_out_b[13]), .A2(n13), .B1(adder[13]), .B2(n11), 
        .C1(n59), .C2(n39), .ZN(n40) );
  INV_X1 U65 ( .A(n40), .ZN(n72) );
  AOI222_X1 U66 ( .A1(data_out_b[12]), .A2(n13), .B1(adder[12]), .B2(n11), 
        .C1(n59), .C2(n41), .ZN(n42) );
  INV_X1 U67 ( .A(n42), .ZN(n73) );
  AOI222_X1 U68 ( .A1(data_out_b[11]), .A2(n13), .B1(adder[11]), .B2(n11), 
        .C1(n59), .C2(n43), .ZN(n44) );
  INV_X1 U69 ( .A(n44), .ZN(n74) );
  AOI222_X1 U70 ( .A1(data_out_b[10]), .A2(n13), .B1(adder[10]), .B2(n11), 
        .C1(n59), .C2(n45), .ZN(n46) );
  INV_X1 U71 ( .A(n46), .ZN(n75) );
  AOI222_X1 U72 ( .A1(data_out_b[8]), .A2(n13), .B1(adder[8]), .B2(n11), .C1(
        n59), .C2(f[8]), .ZN(n47) );
  INV_X1 U73 ( .A(n47), .ZN(n77) );
  AOI222_X1 U74 ( .A1(data_out_b[7]), .A2(n13), .B1(adder[7]), .B2(n11), .C1(
        n59), .C2(f[7]), .ZN(n48) );
  INV_X1 U75 ( .A(n48), .ZN(n78) );
  AOI222_X1 U76 ( .A1(data_out_b[6]), .A2(n13), .B1(adder[6]), .B2(n11), .C1(
        n59), .C2(f[6]), .ZN(n49) );
  INV_X1 U77 ( .A(n49), .ZN(n79) );
  AOI222_X1 U78 ( .A1(data_out_b[5]), .A2(n13), .B1(adder[5]), .B2(n11), .C1(
        n59), .C2(f[5]), .ZN(n50) );
  INV_X1 U79 ( .A(n50), .ZN(n80) );
  AOI222_X1 U80 ( .A1(data_out_b[4]), .A2(n13), .B1(adder[4]), .B2(n11), .C1(
        n59), .C2(f[4]), .ZN(n51) );
  INV_X1 U81 ( .A(n51), .ZN(n81) );
  AOI222_X1 U82 ( .A1(data_out_b[3]), .A2(n13), .B1(adder[3]), .B2(n11), .C1(
        n59), .C2(f[3]), .ZN(n52) );
  INV_X1 U83 ( .A(n52), .ZN(n82) );
  AOI222_X1 U84 ( .A1(data_out_b[2]), .A2(n13), .B1(adder[2]), .B2(n11), .C1(
        n59), .C2(n53), .ZN(n54) );
  INV_X1 U85 ( .A(n54), .ZN(n83) );
  AOI222_X1 U86 ( .A1(data_out_b[1]), .A2(n13), .B1(adder[1]), .B2(n11), .C1(
        n59), .C2(n55), .ZN(n56) );
  INV_X1 U87 ( .A(n56), .ZN(n84) );
  AOI222_X1 U88 ( .A1(data_out_b[0]), .A2(n13), .B1(adder[0]), .B2(n11), .C1(
        n59), .C2(n57), .ZN(n58) );
  INV_X1 U89 ( .A(n58), .ZN(n85) );
  AOI222_X1 U90 ( .A1(data_out_b[9]), .A2(n13), .B1(adder[9]), .B2(n11), .C1(
        n59), .C2(f[9]), .ZN(n60) );
  INV_X1 U91 ( .A(n60), .ZN(n76) );
  NOR4_X1 U92 ( .A1(n43), .A2(n41), .A3(n39), .A4(n38), .ZN(n68) );
  NOR4_X1 U93 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n45), .ZN(n67) );
  NAND4_X1 U94 ( .A1(n64), .A2(n63), .A3(n62), .A4(n61), .ZN(n65) );
  NOR4_X1 U95 ( .A1(n65), .A2(n57), .A3(n55), .A4(n53), .ZN(n66) );
  NAND3_X1 U96 ( .A1(n68), .A2(n67), .A3(n66), .ZN(n70) );
  NAND3_X1 U97 ( .A1(wr_en_y), .A2(n70), .A3(n69), .ZN(n31) );
  OAI22_X1 U98 ( .A1(n151), .A2(n30), .B1(n119), .B2(n31), .ZN(n152) );
  OAI22_X1 U99 ( .A1(n150), .A2(n30), .B1(n118), .B2(n31), .ZN(n153) );
  OAI22_X1 U100 ( .A1(n149), .A2(n30), .B1(n117), .B2(n31), .ZN(n154) );
  OAI22_X1 U101 ( .A1(n141), .A2(n30), .B1(n109), .B2(n31), .ZN(n162) );
  OAI22_X1 U102 ( .A1(n140), .A2(n30), .B1(n108), .B2(n31), .ZN(n163) );
  OAI22_X1 U103 ( .A1(n139), .A2(n30), .B1(n107), .B2(n31), .ZN(n164) );
  OAI22_X1 U104 ( .A1(n138), .A2(n30), .B1(n106), .B2(n31), .ZN(n165) );
  OAI22_X1 U105 ( .A1(n137), .A2(n30), .B1(n105), .B2(n31), .ZN(n166) );
  OAI22_X1 U106 ( .A1(n136), .A2(n30), .B1(n69), .B2(n31), .ZN(n167) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_11_DW_mult_tc_1 ( a, b, 
        product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n9, n12, n13, n16, n18, n19, n21, n23, n25, n27, n29, n31,
         n32, n34, n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n50,
         n52, n53, n54, n55, n56, n57, n58, n59, n62, n63, n64, n65, n67, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n93, n95, n96, n97, n98, n99,
         n101, n103, n104, n105, n106, n107, n109, n111, n112, n113, n114,
         n115, n117, n119, n120, n122, n125, n127, n129, n131, n133, n135,
         n139, n141, n142, n143, n144, n145, n146, n147, n148, n149, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n230, n231, n232, n233, n234, n235, n237, n241, n247, n249, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n418, n419, n420, n421, n422, n423, n424,
         n426, n427, n429, n431, n433, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U148 ( .A(n265), .B(n144), .Z(n145) );
  XOR2_X1 U150 ( .A(n271), .B(n146), .Z(n147) );
  XOR2_X1 U152 ( .A(n148), .B(n301), .Z(n149) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n263), .CI(n291), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n317), .B(n252), .CO(n173), .S(n174) );
  FA_X1 U167 ( .A(n180), .B(n187), .CI(n178), .CO(n175), .S(n176) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U169 ( .A(n193), .B(n282), .CI(n191), .CO(n179), .S(n180) );
  FA_X1 U170 ( .A(n268), .B(n292), .CI(n274), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U172 ( .A(n197), .B(n190), .CI(n188), .CO(n185), .S(n186) );
  FA_X1 U173 ( .A(n199), .B(n201), .CI(n192), .CO(n187), .S(n188) );
  FA_X1 U174 ( .A(n275), .B(n293), .CI(n194), .CO(n189), .S(n190) );
  FA_X1 U175 ( .A(n253), .B(n283), .CI(n305), .CO(n191), .S(n192) );
  HA_X1 U176 ( .A(n269), .B(n319), .CO(n193), .S(n194) );
  FA_X1 U177 ( .A(n205), .B(n200), .CI(n198), .CO(n195), .S(n196) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U179 ( .A(n276), .B(n294), .CI(n284), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n320), .B(n270), .CI(n306), .CO(n201), .S(n202) );
  FA_X1 U183 ( .A(n254), .B(n285), .CI(n295), .CO(n207), .S(n208) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U185 ( .A(n216), .B(n219), .CI(n214), .CO(n211), .S(n212) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n322), .B(n278), .CI(n308), .CO(n215), .S(n216) );
  FA_X1 U188 ( .A(n225), .B(n222), .CI(n220), .CO(n217), .S(n218) );
  FA_X1 U189 ( .A(n255), .B(n309), .CI(n297), .CO(n219), .S(n220) );
  HA_X1 U190 ( .A(n287), .B(n323), .CO(n221), .S(n222) );
  FA_X1 U192 ( .A(n324), .B(n288), .CI(n310), .CO(n225), .S(n226) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  FA_X1 U195 ( .A(n326), .B(n300), .CI(n312), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  INV_X2 U414 ( .A(n542), .ZN(n515) );
  BUF_X1 U415 ( .A(a[6]), .Z(n490) );
  NOR2_X1 U416 ( .A1(n164), .A2(n175), .ZN(n75) );
  NOR2_X1 U417 ( .A1(n176), .A2(n185), .ZN(n78) );
  AND2_X1 U418 ( .A1(n311), .A2(n325), .ZN(n491) );
  OR2_X1 U419 ( .A1(n329), .A2(n258), .ZN(n492) );
  BUF_X1 U420 ( .A(n584), .Z(n493) );
  NAND2_X1 U421 ( .A1(n429), .A2(n27), .ZN(n494) );
  NAND2_X1 U422 ( .A1(n429), .A2(n27), .ZN(n29) );
  BUF_X1 U423 ( .A(n83), .Z(n495) );
  INV_X1 U424 ( .A(n584), .ZN(n582) );
  XNOR2_X1 U425 ( .A(n493), .B(a[4]), .ZN(n431) );
  INV_X1 U426 ( .A(n501), .ZN(n496) );
  INV_X1 U427 ( .A(n501), .ZN(n576) );
  INV_X1 U428 ( .A(n580), .ZN(n497) );
  INV_X2 U429 ( .A(n581), .ZN(n580) );
  BUF_X2 U430 ( .A(n27), .Z(n498) );
  XNOR2_X1 U431 ( .A(a[8]), .B(n19), .ZN(n27) );
  INV_X1 U432 ( .A(n590), .ZN(n499) );
  INV_X1 U433 ( .A(n590), .ZN(n589) );
  XOR2_X1 U434 ( .A(n501), .B(a[2]), .Z(n9) );
  INV_X1 U435 ( .A(n586), .ZN(n500) );
  INV_X1 U436 ( .A(n1), .ZN(n501) );
  XOR2_X1 U437 ( .A(n572), .B(b[13]), .Z(n395) );
  INV_X1 U438 ( .A(n588), .ZN(n502) );
  INV_X1 U439 ( .A(n588), .ZN(n587) );
  BUF_X2 U440 ( .A(n37), .Z(n503) );
  XNOR2_X1 U441 ( .A(n504), .B(n210), .ZN(n206) );
  XNOR2_X1 U442 ( .A(n215), .B(n307), .ZN(n504) );
  INV_X1 U443 ( .A(n550), .ZN(n505) );
  INV_X1 U444 ( .A(n550), .ZN(n585) );
  OAI22_X1 U445 ( .A1(n539), .A2(n389), .B1(n388), .B2(n512), .ZN(n506) );
  BUF_X2 U446 ( .A(n533), .Z(n511) );
  CLKBUF_X1 U447 ( .A(n86), .Z(n507) );
  OR2_X1 U448 ( .A1(n176), .A2(n185), .ZN(n508) );
  XNOR2_X1 U449 ( .A(n509), .B(n166), .ZN(n164) );
  XNOR2_X1 U450 ( .A(n177), .B(n168), .ZN(n509) );
  BUF_X1 U451 ( .A(n12), .Z(n539) );
  OAI21_X1 U452 ( .B1(n113), .B2(n115), .A(n114), .ZN(n510) );
  BUF_X2 U453 ( .A(n533), .Z(n512) );
  XNOR2_X1 U454 ( .A(n577), .B(a[2]), .ZN(n533) );
  OR2_X1 U455 ( .A1(n196), .A2(n203), .ZN(n513) );
  NOR2_X1 U456 ( .A1(n186), .A2(n195), .ZN(n514) );
  NOR2_X1 U457 ( .A1(n186), .A2(n195), .ZN(n82) );
  NOR2_X1 U458 ( .A1(n196), .A2(n203), .ZN(n85) );
  INV_X1 U459 ( .A(n542), .ZN(n16) );
  INV_X1 U460 ( .A(n16), .ZN(n516) );
  XNOR2_X1 U461 ( .A(n226), .B(n517), .ZN(n224) );
  XNOR2_X1 U462 ( .A(n491), .B(n298), .ZN(n517) );
  OR2_X2 U463 ( .A1(n518), .A2(n534), .ZN(n34) );
  XNOR2_X1 U464 ( .A(n589), .B(a[10]), .ZN(n518) );
  INV_X1 U465 ( .A(n534), .ZN(n32) );
  INV_X1 U466 ( .A(n578), .ZN(n577) );
  OR2_X2 U467 ( .A1(n519), .A2(n560), .ZN(n23) );
  XNOR2_X1 U468 ( .A(n585), .B(n490), .ZN(n519) );
  OAI21_X1 U469 ( .B1(n105), .B2(n107), .A(n106), .ZN(n520) );
  AOI21_X2 U470 ( .B1(n567), .B2(n112), .A(n109), .ZN(n107) );
  XOR2_X1 U471 ( .A(n170), .B(n172), .Z(n521) );
  XOR2_X1 U472 ( .A(n521), .B(n179), .Z(n166) );
  NAND2_X1 U473 ( .A1(n170), .A2(n172), .ZN(n522) );
  NAND2_X1 U474 ( .A1(n170), .A2(n179), .ZN(n523) );
  NAND2_X1 U475 ( .A1(n172), .A2(n179), .ZN(n524) );
  NAND3_X1 U476 ( .A1(n522), .A2(n523), .A3(n524), .ZN(n165) );
  NAND2_X1 U477 ( .A1(n177), .A2(n168), .ZN(n525) );
  NAND2_X1 U478 ( .A1(n177), .A2(n166), .ZN(n526) );
  NAND2_X1 U479 ( .A1(n168), .A2(n166), .ZN(n527) );
  NAND3_X1 U480 ( .A1(n525), .A2(n526), .A3(n527), .ZN(n163) );
  INV_X1 U481 ( .A(n560), .ZN(n21) );
  BUF_X2 U482 ( .A(n575), .Z(n528) );
  INV_X1 U483 ( .A(n249), .ZN(n575) );
  OR2_X1 U484 ( .A1(n402), .A2(n575), .ZN(n557) );
  XNOR2_X1 U485 ( .A(n581), .B(a[2]), .ZN(n561) );
  INV_X1 U486 ( .A(n581), .ZN(n579) );
  XNOR2_X1 U487 ( .A(n45), .B(n529), .ZN(product[12]) );
  AND2_X1 U488 ( .A1(n508), .A2(n79), .ZN(n529) );
  BUF_X2 U489 ( .A(n12), .Z(n540) );
  CLKBUF_X1 U490 ( .A(n74), .Z(n530) );
  XNOR2_X1 U491 ( .A(n578), .B(n249), .ZN(n433) );
  XNOR2_X1 U492 ( .A(n88), .B(n531), .ZN(product[10]) );
  NAND2_X1 U493 ( .A1(n513), .A2(n86), .ZN(n531) );
  AOI21_X1 U494 ( .B1(n96), .B2(n563), .A(n93), .ZN(n532) );
  AOI21_X1 U495 ( .B1(n96), .B2(n563), .A(n93), .ZN(n91) );
  XNOR2_X1 U496 ( .A(n588), .B(a[10]), .ZN(n534) );
  OAI21_X1 U497 ( .B1(n532), .B2(n89), .A(n90), .ZN(n535) );
  AOI21_X1 U498 ( .B1(n566), .B2(n520), .A(n101), .ZN(n536) );
  NAND2_X2 U499 ( .A1(n433), .A2(n575), .ZN(n537) );
  NAND2_X1 U500 ( .A1(n433), .A2(n575), .ZN(n6) );
  XOR2_X1 U501 ( .A(n506), .B(n325), .Z(n230) );
  AOI21_X1 U502 ( .B1(n80), .B2(n535), .A(n81), .ZN(n538) );
  BUF_X2 U503 ( .A(n12), .Z(n541) );
  AOI21_X1 U504 ( .B1(n535), .B2(n80), .A(n81), .ZN(n45) );
  NAND2_X1 U505 ( .A1(n9), .A2(n561), .ZN(n12) );
  XNOR2_X1 U506 ( .A(n581), .B(a[4]), .ZN(n542) );
  XOR2_X1 U507 ( .A(n208), .B(n213), .Z(n543) );
  XOR2_X1 U508 ( .A(n543), .B(n206), .Z(n204) );
  NAND2_X1 U509 ( .A1(n215), .A2(n307), .ZN(n544) );
  NAND2_X1 U510 ( .A1(n215), .A2(n210), .ZN(n545) );
  NAND2_X1 U511 ( .A1(n307), .A2(n210), .ZN(n546) );
  NAND3_X1 U512 ( .A1(n544), .A2(n545), .A3(n546), .ZN(n205) );
  NAND2_X1 U513 ( .A1(n208), .A2(n213), .ZN(n547) );
  NAND2_X1 U514 ( .A1(n208), .A2(n206), .ZN(n548) );
  NAND2_X1 U515 ( .A1(n213), .A2(n206), .ZN(n549) );
  NAND3_X1 U516 ( .A1(n547), .A2(n548), .A3(n549), .ZN(n203) );
  INV_X1 U517 ( .A(n19), .ZN(n550) );
  NAND2_X1 U518 ( .A1(n431), .A2(n16), .ZN(n551) );
  NAND2_X1 U519 ( .A1(n431), .A2(n16), .ZN(n552) );
  NAND2_X1 U520 ( .A1(n431), .A2(n16), .ZN(n18) );
  NAND2_X1 U521 ( .A1(n226), .A2(n491), .ZN(n553) );
  NAND2_X1 U522 ( .A1(n226), .A2(n298), .ZN(n554) );
  NAND2_X1 U523 ( .A1(n491), .A2(n298), .ZN(n555) );
  NAND3_X1 U524 ( .A1(n553), .A2(n554), .A3(n555), .ZN(n223) );
  OR2_X1 U525 ( .A1(n6), .A2(n403), .ZN(n556) );
  NAND2_X1 U526 ( .A1(n556), .A2(n557), .ZN(n324) );
  OR2_X1 U527 ( .A1(n29), .A2(n352), .ZN(n558) );
  OR2_X1 U528 ( .A1(n351), .A2(n27), .ZN(n559) );
  NAND2_X1 U529 ( .A1(n558), .A2(n559), .ZN(n277) );
  XNOR2_X1 U530 ( .A(n584), .B(a[6]), .ZN(n560) );
  XNOR2_X1 U531 ( .A(n70), .B(n47), .ZN(product[14]) );
  NAND2_X1 U532 ( .A1(n562), .A2(n69), .ZN(n47) );
  INV_X1 U533 ( .A(n74), .ZN(n72) );
  INV_X1 U534 ( .A(n69), .ZN(n67) );
  NAND2_X1 U535 ( .A1(n73), .A2(n562), .ZN(n64) );
  INV_X1 U536 ( .A(n73), .ZN(n71) );
  NOR2_X1 U537 ( .A1(n514), .A2(n85), .ZN(n80) );
  OAI21_X1 U538 ( .B1(n82), .B2(n86), .A(n83), .ZN(n81) );
  NAND2_X1 U539 ( .A1(n129), .A2(n90), .ZN(n52) );
  INV_X1 U540 ( .A(n89), .ZN(n129) );
  OR2_X1 U541 ( .A1(n152), .A2(n163), .ZN(n562) );
  NAND2_X1 U542 ( .A1(n125), .A2(n76), .ZN(n48) );
  INV_X1 U543 ( .A(n75), .ZN(n125) );
  OAI21_X1 U544 ( .B1(n75), .B2(n79), .A(n76), .ZN(n74) );
  NOR2_X1 U545 ( .A1(n75), .A2(n78), .ZN(n73) );
  XNOR2_X1 U546 ( .A(n84), .B(n50), .ZN(product[11]) );
  NAND2_X1 U547 ( .A1(n127), .A2(n495), .ZN(n50) );
  INV_X1 U548 ( .A(n514), .ZN(n127) );
  NAND2_X1 U549 ( .A1(n152), .A2(n163), .ZN(n69) );
  INV_X1 U550 ( .A(n95), .ZN(n93) );
  OAI21_X1 U551 ( .B1(n113), .B2(n115), .A(n114), .ZN(n112) );
  NAND2_X1 U552 ( .A1(n133), .A2(n106), .ZN(n56) );
  INV_X1 U553 ( .A(n105), .ZN(n133) );
  AOI21_X1 U554 ( .B1(n565), .B2(n120), .A(n117), .ZN(n115) );
  INV_X1 U555 ( .A(n119), .ZN(n117) );
  NAND2_X1 U556 ( .A1(n566), .A2(n103), .ZN(n55) );
  NAND2_X1 U557 ( .A1(n564), .A2(n62), .ZN(n46) );
  AOI21_X1 U558 ( .B1(n530), .B2(n562), .A(n67), .ZN(n65) );
  OAI21_X1 U559 ( .B1(n105), .B2(n107), .A(n106), .ZN(n104) );
  INV_X1 U560 ( .A(n122), .ZN(n120) );
  XNOR2_X1 U561 ( .A(n57), .B(n510), .ZN(product[4]) );
  NAND2_X1 U562 ( .A1(n176), .A2(n185), .ZN(n79) );
  NAND2_X1 U563 ( .A1(n196), .A2(n203), .ZN(n86) );
  NAND2_X1 U564 ( .A1(n186), .A2(n195), .ZN(n83) );
  NAND2_X1 U565 ( .A1(n164), .A2(n175), .ZN(n76) );
  NAND2_X1 U566 ( .A1(n212), .A2(n217), .ZN(n95) );
  OR2_X1 U567 ( .A1(n212), .A2(n217), .ZN(n563) );
  XOR2_X1 U568 ( .A(n58), .B(n115), .Z(product[3]) );
  NAND2_X1 U569 ( .A1(n135), .A2(n114), .ZN(n58) );
  INV_X1 U570 ( .A(n113), .ZN(n135) );
  XNOR2_X1 U571 ( .A(n59), .B(n120), .ZN(product[2]) );
  NAND2_X1 U572 ( .A1(n565), .A2(n119), .ZN(n59) );
  NAND2_X1 U573 ( .A1(n563), .A2(n95), .ZN(n53) );
  NAND2_X1 U574 ( .A1(n131), .A2(n98), .ZN(n54) );
  INV_X1 U575 ( .A(n97), .ZN(n131) );
  NOR2_X1 U576 ( .A1(n234), .A2(n257), .ZN(n113) );
  NAND2_X1 U577 ( .A1(n328), .A2(n314), .ZN(n119) );
  NOR2_X1 U578 ( .A1(n218), .A2(n223), .ZN(n97) );
  NOR2_X1 U579 ( .A1(n228), .A2(n231), .ZN(n105) );
  OR2_X1 U580 ( .A1(n139), .A2(n151), .ZN(n564) );
  OR2_X1 U581 ( .A1(n328), .A2(n314), .ZN(n565) );
  NAND2_X1 U582 ( .A1(n218), .A2(n223), .ZN(n98) );
  NAND2_X1 U583 ( .A1(n228), .A2(n231), .ZN(n106) );
  INV_X1 U584 ( .A(n37), .ZN(n237) );
  OR2_X1 U585 ( .A1(n224), .A2(n227), .ZN(n566) );
  NAND2_X1 U586 ( .A1(n224), .A2(n227), .ZN(n103) );
  INV_X1 U587 ( .A(n41), .ZN(n235) );
  NAND2_X1 U588 ( .A1(n232), .A2(n233), .ZN(n111) );
  OR2_X1 U589 ( .A1(n232), .A2(n233), .ZN(n567) );
  AND2_X1 U590 ( .A1(n492), .A2(n122), .ZN(product[1]) );
  XNOR2_X1 U591 ( .A(n589), .B(a[12]), .ZN(n37) );
  XNOR2_X1 U592 ( .A(n591), .B(a[14]), .ZN(n41) );
  OR2_X1 U593 ( .A1(n574), .A2(n497), .ZN(n392) );
  XNOR2_X1 U594 ( .A(n580), .B(n43), .ZN(n391) );
  OAI22_X1 U595 ( .A1(n39), .A2(n336), .B1(n503), .B2(n335), .ZN(n263) );
  AND2_X1 U596 ( .A1(n574), .A2(n560), .ZN(n288) );
  AND2_X1 U597 ( .A1(n574), .A2(n534), .ZN(n270) );
  XNOR2_X1 U598 ( .A(n583), .B(n43), .ZN(n376) );
  XNOR2_X1 U599 ( .A(n155), .B(n569), .ZN(n139) );
  XNOR2_X1 U600 ( .A(n153), .B(n141), .ZN(n569) );
  XNOR2_X1 U601 ( .A(n157), .B(n570), .ZN(n141) );
  XNOR2_X1 U602 ( .A(n145), .B(n143), .ZN(n570) );
  OAI22_X1 U603 ( .A1(n42), .A2(n594), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U604 ( .A1(n43), .A2(n594), .ZN(n332) );
  XNOR2_X1 U605 ( .A(n499), .B(n43), .ZN(n343) );
  XOR2_X1 U606 ( .A(n587), .B(a[8]), .Z(n429) );
  XNOR2_X1 U607 ( .A(n159), .B(n571), .ZN(n142) );
  XNOR2_X1 U608 ( .A(n315), .B(n261), .ZN(n571) );
  AND2_X1 U609 ( .A1(n574), .A2(n516), .ZN(n300) );
  XNOR2_X1 U610 ( .A(n591), .B(n43), .ZN(n336) );
  AND2_X1 U611 ( .A1(n574), .A2(n247), .ZN(n314) );
  NAND2_X1 U612 ( .A1(n427), .A2(n37), .ZN(n39) );
  XOR2_X1 U613 ( .A(n591), .B(a[12]), .Z(n427) );
  AND2_X1 U614 ( .A1(n574), .A2(n241), .ZN(n278) );
  AND2_X1 U615 ( .A1(n574), .A2(n235), .ZN(n260) );
  OAI22_X1 U616 ( .A1(n39), .A2(n335), .B1(n503), .B2(n334), .ZN(n262) );
  INV_X1 U617 ( .A(n25), .ZN(n588) );
  XNOR2_X1 U618 ( .A(n502), .B(n43), .ZN(n352) );
  NAND2_X1 U619 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U620 ( .A(n593), .B(a[14]), .Z(n426) );
  XNOR2_X1 U621 ( .A(n505), .B(n43), .ZN(n363) );
  OAI22_X1 U622 ( .A1(n39), .A2(n592), .B1(n337), .B2(n503), .ZN(n252) );
  OR2_X1 U623 ( .A1(n43), .A2(n592), .ZN(n337) );
  AND2_X1 U624 ( .A1(n574), .A2(n237), .ZN(n264) );
  AND2_X1 U625 ( .A1(n574), .A2(n249), .ZN(product[0]) );
  OR2_X1 U626 ( .A1(n43), .A2(n590), .ZN(n344) );
  OR2_X1 U627 ( .A1(n43), .A2(n588), .ZN(n353) );
  OR2_X1 U628 ( .A1(n43), .A2(n586), .ZN(n364) );
  OR2_X1 U629 ( .A1(n43), .A2(n493), .ZN(n377) );
  XNOR2_X1 U630 ( .A(n505), .B(b[9]), .ZN(n354) );
  OAI22_X1 U631 ( .A1(n39), .A2(n334), .B1(n503), .B2(n333), .ZN(n261) );
  XNOR2_X1 U632 ( .A(n591), .B(n422), .ZN(n333) );
  XNOR2_X1 U633 ( .A(n583), .B(b[11]), .ZN(n365) );
  XNOR2_X1 U634 ( .A(n591), .B(n424), .ZN(n335) );
  XNOR2_X1 U635 ( .A(n591), .B(n423), .ZN(n334) );
  OAI22_X1 U636 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U637 ( .A(n593), .B(n424), .ZN(n330) );
  XNOR2_X1 U638 ( .A(n593), .B(n43), .ZN(n331) );
  XNOR2_X1 U639 ( .A(n502), .B(n418), .ZN(n345) );
  XNOR2_X1 U640 ( .A(n589), .B(n424), .ZN(n342) );
  XNOR2_X1 U641 ( .A(n500), .B(n424), .ZN(n362) );
  XNOR2_X1 U642 ( .A(n587), .B(n424), .ZN(n351) );
  XNOR2_X1 U643 ( .A(n579), .B(n424), .ZN(n390) );
  XNOR2_X1 U644 ( .A(n582), .B(n424), .ZN(n375) );
  XNOR2_X1 U645 ( .A(n499), .B(n420), .ZN(n338) );
  XNOR2_X1 U646 ( .A(n580), .B(b[13]), .ZN(n378) );
  XNOR2_X1 U647 ( .A(n589), .B(n423), .ZN(n341) );
  XNOR2_X1 U648 ( .A(n499), .B(n422), .ZN(n340) );
  XNOR2_X1 U649 ( .A(n499), .B(n421), .ZN(n339) );
  XNOR2_X1 U650 ( .A(n579), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U651 ( .A(n579), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U652 ( .A(n580), .B(n418), .ZN(n384) );
  XNOR2_X1 U653 ( .A(n580), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U654 ( .A(n580), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U655 ( .A(n580), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U656 ( .A(n580), .B(n419), .ZN(n385) );
  XNOR2_X1 U657 ( .A(n579), .B(n422), .ZN(n388) );
  XNOR2_X1 U658 ( .A(n579), .B(n423), .ZN(n389) );
  XNOR2_X1 U659 ( .A(n587), .B(n423), .ZN(n350) );
  XNOR2_X1 U660 ( .A(n505), .B(n423), .ZN(n361) );
  XNOR2_X1 U661 ( .A(n505), .B(n422), .ZN(n360) );
  XNOR2_X1 U662 ( .A(n582), .B(n423), .ZN(n374) );
  XNOR2_X1 U663 ( .A(n502), .B(n422), .ZN(n349) );
  XNOR2_X1 U664 ( .A(n582), .B(n422), .ZN(n373) );
  XNOR2_X1 U665 ( .A(n583), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U666 ( .A(n583), .B(n418), .ZN(n369) );
  XNOR2_X1 U667 ( .A(n583), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U668 ( .A(n583), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U669 ( .A(n576), .B(b[11]), .ZN(n397) );
  XNOR2_X1 U670 ( .A(n576), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U671 ( .A(n496), .B(b[14]), .ZN(n394) );
  XNOR2_X1 U672 ( .A(n505), .B(n421), .ZN(n359) );
  XNOR2_X1 U673 ( .A(n500), .B(n420), .ZN(n358) );
  XNOR2_X1 U674 ( .A(n580), .B(n421), .ZN(n387) );
  XNOR2_X1 U675 ( .A(n582), .B(n420), .ZN(n371) );
  XNOR2_X1 U676 ( .A(n582), .B(n421), .ZN(n372) );
  XNOR2_X1 U677 ( .A(n587), .B(n421), .ZN(n348) );
  XNOR2_X1 U678 ( .A(n502), .B(n420), .ZN(n347) );
  XNOR2_X1 U679 ( .A(n580), .B(n420), .ZN(n386) );
  XNOR2_X1 U680 ( .A(n582), .B(n419), .ZN(n370) );
  XNOR2_X1 U681 ( .A(n505), .B(n419), .ZN(n357) );
  XNOR2_X1 U682 ( .A(n502), .B(n419), .ZN(n346) );
  XNOR2_X1 U683 ( .A(n500), .B(n418), .ZN(n356) );
  XNOR2_X1 U684 ( .A(n500), .B(b[8]), .ZN(n355) );
  XNOR2_X1 U685 ( .A(n496), .B(b[15]), .ZN(n393) );
  BUF_X1 U686 ( .A(n43), .Z(n574) );
  OAI22_X1 U687 ( .A1(n537), .A2(n395), .B1(n394), .B2(n528), .ZN(n316) );
  OAI22_X1 U688 ( .A1(n537), .A2(n400), .B1(n399), .B2(n528), .ZN(n321) );
  OAI22_X1 U689 ( .A1(n537), .A2(n394), .B1(n393), .B2(n528), .ZN(n315) );
  OAI22_X1 U690 ( .A1(n537), .A2(n401), .B1(n400), .B2(n528), .ZN(n322) );
  OAI22_X1 U691 ( .A1(n537), .A2(n397), .B1(n396), .B2(n528), .ZN(n318) );
  OAI22_X1 U692 ( .A1(n537), .A2(n396), .B1(n395), .B2(n528), .ZN(n317) );
  OAI22_X1 U693 ( .A1(n398), .A2(n537), .B1(n397), .B2(n575), .ZN(n319) );
  OAI22_X1 U694 ( .A1(n6), .A2(n406), .B1(n405), .B2(n528), .ZN(n327) );
  OAI22_X1 U695 ( .A1(n6), .A2(n405), .B1(n404), .B2(n575), .ZN(n326) );
  OAI22_X1 U696 ( .A1(n6), .A2(n404), .B1(n403), .B2(n575), .ZN(n325) );
  OAI22_X1 U697 ( .A1(n399), .A2(n537), .B1(n398), .B2(n575), .ZN(n320) );
  OAI22_X1 U698 ( .A1(n537), .A2(n402), .B1(n401), .B2(n528), .ZN(n323) );
  OAI22_X1 U699 ( .A1(n537), .A2(n408), .B1(n407), .B2(n528), .ZN(n329) );
  OAI22_X1 U700 ( .A1(n537), .A2(n407), .B1(n406), .B2(n528), .ZN(n328) );
  OAI22_X1 U701 ( .A1(n34), .A2(n339), .B1(n338), .B2(n32), .ZN(n265) );
  OAI22_X1 U702 ( .A1(n34), .A2(n340), .B1(n339), .B2(n32), .ZN(n266) );
  OAI22_X1 U703 ( .A1(n34), .A2(n341), .B1(n340), .B2(n32), .ZN(n267) );
  OAI22_X1 U704 ( .A1(n34), .A2(n342), .B1(n341), .B2(n32), .ZN(n268) );
  OAI22_X1 U705 ( .A1(n34), .A2(n343), .B1(n342), .B2(n32), .ZN(n269) );
  OAI22_X1 U706 ( .A1(n34), .A2(n590), .B1(n344), .B2(n32), .ZN(n253) );
  INV_X1 U707 ( .A(n496), .ZN(n572) );
  INV_X1 U708 ( .A(n19), .ZN(n586) );
  INV_X1 U709 ( .A(n1), .ZN(n578) );
  OAI21_X1 U710 ( .B1(n536), .B2(n97), .A(n98), .ZN(n573) );
  OAI21_X1 U711 ( .B1(n99), .B2(n97), .A(n98), .ZN(n96) );
  NAND2_X1 U712 ( .A1(n204), .A2(n211), .ZN(n90) );
  NOR2_X1 U713 ( .A1(n204), .A2(n211), .ZN(n89) );
  OAI22_X1 U714 ( .A1(n494), .A2(n350), .B1(n349), .B2(n498), .ZN(n275) );
  OAI22_X1 U715 ( .A1(n494), .A2(n346), .B1(n345), .B2(n498), .ZN(n271) );
  OAI22_X1 U716 ( .A1(n494), .A2(n347), .B1(n346), .B2(n498), .ZN(n272) );
  OAI22_X1 U717 ( .A1(n494), .A2(n348), .B1(n347), .B2(n498), .ZN(n273) );
  OAI22_X1 U718 ( .A1(n29), .A2(n349), .B1(n348), .B2(n498), .ZN(n274) );
  OAI22_X1 U719 ( .A1(n494), .A2(n351), .B1(n350), .B2(n498), .ZN(n276) );
  OAI22_X1 U720 ( .A1(n29), .A2(n588), .B1(n353), .B2(n27), .ZN(n254) );
  INV_X1 U721 ( .A(n27), .ZN(n241) );
  XNOR2_X1 U722 ( .A(n77), .B(n48), .ZN(product[13]) );
  NAND2_X1 U723 ( .A1(n567), .A2(n111), .ZN(n57) );
  OR2_X1 U724 ( .A1(n43), .A2(n572), .ZN(n409) );
  XNOR2_X1 U725 ( .A(n63), .B(n46), .ZN(product[15]) );
  INV_X1 U726 ( .A(n7), .ZN(n581) );
  XOR2_X1 U727 ( .A(n536), .B(n54), .Z(product[7]) );
  XNOR2_X1 U728 ( .A(n573), .B(n53), .ZN(product[8]) );
  INV_X1 U729 ( .A(n13), .ZN(n584) );
  AOI21_X1 U730 ( .B1(n566), .B2(n104), .A(n101), .ZN(n99) );
  INV_X1 U731 ( .A(n103), .ZN(n101) );
  OAI22_X1 U732 ( .A1(n23), .A2(n356), .B1(n355), .B2(n21), .ZN(n280) );
  OAI22_X1 U733 ( .A1(n23), .A2(n358), .B1(n357), .B2(n21), .ZN(n282) );
  OAI22_X1 U734 ( .A1(n23), .A2(n362), .B1(n21), .B2(n361), .ZN(n286) );
  OAI22_X1 U735 ( .A1(n23), .A2(n360), .B1(n21), .B2(n359), .ZN(n284) );
  OAI22_X1 U736 ( .A1(n23), .A2(n361), .B1(n21), .B2(n360), .ZN(n285) );
  OAI22_X1 U737 ( .A1(n23), .A2(n586), .B1(n21), .B2(n364), .ZN(n255) );
  OAI22_X1 U738 ( .A1(n23), .A2(n355), .B1(n354), .B2(n21), .ZN(n279) );
  OAI22_X1 U739 ( .A1(n23), .A2(n357), .B1(n21), .B2(n356), .ZN(n281) );
  OAI22_X1 U740 ( .A1(n23), .A2(n363), .B1(n362), .B2(n21), .ZN(n287) );
  OAI22_X1 U741 ( .A1(n23), .A2(n359), .B1(n21), .B2(n358), .ZN(n283) );
  OAI21_X1 U742 ( .B1(n87), .B2(n85), .A(n507), .ZN(n84) );
  INV_X1 U743 ( .A(n88), .ZN(n87) );
  OAI21_X1 U744 ( .B1(n91), .B2(n89), .A(n90), .ZN(n88) );
  XNOR2_X1 U745 ( .A(n520), .B(n55), .ZN(product[6]) );
  NAND2_X1 U746 ( .A1(n151), .A2(n139), .ZN(n62) );
  OAI22_X1 U747 ( .A1(n552), .A2(n370), .B1(n369), .B2(n515), .ZN(n293) );
  OAI22_X1 U748 ( .A1(n551), .A2(n367), .B1(n366), .B2(n515), .ZN(n290) );
  OAI22_X1 U749 ( .A1(n552), .A2(n375), .B1(n374), .B2(n515), .ZN(n298) );
  OAI22_X1 U750 ( .A1(n551), .A2(n368), .B1(n367), .B2(n515), .ZN(n291) );
  OAI22_X1 U751 ( .A1(n552), .A2(n372), .B1(n371), .B2(n515), .ZN(n295) );
  OAI22_X1 U752 ( .A1(n552), .A2(n373), .B1(n372), .B2(n515), .ZN(n296) );
  OAI22_X1 U753 ( .A1(n551), .A2(n369), .B1(n368), .B2(n515), .ZN(n292) );
  OAI22_X1 U754 ( .A1(n18), .A2(n371), .B1(n370), .B2(n515), .ZN(n294) );
  OAI22_X1 U755 ( .A1(n18), .A2(n374), .B1(n373), .B2(n515), .ZN(n297) );
  OAI22_X1 U756 ( .A1(n552), .A2(n493), .B1(n377), .B2(n515), .ZN(n256) );
  OAI22_X1 U757 ( .A1(n551), .A2(n376), .B1(n375), .B2(n515), .ZN(n299) );
  OAI22_X1 U758 ( .A1(n551), .A2(n366), .B1(n365), .B2(n515), .ZN(n289) );
  OAI21_X1 U759 ( .B1(n64), .B2(n538), .A(n65), .ZN(n63) );
  OAI21_X1 U760 ( .B1(n538), .B2(n78), .A(n79), .ZN(n77) );
  OAI21_X1 U761 ( .B1(n45), .B2(n71), .A(n72), .ZN(n70) );
  XNOR2_X1 U762 ( .A(n576), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U763 ( .A(n576), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U764 ( .A(n496), .B(n418), .ZN(n401) );
  XNOR2_X1 U765 ( .A(n496), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U766 ( .A(n496), .B(n421), .ZN(n404) );
  XNOR2_X1 U767 ( .A(n496), .B(n422), .ZN(n405) );
  XNOR2_X1 U768 ( .A(n576), .B(n43), .ZN(n408) );
  XNOR2_X1 U769 ( .A(n576), .B(n419), .ZN(n402) );
  XNOR2_X1 U770 ( .A(n496), .B(n420), .ZN(n403) );
  XNOR2_X1 U771 ( .A(n576), .B(n424), .ZN(n407) );
  XNOR2_X1 U772 ( .A(n576), .B(n423), .ZN(n406) );
  XOR2_X1 U773 ( .A(n532), .B(n52), .Z(product[9]) );
  XOR2_X1 U774 ( .A(n56), .B(n107), .Z(product[5]) );
  NAND2_X1 U775 ( .A1(n329), .A2(n258), .ZN(n122) );
  INV_X1 U776 ( .A(n111), .ZN(n109) );
  OAI22_X1 U777 ( .A1(n6), .A2(n572), .B1(n409), .B2(n528), .ZN(n258) );
  OAI22_X1 U778 ( .A1(n540), .A2(n379), .B1(n378), .B2(n511), .ZN(n301) );
  OAI22_X1 U779 ( .A1(n541), .A2(n380), .B1(n379), .B2(n512), .ZN(n302) );
  OAI22_X1 U780 ( .A1(n540), .A2(n385), .B1(n384), .B2(n512), .ZN(n307) );
  OAI22_X1 U781 ( .A1(n540), .A2(n382), .B1(n381), .B2(n512), .ZN(n304) );
  OAI22_X1 U782 ( .A1(n541), .A2(n381), .B1(n380), .B2(n511), .ZN(n303) );
  NAND2_X1 U783 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U784 ( .A1(n541), .A2(n383), .B1(n382), .B2(n512), .ZN(n305) );
  OAI22_X1 U785 ( .A1(n540), .A2(n384), .B1(n383), .B2(n511), .ZN(n306) );
  OAI22_X1 U786 ( .A1(n541), .A2(n386), .B1(n385), .B2(n512), .ZN(n308) );
  OAI22_X1 U787 ( .A1(n540), .A2(n387), .B1(n386), .B2(n511), .ZN(n309) );
  OAI22_X1 U788 ( .A1(n541), .A2(n497), .B1(n392), .B2(n511), .ZN(n257) );
  OAI22_X1 U789 ( .A1(n539), .A2(n389), .B1(n388), .B2(n512), .ZN(n311) );
  OAI22_X1 U790 ( .A1(n540), .A2(n388), .B1(n387), .B2(n512), .ZN(n310) );
  OAI22_X1 U791 ( .A1(n539), .A2(n390), .B1(n389), .B2(n511), .ZN(n312) );
  INV_X1 U792 ( .A(n511), .ZN(n247) );
  OAI22_X1 U793 ( .A1(n541), .A2(n391), .B1(n390), .B2(n512), .ZN(n313) );
  INV_X1 U794 ( .A(n584), .ZN(n583) );
  INV_X1 U795 ( .A(n31), .ZN(n590) );
  INV_X1 U796 ( .A(n592), .ZN(n591) );
  INV_X1 U797 ( .A(n36), .ZN(n592) );
  INV_X1 U798 ( .A(n594), .ZN(n593) );
  INV_X1 U799 ( .A(n40), .ZN(n594) );
  XOR2_X1 U800 ( .A(n259), .B(n251), .Z(n148) );
  XOR2_X1 U801 ( .A(n289), .B(n279), .Z(n146) );
  XOR2_X1 U802 ( .A(n149), .B(n147), .Z(n144) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_11_DW01_add_2 ( A, B, CI, SUM, 
        CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n7, n8, n9, n10, n11, n12, n13, n14, n15, n18, n19,
         n20, n21, n23, n25, n26, n27, n28, n30, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n48, n49, n51, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n71, n72, n73, n74,
         n75, n77, n79, n80, n81, n82, n83, n85, n87, n88, n90, n93, n94, n98,
         n99, n100, n102, n104, n161, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179;

  AOI21_X1 U126 ( .B1(n56), .B2(n64), .A(n57), .ZN(n161) );
  OR2_X2 U127 ( .A1(A[10]), .A2(B[10]), .ZN(n177) );
  NOR2_X1 U128 ( .A1(A[11]), .A2(B[11]), .ZN(n39) );
  AND2_X1 U129 ( .A1(n173), .A2(n90), .ZN(SUM[0]) );
  OR2_X1 U130 ( .A1(A[15]), .A2(B[15]), .ZN(n163) );
  XNOR2_X1 U131 ( .A(n49), .B(n164), .ZN(SUM[10]) );
  AND2_X1 U132 ( .A1(n177), .A2(n48), .ZN(n164) );
  INV_X1 U133 ( .A(n171), .ZN(n48) );
  OR2_X1 U134 ( .A1(A[11]), .A2(B[11]), .ZN(n165) );
  XNOR2_X1 U135 ( .A(n41), .B(n166), .ZN(SUM[11]) );
  AND2_X1 U136 ( .A1(n165), .A2(n40), .ZN(n166) );
  BUF_X1 U137 ( .A(n37), .Z(n167) );
  BUF_X1 U138 ( .A(n170), .Z(n168) );
  NOR2_X1 U139 ( .A1(A[8]), .A2(B[8]), .ZN(n169) );
  AOI21_X2 U140 ( .B1(n42), .B2(n34), .A(n35), .ZN(n172) );
  NOR2_X1 U141 ( .A1(A[12]), .A2(B[12]), .ZN(n170) );
  NOR2_X1 U142 ( .A1(A[12]), .A2(B[12]), .ZN(n36) );
  AND2_X1 U143 ( .A1(A[10]), .A2(B[10]), .ZN(n171) );
  OR2_X1 U144 ( .A1(A[0]), .A2(B[0]), .ZN(n173) );
  INV_X1 U145 ( .A(n161), .ZN(n54) );
  AOI21_X1 U146 ( .B1(n178), .B2(n72), .A(n69), .ZN(n67) );
  INV_X1 U147 ( .A(n71), .ZN(n69) );
  AOI21_X1 U148 ( .B1(n176), .B2(n80), .A(n77), .ZN(n75) );
  AOI21_X1 U149 ( .B1(n175), .B2(n88), .A(n85), .ZN(n83) );
  INV_X1 U150 ( .A(n87), .ZN(n85) );
  OAI21_X1 U151 ( .B1(n83), .B2(n81), .A(n82), .ZN(n80) );
  INV_X1 U152 ( .A(n28), .ZN(n30) );
  OAI21_X1 U153 ( .B1(n75), .B2(n73), .A(n74), .ZN(n72) );
  AOI21_X1 U154 ( .B1(n54), .B2(n174), .A(n51), .ZN(n49) );
  INV_X1 U155 ( .A(n90), .ZN(n88) );
  OAI21_X1 U156 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  INV_X1 U157 ( .A(n53), .ZN(n51) );
  INV_X1 U158 ( .A(n27), .ZN(n93) );
  NAND2_X1 U159 ( .A1(n102), .A2(n74), .ZN(n12) );
  INV_X1 U160 ( .A(n73), .ZN(n102) );
  NAND2_X1 U161 ( .A1(n174), .A2(n53), .ZN(n7) );
  NAND2_X1 U162 ( .A1(n176), .A2(n79), .ZN(n13) );
  NAND2_X1 U163 ( .A1(n99), .A2(n62), .ZN(n9) );
  INV_X1 U164 ( .A(n61), .ZN(n99) );
  NAND2_X1 U165 ( .A1(n104), .A2(n82), .ZN(n14) );
  INV_X1 U166 ( .A(n81), .ZN(n104) );
  NAND2_X1 U167 ( .A1(n98), .A2(n59), .ZN(n8) );
  INV_X1 U168 ( .A(n169), .ZN(n98) );
  NAND2_X1 U169 ( .A1(n100), .A2(n66), .ZN(n10) );
  INV_X1 U170 ( .A(n65), .ZN(n100) );
  NAND2_X1 U171 ( .A1(n178), .A2(n71), .ZN(n11) );
  NAND2_X1 U172 ( .A1(n175), .A2(n87), .ZN(n15) );
  INV_X1 U173 ( .A(n25), .ZN(n23) );
  NAND2_X1 U174 ( .A1(n94), .A2(n167), .ZN(n4) );
  XNOR2_X1 U175 ( .A(n54), .B(n7), .ZN(SUM[9]) );
  XOR2_X1 U176 ( .A(n63), .B(n9), .Z(SUM[7]) );
  XOR2_X1 U177 ( .A(n12), .B(n75), .Z(SUM[4]) );
  XNOR2_X1 U178 ( .A(n13), .B(n80), .ZN(SUM[3]) );
  XNOR2_X1 U179 ( .A(n15), .B(n88), .ZN(SUM[1]) );
  NOR2_X1 U180 ( .A1(A[7]), .A2(B[7]), .ZN(n61) );
  OR2_X1 U181 ( .A1(A[9]), .A2(B[9]), .ZN(n174) );
  NOR2_X1 U182 ( .A1(A[2]), .A2(B[2]), .ZN(n81) );
  NOR2_X1 U183 ( .A1(A[4]), .A2(B[4]), .ZN(n73) );
  NAND2_X1 U184 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  NAND2_X1 U185 ( .A1(A[11]), .A2(B[11]), .ZN(n40) );
  OR2_X1 U186 ( .A1(A[1]), .A2(B[1]), .ZN(n175) );
  OR2_X1 U187 ( .A1(A[3]), .A2(B[3]), .ZN(n176) );
  NOR2_X1 U188 ( .A1(A[8]), .A2(B[8]), .ZN(n58) );
  NAND2_X1 U189 ( .A1(A[12]), .A2(B[12]), .ZN(n37) );
  XNOR2_X1 U190 ( .A(n60), .B(n8), .ZN(SUM[8]) );
  NOR2_X1 U191 ( .A1(A[6]), .A2(B[6]), .ZN(n65) );
  NAND2_X1 U192 ( .A1(A[7]), .A2(B[7]), .ZN(n62) );
  OR2_X1 U193 ( .A1(A[5]), .A2(B[5]), .ZN(n178) );
  NAND2_X1 U194 ( .A1(A[2]), .A2(B[2]), .ZN(n82) );
  NAND2_X1 U195 ( .A1(A[4]), .A2(B[4]), .ZN(n74) );
  NAND2_X1 U196 ( .A1(A[15]), .A2(B[15]), .ZN(n18) );
  NAND2_X1 U197 ( .A1(A[5]), .A2(B[5]), .ZN(n71) );
  NAND2_X1 U198 ( .A1(A[1]), .A2(B[1]), .ZN(n87) );
  NAND2_X1 U199 ( .A1(A[0]), .A2(B[0]), .ZN(n90) );
  NAND2_X1 U200 ( .A1(A[6]), .A2(B[6]), .ZN(n66) );
  NAND2_X1 U201 ( .A1(A[8]), .A2(B[8]), .ZN(n59) );
  XOR2_X1 U202 ( .A(n67), .B(n10), .Z(SUM[6]) );
  XNOR2_X1 U203 ( .A(n11), .B(n72), .ZN(SUM[5]) );
  XOR2_X1 U204 ( .A(n14), .B(n83), .Z(SUM[2]) );
  OR2_X1 U205 ( .A1(A[14]), .A2(B[14]), .ZN(n179) );
  NAND2_X1 U206 ( .A1(n93), .A2(n28), .ZN(n3) );
  OAI21_X1 U207 ( .B1(n41), .B2(n39), .A(n40), .ZN(n38) );
  INV_X1 U208 ( .A(n42), .ZN(n41) );
  NAND2_X1 U209 ( .A1(A[9]), .A2(B[9]), .ZN(n53) );
  NOR2_X1 U210 ( .A1(A[13]), .A2(B[13]), .ZN(n27) );
  NAND2_X1 U211 ( .A1(n163), .A2(n18), .ZN(n1) );
  NAND2_X1 U212 ( .A1(A[14]), .A2(B[14]), .ZN(n25) );
  OAI21_X1 U213 ( .B1(n58), .B2(n62), .A(n59), .ZN(n57) );
  NOR2_X1 U214 ( .A1(n169), .A2(n61), .ZN(n56) );
  INV_X1 U215 ( .A(n168), .ZN(n94) );
  NOR2_X1 U216 ( .A1(n170), .A2(n39), .ZN(n34) );
  OAI21_X1 U217 ( .B1(n36), .B2(n40), .A(n37), .ZN(n35) );
  NAND2_X1 U218 ( .A1(A[3]), .A2(B[3]), .ZN(n79) );
  INV_X1 U219 ( .A(n79), .ZN(n77) );
  OAI21_X1 U220 ( .B1(n67), .B2(n65), .A(n66), .ZN(n64) );
  AOI21_X1 U221 ( .B1(n56), .B2(n64), .A(n57), .ZN(n55) );
  INV_X1 U222 ( .A(n64), .ZN(n63) );
  NAND2_X1 U223 ( .A1(n179), .A2(n25), .ZN(n2) );
  NAND2_X1 U224 ( .A1(n179), .A2(n93), .ZN(n20) );
  AOI21_X1 U225 ( .B1(n179), .B2(n30), .A(n23), .ZN(n21) );
  XNOR2_X1 U226 ( .A(n26), .B(n2), .ZN(SUM[14]) );
  XNOR2_X1 U227 ( .A(n19), .B(n1), .ZN(SUM[15]) );
  NAND2_X1 U228 ( .A1(n177), .A2(n174), .ZN(n43) );
  AOI21_X1 U229 ( .B1(n177), .B2(n51), .A(n171), .ZN(n44) );
  XNOR2_X1 U230 ( .A(n38), .B(n4), .ZN(SUM[12]) );
  XOR2_X1 U231 ( .A(n172), .B(n3), .Z(SUM[13]) );
  OAI21_X1 U232 ( .B1(n172), .B2(n27), .A(n28), .ZN(n26) );
  OAI21_X1 U233 ( .B1(n20), .B2(n172), .A(n21), .ZN(n19) );
  OAI21_X1 U234 ( .B1(n43), .B2(n55), .A(n44), .ZN(n42) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_11 ( clk, clear_acc, 
        data_out_x, data_out, data_out_w, data_out_b, wr_en_y, m_valid, 
        m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [3:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N27, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, n1, n2, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n87, n104, n113, n114, n115, n116, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n21), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n227), .CK(clk), .Q(n26) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n228), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n229), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n230), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n231), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n232), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n233), .CK(clk), .Q(n34) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n234), .CK(clk), .Q(n35) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n235), .CK(clk), .Q(n36) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n236), .CK(clk), .Q(n37) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n237), .CK(clk), .Q(n38) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n238), .CK(clk), .Q(n39) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n239), .CK(clk), .Q(n40) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n240), .CK(clk), .Q(n41) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n241), .CK(clk), .Q(n42) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n242), .CK(clk), .Q(n44) );
  DFF_X1 \f_reg[7]  ( .D(n84), .CK(clk), .Q(f[7]), .QN(n219) );
  DFF_X1 \f_reg[8]  ( .D(n83), .CK(clk), .Q(f[8]), .QN(n220) );
  DFF_X1 \f_reg[9]  ( .D(n82), .CK(clk), .Q(f[9]), .QN(n221) );
  DFF_X1 \f_reg[10]  ( .D(n81), .CK(clk), .Q(n53), .QN(n222) );
  DFF_X1 \f_reg[11]  ( .D(n80), .CK(clk), .Q(n51), .QN(n223) );
  DFF_X1 \f_reg[12]  ( .D(n4), .CK(clk), .Q(n50), .QN(n224) );
  DFF_X1 \f_reg[13]  ( .D(n2), .CK(clk), .Q(n49), .QN(n225) );
  DFF_X1 \f_reg[14]  ( .D(n8), .CK(clk), .Q(n48), .QN(n226) );
  DFF_X1 \f_reg[15]  ( .D(n79), .CK(clk), .Q(f[15]), .QN(n77) );
  DFF_X1 \data_out_reg[15]  ( .D(n168), .CK(clk), .Q(data_out[15]), .QN(n199)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n169), .CK(clk), .Q(data_out[14]), .QN(n198)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n170), .CK(clk), .Q(data_out[13]), .QN(n197)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n171), .CK(clk), .Q(data_out[12]), .QN(n196)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n172), .CK(clk), .Q(data_out[11]), .QN(n195)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n173), .CK(clk), .Q(data_out[10]), .QN(n194)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n174), .CK(clk), .Q(data_out[9]), .QN(n193) );
  DFF_X1 \data_out_reg[8]  ( .D(n175), .CK(clk), .Q(data_out[8]), .QN(n192) );
  DFF_X1 \data_out_reg[7]  ( .D(n176), .CK(clk), .Q(data_out[7]), .QN(n191) );
  DFF_X1 \data_out_reg[6]  ( .D(n177), .CK(clk), .Q(data_out[6]), .QN(n190) );
  DFF_X1 \data_out_reg[5]  ( .D(n178), .CK(clk), .Q(data_out[5]), .QN(n189) );
  DFF_X1 \data_out_reg[4]  ( .D(n179), .CK(clk), .Q(data_out[4]), .QN(n188) );
  DFF_X1 \data_out_reg[3]  ( .D(n180), .CK(clk), .Q(data_out[3]), .QN(n187) );
  DFF_X1 \data_out_reg[2]  ( .D(n181), .CK(clk), .Q(data_out[2]), .QN(n186) );
  DFF_X1 \data_out_reg[1]  ( .D(n182), .CK(clk), .Q(data_out[1]), .QN(n185) );
  DFF_X1 \data_out_reg[0]  ( .D(n183), .CK(clk), .Q(data_out[0]), .QN(n184) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_11_DW_mult_tc_1 mult_960 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_11_DW01_add_2 add_961 ( .A({n206, 
        n205, n204, n203, n202, n201, n215, n214, n213, n212, n211, n210, n209, 
        n208, n207, n200}), .B({f[15], n48, n49, n50, n51, n53, f[9:3], n61, 
        n63, n65}), .CI(1'b0), .SUM(adder) );
  DFF_X1 \f_reg[2]  ( .D(n114), .CK(clk), .Q(n61), .QN(n218) );
  DFF_X1 \f_reg[3]  ( .D(n113), .CK(clk), .Q(f[3]), .QN(n69) );
  DFF_X1 \f_reg[1]  ( .D(n115), .CK(clk), .Q(n63), .QN(n217) );
  DFF_X1 \f_reg[0]  ( .D(n116), .CK(clk), .Q(n65), .QN(n216) );
  DFF_X1 \f_reg[4]  ( .D(n104), .CK(clk), .Q(f[4]), .QN(n70) );
  DFF_X1 \f_reg[5]  ( .D(n87), .CK(clk), .Q(f[5]), .QN(n71) );
  DFF_X1 \f_reg[6]  ( .D(n85), .CK(clk), .Q(f[6]), .QN(n72) );
  DFF_X2 delay_reg ( .D(N27), .CK(clk), .Q(n1), .QN(n243) );
  AND2_X2 U3 ( .A1(n47), .A2(n22), .ZN(n19) );
  MUX2_X2 U4 ( .A(N41), .B(n29), .S(n1), .Z(n203) );
  MUX2_X2 U5 ( .A(n32), .B(N40), .S(n243), .Z(n202) );
  NAND3_X1 U6 ( .A1(n6), .A2(n5), .A3(n7), .ZN(n2) );
  NAND3_X1 U8 ( .A1(n11), .A2(n10), .A3(n12), .ZN(n4) );
  MUX2_X2 U9 ( .A(n35), .B(N37), .S(n243), .Z(n214) );
  NAND2_X1 U10 ( .A1(data_out_b[13]), .A2(n21), .ZN(n5) );
  NAND2_X1 U11 ( .A1(adder[13]), .A2(n19), .ZN(n6) );
  NAND2_X1 U12 ( .A1(n67), .A2(n49), .ZN(n7) );
  NAND3_X1 U13 ( .A1(n14), .A2(n13), .A3(n15), .ZN(n8) );
  AND2_X1 U14 ( .A1(n18), .A2(n16), .ZN(n9) );
  NAND2_X1 U15 ( .A1(n17), .A2(n9), .ZN(n79) );
  NAND2_X1 U16 ( .A1(data_out_b[12]), .A2(n21), .ZN(n10) );
  NAND2_X1 U17 ( .A1(adder[12]), .A2(n19), .ZN(n11) );
  NAND2_X1 U18 ( .A1(n67), .A2(n50), .ZN(n12) );
  NAND2_X1 U19 ( .A1(data_out_b[14]), .A2(n21), .ZN(n13) );
  NAND2_X1 U20 ( .A1(adder[14]), .A2(n19), .ZN(n14) );
  NAND2_X1 U21 ( .A1(n67), .A2(n48), .ZN(n15) );
  NAND2_X1 U22 ( .A1(data_out_b[15]), .A2(n21), .ZN(n16) );
  NAND2_X1 U23 ( .A1(adder[15]), .A2(n19), .ZN(n17) );
  NAND2_X1 U24 ( .A1(n67), .A2(f[15]), .ZN(n18) );
  INV_X2 U25 ( .A(n47), .ZN(n67) );
  INV_X1 U26 ( .A(n22), .ZN(n21) );
  INV_X1 U27 ( .A(clear_acc), .ZN(n22) );
  NAND2_X1 U28 ( .A1(n20), .A2(N27), .ZN(n245) );
  OAI22_X1 U29 ( .A1(n187), .A2(n245), .B1(n69), .B2(n244), .ZN(n180) );
  OAI22_X1 U30 ( .A1(n188), .A2(n245), .B1(n70), .B2(n244), .ZN(n179) );
  OAI22_X1 U31 ( .A1(n189), .A2(n245), .B1(n71), .B2(n244), .ZN(n178) );
  OAI22_X1 U32 ( .A1(n190), .A2(n245), .B1(n72), .B2(n244), .ZN(n177) );
  OAI22_X1 U33 ( .A1(n191), .A2(n245), .B1(n219), .B2(n244), .ZN(n176) );
  OAI22_X1 U34 ( .A1(n192), .A2(n245), .B1(n220), .B2(n244), .ZN(n175) );
  OAI22_X1 U35 ( .A1(n193), .A2(n245), .B1(n221), .B2(n244), .ZN(n174) );
  INV_X1 U36 ( .A(n25), .ZN(n43) );
  INV_X1 U37 ( .A(wr_en_y), .ZN(n20) );
  AND2_X1 U38 ( .A1(sel[0]), .A2(sel[1]), .ZN(n24) );
  INV_X1 U39 ( .A(m_ready), .ZN(n23) );
  NAND2_X1 U40 ( .A1(m_valid), .A2(n23), .ZN(n45) );
  OAI211_X1 U41 ( .C1(sel[2]), .C2(n24), .A(sel[3]), .B(n45), .ZN(N27) );
  NAND2_X1 U42 ( .A1(clear_acc_delay), .A2(n243), .ZN(n25) );
  MUX2_X1 U43 ( .A(n26), .B(N44), .S(n43), .Z(n227) );
  MUX2_X1 U44 ( .A(n26), .B(N44), .S(n243), .Z(n206) );
  MUX2_X1 U45 ( .A(n27), .B(N43), .S(n43), .Z(n228) );
  MUX2_X1 U46 ( .A(n27), .B(N43), .S(n243), .Z(n205) );
  MUX2_X1 U47 ( .A(n28), .B(N42), .S(n43), .Z(n229) );
  MUX2_X1 U48 ( .A(n28), .B(N42), .S(n243), .Z(n204) );
  MUX2_X1 U49 ( .A(n29), .B(N41), .S(n43), .Z(n230) );
  MUX2_X1 U50 ( .A(n32), .B(N40), .S(n43), .Z(n231) );
  MUX2_X1 U51 ( .A(n33), .B(N39), .S(n43), .Z(n232) );
  MUX2_X1 U52 ( .A(n33), .B(N39), .S(n243), .Z(n201) );
  MUX2_X1 U53 ( .A(n34), .B(N38), .S(n43), .Z(n233) );
  MUX2_X1 U54 ( .A(n34), .B(N38), .S(n243), .Z(n215) );
  MUX2_X1 U55 ( .A(n35), .B(N37), .S(n43), .Z(n234) );
  MUX2_X1 U56 ( .A(n36), .B(N36), .S(n43), .Z(n235) );
  MUX2_X1 U57 ( .A(n36), .B(N36), .S(n243), .Z(n213) );
  MUX2_X1 U58 ( .A(n37), .B(N35), .S(n43), .Z(n236) );
  MUX2_X1 U59 ( .A(n37), .B(N35), .S(n243), .Z(n212) );
  MUX2_X1 U60 ( .A(n38), .B(N34), .S(n43), .Z(n237) );
  MUX2_X1 U61 ( .A(n38), .B(N34), .S(n243), .Z(n211) );
  MUX2_X1 U62 ( .A(n39), .B(N33), .S(n43), .Z(n238) );
  MUX2_X1 U63 ( .A(n39), .B(N33), .S(n243), .Z(n210) );
  MUX2_X1 U64 ( .A(n40), .B(N32), .S(n43), .Z(n239) );
  MUX2_X1 U65 ( .A(n40), .B(N32), .S(n243), .Z(n209) );
  MUX2_X1 U66 ( .A(n41), .B(N31), .S(n43), .Z(n240) );
  MUX2_X1 U67 ( .A(n41), .B(N31), .S(n243), .Z(n208) );
  MUX2_X1 U68 ( .A(n42), .B(N30), .S(n43), .Z(n241) );
  MUX2_X1 U69 ( .A(n42), .B(N30), .S(n243), .Z(n207) );
  MUX2_X1 U70 ( .A(n44), .B(N29), .S(n43), .Z(n242) );
  MUX2_X1 U71 ( .A(n44), .B(N29), .S(n243), .Z(n200) );
  INV_X1 U72 ( .A(n45), .ZN(n46) );
  OAI21_X1 U73 ( .B1(n46), .B2(n1), .A(n22), .ZN(n47) );
  AOI222_X1 U74 ( .A1(data_out_b[11]), .A2(n21), .B1(adder[11]), .B2(n19), 
        .C1(n67), .C2(n51), .ZN(n52) );
  INV_X1 U75 ( .A(n52), .ZN(n80) );
  AOI222_X1 U76 ( .A1(data_out_b[10]), .A2(n21), .B1(adder[10]), .B2(n19), 
        .C1(n67), .C2(n53), .ZN(n54) );
  INV_X1 U77 ( .A(n54), .ZN(n81) );
  AOI222_X1 U78 ( .A1(data_out_b[8]), .A2(n21), .B1(adder[8]), .B2(n19), .C1(
        n67), .C2(f[8]), .ZN(n55) );
  INV_X1 U79 ( .A(n55), .ZN(n83) );
  AOI222_X1 U80 ( .A1(data_out_b[7]), .A2(n21), .B1(adder[7]), .B2(n19), .C1(
        n67), .C2(f[7]), .ZN(n56) );
  INV_X1 U81 ( .A(n56), .ZN(n84) );
  AOI222_X1 U82 ( .A1(data_out_b[6]), .A2(n21), .B1(adder[6]), .B2(n19), .C1(
        n67), .C2(f[6]), .ZN(n57) );
  INV_X1 U83 ( .A(n57), .ZN(n85) );
  AOI222_X1 U84 ( .A1(data_out_b[5]), .A2(n21), .B1(adder[5]), .B2(n19), .C1(
        n67), .C2(f[5]), .ZN(n58) );
  INV_X1 U85 ( .A(n58), .ZN(n87) );
  AOI222_X1 U86 ( .A1(data_out_b[4]), .A2(n21), .B1(adder[4]), .B2(n19), .C1(
        n67), .C2(f[4]), .ZN(n59) );
  INV_X1 U87 ( .A(n59), .ZN(n104) );
  AOI222_X1 U88 ( .A1(data_out_b[3]), .A2(n21), .B1(adder[3]), .B2(n19), .C1(
        n67), .C2(f[3]), .ZN(n60) );
  INV_X1 U89 ( .A(n60), .ZN(n113) );
  AOI222_X1 U90 ( .A1(data_out_b[2]), .A2(n21), .B1(adder[2]), .B2(n19), .C1(
        n67), .C2(n61), .ZN(n62) );
  INV_X1 U91 ( .A(n62), .ZN(n114) );
  AOI222_X1 U92 ( .A1(data_out_b[1]), .A2(n21), .B1(adder[1]), .B2(n19), .C1(
        n67), .C2(n63), .ZN(n64) );
  INV_X1 U93 ( .A(n64), .ZN(n115) );
  AOI222_X1 U94 ( .A1(data_out_b[0]), .A2(n21), .B1(adder[0]), .B2(n19), .C1(
        n67), .C2(n65), .ZN(n66) );
  INV_X1 U95 ( .A(n66), .ZN(n116) );
  AOI222_X1 U96 ( .A1(data_out_b[9]), .A2(n21), .B1(adder[9]), .B2(n19), .C1(
        n67), .C2(f[9]), .ZN(n68) );
  INV_X1 U97 ( .A(n68), .ZN(n82) );
  NOR4_X1 U98 ( .A1(n51), .A2(n50), .A3(n49), .A4(n48), .ZN(n76) );
  NOR4_X1 U99 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n53), .ZN(n75) );
  NAND4_X1 U100 ( .A1(n72), .A2(n71), .A3(n70), .A4(n69), .ZN(n73) );
  NOR4_X1 U101 ( .A1(n73), .A2(n65), .A3(n63), .A4(n61), .ZN(n74) );
  NAND3_X1 U102 ( .A1(n76), .A2(n75), .A3(n74), .ZN(n78) );
  NAND3_X1 U103 ( .A1(wr_en_y), .A2(n78), .A3(n77), .ZN(n244) );
  OAI22_X1 U104 ( .A1(n184), .A2(n245), .B1(n216), .B2(n244), .ZN(n183) );
  OAI22_X1 U105 ( .A1(n185), .A2(n245), .B1(n217), .B2(n244), .ZN(n182) );
  OAI22_X1 U106 ( .A1(n186), .A2(n245), .B1(n218), .B2(n244), .ZN(n181) );
  OAI22_X1 U107 ( .A1(n194), .A2(n245), .B1(n222), .B2(n244), .ZN(n173) );
  OAI22_X1 U108 ( .A1(n195), .A2(n245), .B1(n223), .B2(n244), .ZN(n172) );
  OAI22_X1 U109 ( .A1(n196), .A2(n245), .B1(n224), .B2(n244), .ZN(n171) );
  OAI22_X1 U110 ( .A1(n197), .A2(n245), .B1(n225), .B2(n244), .ZN(n170) );
  OAI22_X1 U111 ( .A1(n198), .A2(n245), .B1(n226), .B2(n244), .ZN(n169) );
  OAI22_X1 U112 ( .A1(n199), .A2(n245), .B1(n77), .B2(n244), .ZN(n168) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_10_DW_mult_tc_1 ( a, b, 
        product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n9, n12, n13, n16, n18, n19, n21, n23, n25, n27, n29, n31,
         n32, n34, n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n50,
         n52, n53, n54, n55, n56, n57, n58, n59, n62, n63, n64, n65, n67, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n93, n95, n97, n98, n99, n103,
         n104, n105, n106, n107, n109, n111, n112, n113, n114, n115, n117,
         n119, n120, n122, n127, n131, n133, n135, n139, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n237, n245, n247, n249, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n418, n419, n420, n421, n422, n423, n424, n426, n427, n429,
         n433, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U148 ( .A(n265), .B(n144), .Z(n145) );
  XOR2_X1 U150 ( .A(n271), .B(n146), .Z(n147) );
  XOR2_X1 U152 ( .A(n301), .B(n148), .Z(n149) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U161 ( .A(n177), .B(n168), .CI(n166), .CO(n163), .S(n164) );
  FA_X1 U162 ( .A(n170), .B(n172), .CI(n179), .CO(n165), .S(n166) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n263), .CI(n291), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n317), .B(n252), .CO(n173), .S(n174) );
  FA_X1 U167 ( .A(n180), .B(n187), .CI(n178), .CO(n175), .S(n176) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U169 ( .A(n193), .B(n282), .CI(n191), .CO(n179), .S(n180) );
  FA_X1 U170 ( .A(n268), .B(n274), .CI(n292), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U172 ( .A(n197), .B(n190), .CI(n188), .CO(n185), .S(n186) );
  FA_X1 U173 ( .A(n199), .B(n201), .CI(n192), .CO(n187), .S(n188) );
  FA_X1 U174 ( .A(n275), .B(n293), .CI(n194), .CO(n189), .S(n190) );
  FA_X1 U175 ( .A(n305), .B(n253), .CI(n283), .CO(n191), .S(n192) );
  HA_X1 U176 ( .A(n269), .B(n319), .CO(n193), .S(n194) );
  FA_X1 U177 ( .A(n205), .B(n200), .CI(n198), .CO(n195), .S(n196) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U179 ( .A(n284), .B(n276), .CI(n294), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n320), .B(n270), .CI(n306), .CO(n201), .S(n202) );
  FA_X1 U182 ( .A(n215), .B(n307), .CI(n210), .CO(n205), .S(n206) );
  FA_X1 U183 ( .A(n254), .B(n285), .CI(n295), .CO(n207), .S(n208) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U185 ( .A(n216), .B(n219), .CI(n214), .CO(n211), .S(n212) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n322), .B(n278), .CI(n308), .CO(n215), .S(n216) );
  HA_X1 U190 ( .A(n287), .B(n323), .CO(n221), .S(n222) );
  FA_X1 U191 ( .A(n229), .B(n298), .CI(n226), .CO(n223), .S(n224) );
  FA_X1 U192 ( .A(n324), .B(n288), .CI(n310), .CO(n225), .S(n226) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  HA_X1 U194 ( .A(n311), .B(n325), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n326), .B(n312), .CI(n300), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  INV_X1 U414 ( .A(n491), .ZN(n490) );
  CLKBUF_X2 U415 ( .A(n7), .Z(n491) );
  XOR2_X1 U416 ( .A(n13), .B(a[6]), .Z(n553) );
  BUF_X4 U417 ( .A(n9), .Z(n566) );
  CLKBUF_X3 U418 ( .A(n19), .Z(n544) );
  NOR2_X1 U419 ( .A1(n218), .A2(n223), .ZN(n97) );
  OR2_X1 U420 ( .A1(n164), .A2(n175), .ZN(n492) );
  OR2_X1 U421 ( .A1(n329), .A2(n258), .ZN(n493) );
  OR2_X1 U422 ( .A1(n224), .A2(n227), .ZN(n494) );
  OR2_X1 U423 ( .A1(n224), .A2(n227), .ZN(n559) );
  XNOR2_X1 U424 ( .A(n45), .B(n495), .ZN(product[12]) );
  AND2_X1 U425 ( .A1(n531), .A2(n79), .ZN(n495) );
  AND2_X1 U426 ( .A1(n224), .A2(n227), .ZN(n496) );
  BUF_X1 U427 ( .A(n16), .Z(n536) );
  BUF_X2 U428 ( .A(n16), .Z(n565) );
  INV_X1 U429 ( .A(n1), .ZN(n497) );
  INV_X1 U430 ( .A(n1), .ZN(n572) );
  OR2_X1 U431 ( .A1(n196), .A2(n203), .ZN(n498) );
  INV_X1 U432 ( .A(n537), .ZN(n499) );
  NOR2_X1 U433 ( .A1(n164), .A2(n175), .ZN(n500) );
  NOR2_X1 U434 ( .A1(n164), .A2(n175), .ZN(n75) );
  XNOR2_X1 U435 ( .A(n577), .B(a[4]), .ZN(n554) );
  INV_X1 U436 ( .A(n580), .ZN(n501) );
  INV_X1 U437 ( .A(n580), .ZN(n579) );
  INV_X1 U438 ( .A(n545), .ZN(n502) );
  INV_X1 U439 ( .A(n539), .ZN(n503) );
  INV_X1 U440 ( .A(n553), .ZN(n504) );
  NAND2_X1 U441 ( .A1(n525), .A2(n526), .ZN(n505) );
  NAND2_X1 U442 ( .A1(n525), .A2(n526), .ZN(n506) );
  NAND2_X1 U443 ( .A1(n525), .A2(n526), .ZN(n12) );
  OR2_X2 U444 ( .A1(n527), .A2(n553), .ZN(n507) );
  OR2_X1 U445 ( .A1(n527), .A2(n553), .ZN(n23) );
  NAND2_X1 U446 ( .A1(n554), .A2(n536), .ZN(n508) );
  NAND2_X1 U447 ( .A1(n554), .A2(n536), .ZN(n509) );
  NAND2_X1 U448 ( .A1(n554), .A2(n536), .ZN(n18) );
  CLKBUF_X1 U449 ( .A(n74), .Z(n510) );
  XOR2_X1 U450 ( .A(n255), .B(n309), .Z(n511) );
  XOR2_X1 U451 ( .A(n511), .B(n297), .Z(n220) );
  XOR2_X1 U452 ( .A(n225), .B(n222), .Z(n512) );
  XOR2_X1 U453 ( .A(n512), .B(n220), .Z(n218) );
  NAND2_X1 U454 ( .A1(n255), .A2(n309), .ZN(n513) );
  NAND2_X1 U455 ( .A1(n255), .A2(n297), .ZN(n514) );
  NAND2_X1 U456 ( .A1(n309), .A2(n297), .ZN(n515) );
  NAND3_X1 U457 ( .A1(n513), .A2(n514), .A3(n515), .ZN(n219) );
  NAND2_X1 U458 ( .A1(n225), .A2(n222), .ZN(n516) );
  NAND2_X1 U459 ( .A1(n225), .A2(n220), .ZN(n517) );
  NAND2_X1 U460 ( .A1(n222), .A2(n220), .ZN(n518) );
  NAND3_X1 U461 ( .A1(n516), .A2(n517), .A3(n518), .ZN(n217) );
  OR2_X2 U462 ( .A1(n519), .A2(n546), .ZN(n34) );
  XNOR2_X1 U463 ( .A(n581), .B(a[10]), .ZN(n519) );
  XOR2_X1 U464 ( .A(n208), .B(n213), .Z(n520) );
  XOR2_X1 U465 ( .A(n206), .B(n520), .Z(n204) );
  NAND2_X1 U466 ( .A1(n206), .A2(n208), .ZN(n521) );
  NAND2_X1 U467 ( .A1(n206), .A2(n213), .ZN(n522) );
  NAND2_X1 U468 ( .A1(n208), .A2(n213), .ZN(n523) );
  NAND3_X1 U469 ( .A1(n521), .A2(n522), .A3(n523), .ZN(n203) );
  NOR2_X2 U470 ( .A1(n228), .A2(n231), .ZN(n105) );
  CLKBUF_X1 U471 ( .A(n85), .Z(n524) );
  XNOR2_X1 U472 ( .A(n574), .B(a[2]), .ZN(n525) );
  XOR2_X1 U473 ( .A(n572), .B(a[2]), .Z(n526) );
  XNOR2_X1 U474 ( .A(n544), .B(a[6]), .ZN(n527) );
  BUF_X1 U475 ( .A(n573), .Z(n528) );
  BUF_X1 U476 ( .A(n573), .Z(n529) );
  BUF_X1 U477 ( .A(n573), .Z(n530) );
  OR2_X1 U478 ( .A1(n176), .A2(n185), .ZN(n531) );
  OR2_X1 U479 ( .A1(n204), .A2(n211), .ZN(n532) );
  AOI21_X1 U480 ( .B1(n104), .B2(n494), .A(n496), .ZN(n533) );
  AOI21_X1 U481 ( .B1(n104), .B2(n559), .A(n496), .ZN(n99) );
  INV_X1 U482 ( .A(n570), .ZN(n534) );
  INV_X2 U483 ( .A(n497), .ZN(n570) );
  BUF_X2 U484 ( .A(n569), .Z(n535) );
  INV_X1 U485 ( .A(n249), .ZN(n569) );
  INV_X1 U486 ( .A(n577), .ZN(n537) );
  AOI21_X2 U487 ( .B1(n557), .B2(n112), .A(n109), .ZN(n107) );
  INV_X1 U488 ( .A(n553), .ZN(n21) );
  OAI21_X1 U489 ( .B1(n105), .B2(n107), .A(n106), .ZN(n538) );
  INV_X1 U490 ( .A(n545), .ZN(n27) );
  INV_X1 U491 ( .A(n546), .ZN(n32) );
  INV_X1 U492 ( .A(n582), .ZN(n539) );
  INV_X1 U493 ( .A(n582), .ZN(n540) );
  OAI21_X1 U494 ( .B1(n99), .B2(n97), .A(n98), .ZN(n541) );
  OAI21_X1 U495 ( .B1(n533), .B2(n97), .A(n98), .ZN(n542) );
  NAND2_X1 U496 ( .A1(n433), .A2(n569), .ZN(n543) );
  INV_X1 U497 ( .A(n572), .ZN(n571) );
  XOR2_X1 U498 ( .A(n574), .B(a[4]), .Z(n16) );
  XNOR2_X1 U499 ( .A(n578), .B(a[8]), .ZN(n545) );
  XNOR2_X1 U500 ( .A(n580), .B(a[10]), .ZN(n546) );
  XNOR2_X1 U501 ( .A(n88), .B(n547), .ZN(product[10]) );
  NAND2_X1 U502 ( .A1(n498), .A2(n86), .ZN(n547) );
  NAND2_X2 U503 ( .A1(n429), .A2(n27), .ZN(n29) );
  XOR2_X1 U504 ( .A(n572), .B(a[2]), .Z(n9) );
  XNOR2_X1 U505 ( .A(n497), .B(n249), .ZN(n433) );
  OAI21_X1 U506 ( .B1(n89), .B2(n549), .A(n90), .ZN(n548) );
  AOI21_X1 U507 ( .B1(n541), .B2(n556), .A(n93), .ZN(n549) );
  OAI21_X1 U508 ( .B1(n91), .B2(n89), .A(n90), .ZN(n88) );
  NOR2_X2 U509 ( .A1(n186), .A2(n195), .ZN(n82) );
  NAND2_X1 U510 ( .A1(n433), .A2(n569), .ZN(n550) );
  NAND2_X1 U511 ( .A1(n433), .A2(n569), .ZN(n551) );
  AOI21_X1 U512 ( .B1(n548), .B2(n80), .A(n81), .ZN(n552) );
  BUF_X1 U513 ( .A(n43), .Z(n567) );
  NAND2_X1 U514 ( .A1(n555), .A2(n69), .ZN(n47) );
  INV_X1 U515 ( .A(n73), .ZN(n71) );
  AOI21_X1 U516 ( .B1(n510), .B2(n555), .A(n67), .ZN(n65) );
  INV_X1 U517 ( .A(n69), .ZN(n67) );
  INV_X1 U518 ( .A(n74), .ZN(n72) );
  NAND2_X1 U519 ( .A1(n73), .A2(n555), .ZN(n64) );
  INV_X1 U520 ( .A(n95), .ZN(n93) );
  XNOR2_X1 U521 ( .A(n84), .B(n50), .ZN(product[11]) );
  NAND2_X1 U522 ( .A1(n127), .A2(n83), .ZN(n50) );
  INV_X1 U523 ( .A(n82), .ZN(n127) );
  NAND2_X1 U524 ( .A1(n532), .A2(n90), .ZN(n52) );
  OR2_X1 U525 ( .A1(n152), .A2(n163), .ZN(n555) );
  OAI21_X1 U526 ( .B1(n500), .B2(n79), .A(n76), .ZN(n74) );
  NAND2_X1 U527 ( .A1(n492), .A2(n76), .ZN(n48) );
  NOR2_X1 U528 ( .A1(n75), .A2(n78), .ZN(n73) );
  NAND2_X1 U529 ( .A1(n152), .A2(n163), .ZN(n69) );
  NOR2_X1 U530 ( .A1(n82), .A2(n85), .ZN(n80) );
  NAND2_X1 U531 ( .A1(n556), .A2(n95), .ZN(n53) );
  INV_X1 U532 ( .A(n119), .ZN(n117) );
  NAND2_X1 U533 ( .A1(n133), .A2(n106), .ZN(n56) );
  INV_X1 U534 ( .A(n105), .ZN(n133) );
  NAND2_X1 U535 ( .A1(n131), .A2(n98), .ZN(n54) );
  INV_X1 U536 ( .A(n97), .ZN(n131) );
  INV_X1 U537 ( .A(n111), .ZN(n109) );
  NOR2_X1 U538 ( .A1(n176), .A2(n185), .ZN(n78) );
  NOR2_X1 U539 ( .A1(n196), .A2(n203), .ZN(n85) );
  NAND2_X1 U540 ( .A1(n557), .A2(n111), .ZN(n57) );
  NAND2_X1 U541 ( .A1(n494), .A2(n103), .ZN(n55) );
  NAND2_X1 U542 ( .A1(n558), .A2(n119), .ZN(n59) );
  OAI21_X1 U543 ( .B1(n113), .B2(n115), .A(n114), .ZN(n112) );
  NAND2_X1 U544 ( .A1(n176), .A2(n185), .ZN(n79) );
  NAND2_X1 U545 ( .A1(n164), .A2(n175), .ZN(n76) );
  NAND2_X1 U546 ( .A1(n212), .A2(n217), .ZN(n95) );
  NAND2_X1 U547 ( .A1(n186), .A2(n195), .ZN(n83) );
  OR2_X1 U548 ( .A1(n212), .A2(n217), .ZN(n556) );
  NAND2_X1 U549 ( .A1(n204), .A2(n211), .ZN(n90) );
  NAND2_X1 U550 ( .A1(n196), .A2(n203), .ZN(n86) );
  XOR2_X1 U551 ( .A(n58), .B(n115), .Z(product[3]) );
  NAND2_X1 U552 ( .A1(n135), .A2(n114), .ZN(n58) );
  INV_X1 U553 ( .A(n113), .ZN(n135) );
  NAND2_X1 U554 ( .A1(n328), .A2(n314), .ZN(n119) );
  XNOR2_X1 U555 ( .A(n63), .B(n46), .ZN(product[15]) );
  NAND2_X1 U556 ( .A1(n560), .A2(n62), .ZN(n46) );
  OR2_X1 U557 ( .A1(n232), .A2(n233), .ZN(n557) );
  NAND2_X1 U558 ( .A1(n218), .A2(n223), .ZN(n98) );
  INV_X1 U559 ( .A(n37), .ZN(n237) );
  NAND2_X1 U560 ( .A1(n232), .A2(n233), .ZN(n111) );
  NAND2_X1 U561 ( .A1(n224), .A2(n227), .ZN(n103) );
  OR2_X1 U562 ( .A1(n328), .A2(n314), .ZN(n558) );
  INV_X1 U563 ( .A(n41), .ZN(n235) );
  OR2_X1 U564 ( .A1(n151), .A2(n139), .ZN(n560) );
  AND2_X1 U565 ( .A1(n493), .A2(n122), .ZN(product[1]) );
  XNOR2_X1 U566 ( .A(n581), .B(a[12]), .ZN(n37) );
  XNOR2_X1 U567 ( .A(n583), .B(a[14]), .ZN(n41) );
  NAND2_X1 U568 ( .A1(n433), .A2(n569), .ZN(n6) );
  OR2_X1 U569 ( .A1(n567), .A2(n490), .ZN(n392) );
  XNOR2_X1 U570 ( .A(n501), .B(n567), .ZN(n352) );
  AND2_X1 U571 ( .A1(n568), .A2(n553), .ZN(n288) );
  AND2_X1 U572 ( .A1(n568), .A2(n245), .ZN(n300) );
  XNOR2_X1 U573 ( .A(n155), .B(n562), .ZN(n139) );
  XNOR2_X1 U574 ( .A(n153), .B(n141), .ZN(n562) );
  XNOR2_X1 U575 ( .A(n157), .B(n563), .ZN(n141) );
  XNOR2_X1 U576 ( .A(n145), .B(n143), .ZN(n563) );
  OAI22_X1 U577 ( .A1(n39), .A2(n336), .B1(n37), .B2(n335), .ZN(n263) );
  OAI22_X1 U578 ( .A1(n39), .A2(n584), .B1(n337), .B2(n37), .ZN(n252) );
  OR2_X1 U579 ( .A1(n567), .A2(n584), .ZN(n337) );
  OAI22_X1 U580 ( .A1(n34), .A2(n343), .B1(n342), .B2(n32), .ZN(n269) );
  XNOR2_X1 U581 ( .A(n540), .B(n567), .ZN(n343) );
  OAI22_X1 U582 ( .A1(n42), .A2(n586), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U583 ( .A1(n567), .A2(n586), .ZN(n332) );
  XOR2_X1 U584 ( .A(n579), .B(a[8]), .Z(n429) );
  XNOR2_X1 U585 ( .A(n159), .B(n564), .ZN(n142) );
  XNOR2_X1 U586 ( .A(n315), .B(n261), .ZN(n564) );
  XNOR2_X1 U587 ( .A(n583), .B(n567), .ZN(n336) );
  AND2_X1 U588 ( .A1(n568), .A2(n247), .ZN(n314) );
  NAND2_X1 U589 ( .A1(n427), .A2(n37), .ZN(n39) );
  XOR2_X1 U590 ( .A(n583), .B(a[12]), .Z(n427) );
  AND2_X1 U591 ( .A1(n568), .A2(n545), .ZN(n278) );
  OAI22_X1 U592 ( .A1(n34), .A2(n342), .B1(n341), .B2(n32), .ZN(n268) );
  OAI22_X1 U593 ( .A1(n34), .A2(n341), .B1(n340), .B2(n32), .ZN(n267) );
  XNOR2_X1 U594 ( .A(n576), .B(n567), .ZN(n376) );
  AND2_X1 U595 ( .A1(n568), .A2(n546), .ZN(n270) );
  AND2_X1 U596 ( .A1(n568), .A2(n235), .ZN(n260) );
  OAI22_X1 U597 ( .A1(n39), .A2(n335), .B1(n37), .B2(n334), .ZN(n262) );
  INV_X1 U598 ( .A(n25), .ZN(n580) );
  OAI22_X1 U599 ( .A1(n34), .A2(n503), .B1(n344), .B2(n32), .ZN(n253) );
  OAI22_X1 U600 ( .A1(n34), .A2(n340), .B1(n339), .B2(n32), .ZN(n266) );
  NAND2_X1 U601 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U602 ( .A(n585), .B(a[14]), .Z(n426) );
  INV_X1 U603 ( .A(n13), .ZN(n577) );
  INV_X1 U604 ( .A(n7), .ZN(n574) );
  XNOR2_X1 U605 ( .A(n544), .B(n567), .ZN(n363) );
  AND2_X1 U606 ( .A1(n568), .A2(n237), .ZN(n264) );
  OR2_X1 U607 ( .A1(n567), .A2(n503), .ZN(n344) );
  AND2_X1 U608 ( .A1(n568), .A2(n249), .ZN(product[0]) );
  OR2_X1 U609 ( .A1(n567), .A2(n580), .ZN(n353) );
  OR2_X1 U610 ( .A1(n567), .A2(n578), .ZN(n364) );
  OR2_X1 U611 ( .A1(n567), .A2(n499), .ZN(n377) );
  XNOR2_X1 U612 ( .A(n544), .B(b[9]), .ZN(n354) );
  OAI22_X1 U613 ( .A1(n39), .A2(n334), .B1(n37), .B2(n333), .ZN(n261) );
  XNOR2_X1 U614 ( .A(n583), .B(n422), .ZN(n333) );
  XNOR2_X1 U615 ( .A(n576), .B(b[11]), .ZN(n365) );
  XNOR2_X1 U616 ( .A(n540), .B(n424), .ZN(n342) );
  XNOR2_X1 U617 ( .A(n539), .B(n423), .ZN(n341) );
  XNOR2_X1 U618 ( .A(n539), .B(n422), .ZN(n340) );
  XNOR2_X1 U619 ( .A(n540), .B(n421), .ZN(n339) );
  XNOR2_X1 U620 ( .A(n583), .B(n423), .ZN(n334) );
  XNOR2_X1 U621 ( .A(n583), .B(n424), .ZN(n335) );
  OAI22_X1 U622 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U623 ( .A(n585), .B(n424), .ZN(n330) );
  XNOR2_X1 U624 ( .A(n585), .B(n567), .ZN(n331) );
  XNOR2_X1 U625 ( .A(n501), .B(n418), .ZN(n345) );
  OAI22_X1 U626 ( .A1(n34), .A2(n339), .B1(n338), .B2(n32), .ZN(n265) );
  XNOR2_X1 U627 ( .A(n539), .B(n420), .ZN(n338) );
  XNOR2_X1 U628 ( .A(n529), .B(b[13]), .ZN(n378) );
  XNOR2_X1 U629 ( .A(n544), .B(n424), .ZN(n362) );
  XNOR2_X1 U630 ( .A(n579), .B(n424), .ZN(n351) );
  XNOR2_X1 U631 ( .A(n528), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U632 ( .A(n528), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U633 ( .A(n529), .B(n418), .ZN(n384) );
  XNOR2_X1 U634 ( .A(n530), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U635 ( .A(n530), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U636 ( .A(n530), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U637 ( .A(n529), .B(n419), .ZN(n385) );
  XNOR2_X1 U638 ( .A(n576), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U639 ( .A(n576), .B(n418), .ZN(n369) );
  XNOR2_X1 U640 ( .A(n576), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U641 ( .A(n576), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U642 ( .A(n579), .B(n423), .ZN(n350) );
  XNOR2_X1 U643 ( .A(n501), .B(n422), .ZN(n349) );
  XNOR2_X1 U644 ( .A(n544), .B(n423), .ZN(n361) );
  XNOR2_X1 U645 ( .A(n544), .B(n422), .ZN(n360) );
  XNOR2_X1 U646 ( .A(n570), .B(b[11]), .ZN(n397) );
  XNOR2_X1 U647 ( .A(n570), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U648 ( .A(n570), .B(b[13]), .ZN(n395) );
  XNOR2_X1 U649 ( .A(n570), .B(b[14]), .ZN(n394) );
  XNOR2_X1 U650 ( .A(n544), .B(n421), .ZN(n359) );
  XNOR2_X1 U651 ( .A(n544), .B(n420), .ZN(n358) );
  XNOR2_X1 U652 ( .A(n501), .B(n421), .ZN(n348) );
  XNOR2_X1 U653 ( .A(n579), .B(n420), .ZN(n347) );
  XNOR2_X1 U654 ( .A(n544), .B(n418), .ZN(n356) );
  XNOR2_X1 U655 ( .A(n501), .B(n419), .ZN(n346) );
  XNOR2_X1 U656 ( .A(n544), .B(n419), .ZN(n357) );
  XNOR2_X1 U657 ( .A(n544), .B(b[8]), .ZN(n355) );
  XNOR2_X1 U658 ( .A(n570), .B(b[15]), .ZN(n393) );
  BUF_X1 U659 ( .A(n43), .Z(n568) );
  OAI22_X1 U660 ( .A1(n551), .A2(n395), .B1(n394), .B2(n535), .ZN(n316) );
  OAI22_X1 U661 ( .A1(n543), .A2(n394), .B1(n393), .B2(n535), .ZN(n315) );
  OAI22_X1 U662 ( .A1(n550), .A2(n404), .B1(n403), .B2(n569), .ZN(n325) );
  OAI22_X1 U663 ( .A1(n551), .A2(n401), .B1(n400), .B2(n535), .ZN(n322) );
  OAI22_X1 U664 ( .A1(n543), .A2(n400), .B1(n399), .B2(n535), .ZN(n321) );
  OAI22_X1 U665 ( .A1(n551), .A2(n406), .B1(n405), .B2(n535), .ZN(n327) );
  OAI22_X1 U666 ( .A1(n550), .A2(n396), .B1(n395), .B2(n535), .ZN(n317) );
  OAI22_X1 U667 ( .A1(n6), .A2(n397), .B1(n396), .B2(n535), .ZN(n318) );
  OAI22_X1 U668 ( .A1(n551), .A2(n399), .B1(n398), .B2(n569), .ZN(n320) );
  OAI22_X1 U669 ( .A1(n550), .A2(n398), .B1(n397), .B2(n535), .ZN(n319) );
  OAI22_X1 U670 ( .A1(n543), .A2(n408), .B1(n407), .B2(n535), .ZN(n329) );
  OAI22_X1 U671 ( .A1(n551), .A2(n405), .B1(n404), .B2(n569), .ZN(n326) );
  OAI22_X1 U672 ( .A1(n6), .A2(n402), .B1(n401), .B2(n535), .ZN(n323) );
  OAI22_X1 U673 ( .A1(n6), .A2(n403), .B1(n402), .B2(n569), .ZN(n324) );
  OAI22_X1 U674 ( .A1(n550), .A2(n407), .B1(n406), .B2(n535), .ZN(n328) );
  NAND2_X1 U675 ( .A1(n228), .A2(n231), .ZN(n106) );
  INV_X1 U676 ( .A(n19), .ZN(n578) );
  OAI21_X1 U677 ( .B1(n87), .B2(n524), .A(n86), .ZN(n84) );
  NOR2_X1 U678 ( .A1(n204), .A2(n211), .ZN(n89) );
  OAI22_X1 U679 ( .A1(n29), .A2(n350), .B1(n349), .B2(n502), .ZN(n275) );
  OAI22_X1 U680 ( .A1(n29), .A2(n346), .B1(n345), .B2(n502), .ZN(n271) );
  OAI22_X1 U681 ( .A1(n29), .A2(n347), .B1(n346), .B2(n502), .ZN(n272) );
  OAI22_X1 U682 ( .A1(n29), .A2(n349), .B1(n348), .B2(n502), .ZN(n274) );
  OAI22_X1 U683 ( .A1(n29), .A2(n351), .B1(n350), .B2(n502), .ZN(n276) );
  OAI22_X1 U684 ( .A1(n29), .A2(n348), .B1(n347), .B2(n502), .ZN(n273) );
  OAI22_X1 U685 ( .A1(n29), .A2(n580), .B1(n353), .B2(n502), .ZN(n254) );
  OAI22_X1 U686 ( .A1(n29), .A2(n352), .B1(n351), .B2(n502), .ZN(n277) );
  INV_X1 U687 ( .A(n88), .ZN(n87) );
  XNOR2_X1 U688 ( .A(n59), .B(n120), .ZN(product[2]) );
  AOI21_X1 U689 ( .B1(n558), .B2(n120), .A(n117), .ZN(n115) );
  XNOR2_X1 U690 ( .A(n537), .B(n424), .ZN(n375) );
  XNOR2_X1 U691 ( .A(n575), .B(n419), .ZN(n370) );
  XNOR2_X1 U692 ( .A(n575), .B(n420), .ZN(n371) );
  XNOR2_X1 U693 ( .A(n537), .B(n423), .ZN(n374) );
  XNOR2_X1 U694 ( .A(n537), .B(n422), .ZN(n373) );
  XNOR2_X1 U695 ( .A(n575), .B(n421), .ZN(n372) );
  XNOR2_X1 U696 ( .A(n77), .B(n48), .ZN(product[13]) );
  OAI21_X1 U697 ( .B1(n105), .B2(n107), .A(n106), .ZN(n104) );
  XOR2_X1 U698 ( .A(n56), .B(n107), .Z(product[5]) );
  NOR2_X1 U699 ( .A1(n234), .A2(n257), .ZN(n113) );
  XNOR2_X1 U700 ( .A(n57), .B(n112), .ZN(product[4]) );
  AOI21_X1 U701 ( .B1(n541), .B2(n556), .A(n93), .ZN(n91) );
  OAI22_X1 U702 ( .A1(n507), .A2(n356), .B1(n355), .B2(n504), .ZN(n280) );
  OAI22_X1 U703 ( .A1(n507), .A2(n358), .B1(n357), .B2(n504), .ZN(n282) );
  OAI22_X1 U704 ( .A1(n507), .A2(n355), .B1(n354), .B2(n504), .ZN(n279) );
  OAI22_X1 U705 ( .A1(n507), .A2(n360), .B1(n359), .B2(n21), .ZN(n284) );
  OAI22_X1 U706 ( .A1(n507), .A2(n362), .B1(n361), .B2(n504), .ZN(n286) );
  OAI22_X1 U707 ( .A1(n507), .A2(n361), .B1(n360), .B2(n504), .ZN(n285) );
  OAI22_X1 U708 ( .A1(n23), .A2(n578), .B1(n364), .B2(n21), .ZN(n255) );
  OAI22_X1 U709 ( .A1(n507), .A2(n357), .B1(n356), .B2(n504), .ZN(n281) );
  OAI22_X1 U710 ( .A1(n23), .A2(n363), .B1(n362), .B2(n21), .ZN(n287) );
  OAI22_X1 U711 ( .A1(n23), .A2(n359), .B1(n358), .B2(n21), .ZN(n283) );
  OR2_X1 U712 ( .A1(n567), .A2(n534), .ZN(n409) );
  OAI21_X1 U713 ( .B1(n82), .B2(n86), .A(n83), .ZN(n81) );
  XNOR2_X1 U714 ( .A(n55), .B(n538), .ZN(product[6]) );
  NAND2_X1 U715 ( .A1(n151), .A2(n139), .ZN(n62) );
  OAI22_X1 U716 ( .A1(n509), .A2(n370), .B1(n369), .B2(n565), .ZN(n293) );
  OAI22_X1 U717 ( .A1(n508), .A2(n367), .B1(n366), .B2(n565), .ZN(n290) );
  OAI22_X1 U718 ( .A1(n508), .A2(n375), .B1(n374), .B2(n565), .ZN(n298) );
  OAI22_X1 U719 ( .A1(n18), .A2(n368), .B1(n367), .B2(n565), .ZN(n291) );
  OAI22_X1 U720 ( .A1(n509), .A2(n372), .B1(n371), .B2(n565), .ZN(n295) );
  OAI22_X1 U721 ( .A1(n508), .A2(n373), .B1(n372), .B2(n565), .ZN(n296) );
  OAI22_X1 U722 ( .A1(n508), .A2(n376), .B1(n375), .B2(n565), .ZN(n299) );
  OAI22_X1 U723 ( .A1(n509), .A2(n499), .B1(n377), .B2(n565), .ZN(n256) );
  OAI22_X1 U724 ( .A1(n509), .A2(n369), .B1(n368), .B2(n565), .ZN(n292) );
  OAI22_X1 U725 ( .A1(n508), .A2(n371), .B1(n370), .B2(n565), .ZN(n294) );
  OAI22_X1 U726 ( .A1(n509), .A2(n374), .B1(n373), .B2(n565), .ZN(n297) );
  OAI22_X1 U727 ( .A1(n18), .A2(n366), .B1(n365), .B2(n565), .ZN(n289) );
  XNOR2_X1 U728 ( .A(n491), .B(n420), .ZN(n386) );
  INV_X1 U729 ( .A(n536), .ZN(n245) );
  XNOR2_X1 U730 ( .A(n491), .B(n422), .ZN(n388) );
  XNOR2_X1 U731 ( .A(n491), .B(n421), .ZN(n387) );
  XNOR2_X1 U732 ( .A(n491), .B(n567), .ZN(n391) );
  XNOR2_X1 U733 ( .A(n491), .B(n423), .ZN(n389) );
  XNOR2_X1 U734 ( .A(n491), .B(n424), .ZN(n390) );
  XNOR2_X1 U735 ( .A(n570), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U736 ( .A(n571), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U737 ( .A(n571), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U738 ( .A(n570), .B(n418), .ZN(n401) );
  XNOR2_X1 U739 ( .A(n571), .B(n419), .ZN(n402) );
  XNOR2_X1 U740 ( .A(n571), .B(n420), .ZN(n403) );
  XNOR2_X1 U741 ( .A(n571), .B(n422), .ZN(n405) );
  XNOR2_X1 U742 ( .A(n571), .B(n421), .ZN(n404) );
  XNOR2_X1 U743 ( .A(n570), .B(n567), .ZN(n408) );
  XNOR2_X1 U744 ( .A(n570), .B(n423), .ZN(n406) );
  XNOR2_X1 U745 ( .A(n570), .B(n424), .ZN(n407) );
  XOR2_X1 U746 ( .A(n549), .B(n52), .Z(product[9]) );
  OAI21_X1 U747 ( .B1(n552), .B2(n71), .A(n72), .ZN(n70) );
  OAI21_X1 U748 ( .B1(n45), .B2(n78), .A(n79), .ZN(n77) );
  XNOR2_X1 U749 ( .A(n70), .B(n47), .ZN(product[14]) );
  OAI21_X1 U750 ( .B1(n64), .B2(n552), .A(n65), .ZN(n63) );
  AOI21_X1 U751 ( .B1(n80), .B2(n548), .A(n81), .ZN(n45) );
  XNOR2_X1 U752 ( .A(n53), .B(n542), .ZN(product[8]) );
  INV_X1 U753 ( .A(n122), .ZN(n120) );
  NAND2_X1 U754 ( .A1(n329), .A2(n258), .ZN(n122) );
  OAI22_X1 U755 ( .A1(n550), .A2(n534), .B1(n409), .B2(n569), .ZN(n258) );
  XOR2_X1 U756 ( .A(n533), .B(n54), .Z(product[7]) );
  OAI22_X1 U757 ( .A1(n506), .A2(n379), .B1(n378), .B2(n566), .ZN(n301) );
  OAI22_X1 U758 ( .A1(n505), .A2(n380), .B1(n379), .B2(n566), .ZN(n302) );
  OAI22_X1 U759 ( .A1(n505), .A2(n385), .B1(n384), .B2(n566), .ZN(n307) );
  OAI22_X1 U760 ( .A1(n506), .A2(n382), .B1(n381), .B2(n566), .ZN(n304) );
  OAI22_X1 U761 ( .A1(n505), .A2(n381), .B1(n380), .B2(n566), .ZN(n303) );
  NAND2_X1 U762 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U763 ( .A1(n505), .A2(n383), .B1(n382), .B2(n566), .ZN(n305) );
  OAI22_X1 U764 ( .A1(n505), .A2(n384), .B1(n383), .B2(n566), .ZN(n306) );
  OAI22_X1 U765 ( .A1(n505), .A2(n386), .B1(n385), .B2(n566), .ZN(n308) );
  OAI22_X1 U766 ( .A1(n506), .A2(n387), .B1(n386), .B2(n566), .ZN(n309) );
  OAI22_X1 U767 ( .A1(n506), .A2(n490), .B1(n392), .B2(n566), .ZN(n257) );
  OAI22_X1 U768 ( .A1(n12), .A2(n389), .B1(n388), .B2(n566), .ZN(n311) );
  OAI22_X1 U769 ( .A1(n12), .A2(n388), .B1(n387), .B2(n566), .ZN(n310) );
  OAI22_X1 U770 ( .A1(n12), .A2(n390), .B1(n389), .B2(n566), .ZN(n312) );
  INV_X1 U771 ( .A(n566), .ZN(n247) );
  OAI22_X1 U772 ( .A1(n506), .A2(n391), .B1(n390), .B2(n566), .ZN(n313) );
  INV_X1 U773 ( .A(n574), .ZN(n573) );
  INV_X1 U774 ( .A(n577), .ZN(n575) );
  INV_X1 U775 ( .A(n577), .ZN(n576) );
  INV_X1 U776 ( .A(n582), .ZN(n581) );
  INV_X1 U777 ( .A(n31), .ZN(n582) );
  INV_X1 U778 ( .A(n584), .ZN(n583) );
  INV_X1 U779 ( .A(n36), .ZN(n584) );
  INV_X1 U780 ( .A(n586), .ZN(n585) );
  INV_X1 U781 ( .A(n40), .ZN(n586) );
  XOR2_X1 U782 ( .A(n259), .B(n251), .Z(n148) );
  XOR2_X1 U783 ( .A(n289), .B(n279), .Z(n146) );
  XOR2_X1 U784 ( .A(n149), .B(n147), .Z(n144) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_10_DW01_add_2 ( A, B, CI, SUM, 
        CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n7, n8, n9, n10, n11, n12, n13, n14, n15, n18, n19,
         n20, n21, n23, n25, n26, n27, n28, n30, n33, n34, n35, n36, n37, n38,
         n39, n40, n42, n43, n44, n48, n49, n51, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n71, n72, n73, n74,
         n75, n77, n79, n80, n81, n82, n83, n85, n87, n88, n90, n93, n94, n98,
         n99, n100, n102, n104, n161, n162, n163, n164, n165, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185;

  NOR2_X1 U126 ( .A1(A[8]), .A2(B[8]), .ZN(n161) );
  NOR2_X1 U127 ( .A1(A[8]), .A2(B[8]), .ZN(n58) );
  XNOR2_X1 U128 ( .A(n49), .B(n162), .ZN(SUM[10]) );
  AND2_X1 U129 ( .A1(n171), .A2(n48), .ZN(n162) );
  XNOR2_X1 U130 ( .A(n174), .B(n163), .ZN(SUM[11]) );
  NAND2_X1 U131 ( .A1(n165), .A2(n40), .ZN(n163) );
  OAI21_X1 U132 ( .B1(n43), .B2(n55), .A(n44), .ZN(n164) );
  OR2_X1 U133 ( .A1(A[11]), .A2(B[11]), .ZN(n165) );
  NOR2_X1 U134 ( .A1(A[11]), .A2(B[11]), .ZN(n39) );
  AND2_X1 U135 ( .A1(n178), .A2(n90), .ZN(SUM[0]) );
  OR2_X1 U136 ( .A1(A[15]), .A2(B[15]), .ZN(n167) );
  AOI21_X1 U137 ( .B1(n56), .B2(n64), .A(n57), .ZN(n168) );
  AOI21_X1 U138 ( .B1(n56), .B2(n64), .A(n57), .ZN(n169) );
  AOI21_X1 U139 ( .B1(n56), .B2(n64), .A(n57), .ZN(n55) );
  BUF_X1 U140 ( .A(n27), .Z(n170) );
  OR2_X1 U141 ( .A1(A[10]), .A2(B[10]), .ZN(n171) );
  OR2_X1 U142 ( .A1(A[10]), .A2(B[10]), .ZN(n172) );
  OR2_X1 U143 ( .A1(A[10]), .A2(B[10]), .ZN(n182) );
  AOI21_X1 U144 ( .B1(n172), .B2(n51), .A(n176), .ZN(n173) );
  OAI21_X1 U145 ( .B1(n43), .B2(n55), .A(n44), .ZN(n174) );
  NOR2_X1 U146 ( .A1(A[12]), .A2(B[12]), .ZN(n175) );
  NOR2_X1 U147 ( .A1(A[12]), .A2(B[12]), .ZN(n36) );
  AND2_X1 U148 ( .A1(A[10]), .A2(B[10]), .ZN(n176) );
  INV_X1 U149 ( .A(n42), .ZN(n177) );
  OR2_X1 U150 ( .A1(A[0]), .A2(B[0]), .ZN(n178) );
  INV_X1 U151 ( .A(n64), .ZN(n63) );
  INV_X1 U152 ( .A(n168), .ZN(n54) );
  AOI21_X1 U153 ( .B1(n179), .B2(n72), .A(n69), .ZN(n67) );
  INV_X1 U154 ( .A(n71), .ZN(n69) );
  AOI21_X1 U155 ( .B1(n181), .B2(n88), .A(n85), .ZN(n83) );
  INV_X1 U156 ( .A(n87), .ZN(n85) );
  AOI21_X1 U157 ( .B1(n183), .B2(n80), .A(n77), .ZN(n75) );
  INV_X1 U158 ( .A(n79), .ZN(n77) );
  OAI21_X1 U159 ( .B1(n67), .B2(n65), .A(n66), .ZN(n64) );
  OAI21_X1 U160 ( .B1(n83), .B2(n81), .A(n82), .ZN(n80) );
  AOI21_X1 U161 ( .B1(n54), .B2(n180), .A(n51), .ZN(n49) );
  NAND2_X1 U162 ( .A1(n98), .A2(n59), .ZN(n8) );
  INV_X1 U163 ( .A(n90), .ZN(n88) );
  OAI21_X1 U164 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  INV_X1 U165 ( .A(n53), .ZN(n51) );
  NAND2_X1 U166 ( .A1(n100), .A2(n66), .ZN(n10) );
  INV_X1 U167 ( .A(n65), .ZN(n100) );
  NAND2_X1 U168 ( .A1(n179), .A2(n71), .ZN(n11) );
  NAND2_X1 U169 ( .A1(n99), .A2(n62), .ZN(n9) );
  INV_X1 U170 ( .A(n61), .ZN(n99) );
  NAND2_X1 U171 ( .A1(n180), .A2(n53), .ZN(n7) );
  NAND2_X1 U172 ( .A1(n104), .A2(n82), .ZN(n14) );
  INV_X1 U173 ( .A(n81), .ZN(n104) );
  NAND2_X1 U174 ( .A1(n181), .A2(n87), .ZN(n15) );
  NAND2_X1 U175 ( .A1(n183), .A2(n79), .ZN(n13) );
  NAND2_X1 U176 ( .A1(n102), .A2(n74), .ZN(n12) );
  INV_X1 U177 ( .A(n73), .ZN(n102) );
  NAND2_X1 U178 ( .A1(n37), .A2(n94), .ZN(n4) );
  XNOR2_X1 U179 ( .A(n54), .B(n7), .ZN(SUM[9]) );
  XOR2_X1 U180 ( .A(n63), .B(n9), .Z(SUM[7]) );
  XNOR2_X1 U181 ( .A(n15), .B(n88), .ZN(SUM[1]) );
  OR2_X1 U182 ( .A1(A[5]), .A2(B[5]), .ZN(n179) );
  NOR2_X1 U183 ( .A1(A[7]), .A2(B[7]), .ZN(n61) );
  OR2_X1 U184 ( .A1(A[9]), .A2(B[9]), .ZN(n180) );
  NOR2_X1 U185 ( .A1(A[2]), .A2(B[2]), .ZN(n81) );
  NOR2_X1 U186 ( .A1(A[6]), .A2(B[6]), .ZN(n65) );
  NAND2_X1 U187 ( .A1(A[11]), .A2(B[11]), .ZN(n40) );
  OR2_X1 U188 ( .A1(A[1]), .A2(B[1]), .ZN(n181) );
  NAND2_X1 U189 ( .A1(A[3]), .A2(B[3]), .ZN(n79) );
  NOR2_X1 U190 ( .A1(A[13]), .A2(B[13]), .ZN(n27) );
  XNOR2_X1 U191 ( .A(n11), .B(n72), .ZN(SUM[5]) );
  XNOR2_X1 U192 ( .A(n60), .B(n8), .ZN(SUM[8]) );
  NOR2_X1 U193 ( .A1(A[4]), .A2(B[4]), .ZN(n73) );
  NAND2_X1 U194 ( .A1(A[7]), .A2(B[7]), .ZN(n62) );
  OR2_X1 U195 ( .A1(A[3]), .A2(B[3]), .ZN(n183) );
  NAND2_X1 U196 ( .A1(A[2]), .A2(B[2]), .ZN(n82) );
  NAND2_X1 U197 ( .A1(A[6]), .A2(B[6]), .ZN(n66) );
  NAND2_X1 U198 ( .A1(A[9]), .A2(B[9]), .ZN(n53) );
  NAND2_X1 U199 ( .A1(A[1]), .A2(B[1]), .ZN(n87) );
  NAND2_X1 U200 ( .A1(A[0]), .A2(B[0]), .ZN(n90) );
  NAND2_X1 U201 ( .A1(A[8]), .A2(B[8]), .ZN(n59) );
  NAND2_X1 U202 ( .A1(A[4]), .A2(B[4]), .ZN(n74) );
  NAND2_X1 U203 ( .A1(A[12]), .A2(B[12]), .ZN(n37) );
  XOR2_X1 U204 ( .A(n10), .B(n67), .Z(SUM[6]) );
  XNOR2_X1 U205 ( .A(n13), .B(n80), .ZN(SUM[3]) );
  XOR2_X1 U206 ( .A(n14), .B(n83), .Z(SUM[2]) );
  OR2_X1 U207 ( .A1(A[14]), .A2(B[14]), .ZN(n184) );
  NAND2_X1 U208 ( .A1(n167), .A2(n18), .ZN(n1) );
  XOR2_X1 U209 ( .A(n12), .B(n75), .Z(SUM[4]) );
  NAND2_X1 U210 ( .A1(A[5]), .A2(B[5]), .ZN(n71) );
  NAND2_X1 U211 ( .A1(n184), .A2(n25), .ZN(n2) );
  INV_X1 U212 ( .A(n25), .ZN(n23) );
  NAND2_X1 U213 ( .A1(n184), .A2(n93), .ZN(n20) );
  NAND2_X1 U214 ( .A1(n93), .A2(n28), .ZN(n3) );
  XNOR2_X1 U215 ( .A(n38), .B(n4), .ZN(SUM[12]) );
  AOI21_X1 U216 ( .B1(n164), .B2(n34), .A(n35), .ZN(n185) );
  AOI21_X1 U217 ( .B1(n164), .B2(n34), .A(n35), .ZN(n33) );
  NAND2_X1 U218 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  INV_X1 U219 ( .A(n27), .ZN(n93) );
  INV_X1 U220 ( .A(n161), .ZN(n98) );
  NOR2_X1 U221 ( .A1(n161), .A2(n61), .ZN(n56) );
  OAI21_X1 U222 ( .B1(n58), .B2(n62), .A(n59), .ZN(n57) );
  AOI21_X1 U223 ( .B1(n184), .B2(n30), .A(n23), .ZN(n21) );
  INV_X1 U224 ( .A(n28), .ZN(n30) );
  INV_X1 U225 ( .A(n175), .ZN(n94) );
  NOR2_X1 U226 ( .A1(n175), .A2(n39), .ZN(n34) );
  OAI21_X1 U227 ( .B1(n36), .B2(n40), .A(n37), .ZN(n35) );
  OAI21_X1 U228 ( .B1(n75), .B2(n73), .A(n74), .ZN(n72) );
  NAND2_X1 U229 ( .A1(A[14]), .A2(B[14]), .ZN(n25) );
  OAI21_X1 U230 ( .B1(n177), .B2(n39), .A(n40), .ZN(n38) );
  AOI21_X1 U231 ( .B1(n51), .B2(n182), .A(n176), .ZN(n44) );
  NAND2_X1 U232 ( .A1(A[15]), .A2(B[15]), .ZN(n18) );
  OAI21_X1 U233 ( .B1(n43), .B2(n169), .A(n173), .ZN(n42) );
  XNOR2_X1 U234 ( .A(n19), .B(n1), .ZN(SUM[15]) );
  NAND2_X1 U235 ( .A1(n171), .A2(n180), .ZN(n43) );
  XNOR2_X1 U236 ( .A(n26), .B(n2), .ZN(SUM[14]) );
  XOR2_X1 U237 ( .A(n185), .B(n3), .Z(SUM[13]) );
  OAI21_X1 U238 ( .B1(n33), .B2(n170), .A(n28), .ZN(n26) );
  OAI21_X1 U239 ( .B1(n185), .B2(n20), .A(n21), .ZN(n19) );
  NAND2_X1 U240 ( .A1(A[10]), .A2(B[10]), .ZN(n48) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_10 ( clk, clear_acc, 
        data_out_x, data_out, data_out_w, data_out_b, wr_en_y, m_valid, 
        m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [3:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N27, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, n1, n2, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n87, n104, n113, n114, n115, n116, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n22), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n228), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n229), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n230), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n231), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n232), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n233), .CK(clk), .Q(n34) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n234), .CK(clk), .Q(n35) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n235), .CK(clk), .Q(n36) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n236), .CK(clk), .Q(n37) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n237), .CK(clk), .Q(n38) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n238), .CK(clk), .Q(n39) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n239), .CK(clk), .Q(n40) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n240), .CK(clk), .Q(n41) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n241), .CK(clk), .Q(n42) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n242), .CK(clk), .Q(n43) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n243), .CK(clk), .Q(n45) );
  DFF_X1 \f_reg[7]  ( .D(n85), .CK(clk), .Q(f[7]), .QN(n220) );
  DFF_X1 \f_reg[8]  ( .D(n84), .CK(clk), .Q(f[8]), .QN(n221) );
  DFF_X1 \f_reg[9]  ( .D(n83), .CK(clk), .Q(f[9]), .QN(n222) );
  DFF_X1 \f_reg[10]  ( .D(n82), .CK(clk), .Q(n54), .QN(n223) );
  DFF_X1 \f_reg[11]  ( .D(n81), .CK(clk), .Q(n52), .QN(n224) );
  DFF_X1 \f_reg[12]  ( .D(n1), .CK(clk), .Q(n51), .QN(n225) );
  DFF_X1 \f_reg[13]  ( .D(n4), .CK(clk), .Q(n50), .QN(n226) );
  DFF_X1 \f_reg[14]  ( .D(n5), .CK(clk), .Q(n49), .QN(n227) );
  DFF_X1 \f_reg[15]  ( .D(n80), .CK(clk), .Q(f[15]), .QN(n78) );
  DFF_X1 \data_out_reg[15]  ( .D(n169), .CK(clk), .Q(data_out[15]), .QN(n200)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n170), .CK(clk), .Q(data_out[14]), .QN(n199)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n171), .CK(clk), .Q(data_out[13]), .QN(n198)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n172), .CK(clk), .Q(data_out[12]), .QN(n197)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n173), .CK(clk), .Q(data_out[11]), .QN(n196)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n174), .CK(clk), .Q(data_out[10]), .QN(n195)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n175), .CK(clk), .Q(data_out[9]), .QN(n194) );
  DFF_X1 \data_out_reg[8]  ( .D(n176), .CK(clk), .Q(data_out[8]), .QN(n193) );
  DFF_X1 \data_out_reg[7]  ( .D(n177), .CK(clk), .Q(data_out[7]), .QN(n192) );
  DFF_X1 \data_out_reg[6]  ( .D(n178), .CK(clk), .Q(data_out[6]), .QN(n191) );
  DFF_X1 \data_out_reg[5]  ( .D(n179), .CK(clk), .Q(data_out[5]), .QN(n190) );
  DFF_X1 \data_out_reg[4]  ( .D(n180), .CK(clk), .Q(data_out[4]), .QN(n189) );
  DFF_X1 \data_out_reg[3]  ( .D(n181), .CK(clk), .Q(data_out[3]), .QN(n188) );
  DFF_X1 \data_out_reg[2]  ( .D(n182), .CK(clk), .Q(data_out[2]), .QN(n187) );
  DFF_X1 \data_out_reg[1]  ( .D(n183), .CK(clk), .Q(data_out[1]), .QN(n186) );
  DFF_X1 \data_out_reg[0]  ( .D(n184), .CK(clk), .Q(data_out[0]), .QN(n185) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_10_DW_mult_tc_1 mult_960 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_10_DW01_add_2 add_961 ( .A({n207, 
        n206, n205, n204, n203, n202, n216, n215, n214, n213, n212, n211, n210, 
        n209, n208, n201}), .B({f[15], n49, n50, n51, n52, n54, f[9:3], n62, 
        n64, n66}), .CI(1'b0), .SUM(adder) );
  DFF_X1 \f_reg[3]  ( .D(n114), .CK(clk), .Q(f[3]), .QN(n70) );
  DFF_X1 \f_reg[2]  ( .D(n115), .CK(clk), .Q(n62), .QN(n219) );
  DFF_X1 \f_reg[0]  ( .D(n168), .CK(clk), .Q(n66), .QN(n217) );
  DFF_X1 \f_reg[1]  ( .D(n116), .CK(clk), .Q(n64), .QN(n218) );
  DFF_X1 \f_reg[4]  ( .D(n113), .CK(clk), .Q(f[4]), .QN(n71) );
  DFF_X1 \f_reg[5]  ( .D(n104), .CK(clk), .Q(f[5]), .QN(n72) );
  DFF_X1 \f_reg[6]  ( .D(n87), .CK(clk), .Q(f[6]), .QN(n73) );
  DFF_X2 delay_reg ( .D(N27), .CK(clk), .Q(n2), .QN(n244) );
  MUX2_X2 U3 ( .A(n33), .B(N40), .S(n244), .Z(n203) );
  AND2_X2 U4 ( .A1(n48), .A2(n23), .ZN(n19) );
  MUX2_X2 U5 ( .A(n36), .B(N37), .S(n244), .Z(n215) );
  MUX2_X2 U6 ( .A(n29), .B(N42), .S(n244), .Z(n205) );
  MUX2_X2 U8 ( .A(N41), .B(n32), .S(n2), .Z(n204) );
  NAND3_X1 U9 ( .A1(n10), .A2(n9), .A3(n11), .ZN(n1) );
  MUX2_X2 U10 ( .A(N39), .B(n34), .S(n2), .Z(n202) );
  MUX2_X1 U11 ( .A(N38), .B(n35), .S(n2), .Z(n216) );
  NAND3_X1 U12 ( .A1(n7), .A2(n6), .A3(n8), .ZN(n4) );
  NAND3_X1 U13 ( .A1(n17), .A2(n16), .A3(n18), .ZN(n5) );
  NAND2_X1 U14 ( .A1(data_out_b[13]), .A2(n22), .ZN(n6) );
  NAND2_X1 U15 ( .A1(adder[13]), .A2(n19), .ZN(n7) );
  NAND2_X1 U16 ( .A1(n68), .A2(n50), .ZN(n8) );
  NAND2_X1 U17 ( .A1(data_out_b[12]), .A2(n22), .ZN(n9) );
  NAND2_X1 U18 ( .A1(adder[12]), .A2(n19), .ZN(n10) );
  NAND2_X1 U19 ( .A1(n68), .A2(n51), .ZN(n11) );
  AND2_X1 U20 ( .A1(n15), .A2(n13), .ZN(n12) );
  NAND2_X1 U21 ( .A1(n14), .A2(n12), .ZN(n80) );
  NAND2_X1 U22 ( .A1(data_out_b[15]), .A2(n22), .ZN(n13) );
  NAND2_X1 U23 ( .A1(adder[15]), .A2(n19), .ZN(n14) );
  NAND2_X1 U24 ( .A1(n68), .A2(f[15]), .ZN(n15) );
  INV_X2 U25 ( .A(n48), .ZN(n68) );
  NAND2_X1 U26 ( .A1(data_out_b[14]), .A2(n22), .ZN(n16) );
  NAND2_X1 U27 ( .A1(adder[14]), .A2(n19), .ZN(n17) );
  NAND2_X1 U28 ( .A1(n68), .A2(n49), .ZN(n18) );
  INV_X1 U29 ( .A(n23), .ZN(n22) );
  INV_X1 U30 ( .A(clear_acc), .ZN(n23) );
  NAND2_X1 U31 ( .A1(n21), .A2(N27), .ZN(n246) );
  OAI22_X1 U32 ( .A1(n188), .A2(n246), .B1(n70), .B2(n245), .ZN(n181) );
  OAI22_X1 U33 ( .A1(n189), .A2(n246), .B1(n71), .B2(n245), .ZN(n180) );
  OAI22_X1 U34 ( .A1(n190), .A2(n246), .B1(n72), .B2(n245), .ZN(n179) );
  OAI22_X1 U35 ( .A1(n191), .A2(n246), .B1(n73), .B2(n245), .ZN(n178) );
  OAI22_X1 U36 ( .A1(n192), .A2(n246), .B1(n220), .B2(n245), .ZN(n177) );
  OAI22_X1 U37 ( .A1(n193), .A2(n246), .B1(n221), .B2(n245), .ZN(n176) );
  OAI22_X1 U38 ( .A1(n194), .A2(n246), .B1(n222), .B2(n245), .ZN(n175) );
  INV_X1 U39 ( .A(n26), .ZN(n44) );
  MUX2_X1 U40 ( .A(n41), .B(N32), .S(n244), .Z(n210) );
  CLKBUF_X1 U41 ( .A(N42), .Z(n20) );
  INV_X1 U42 ( .A(wr_en_y), .ZN(n21) );
  AND2_X1 U43 ( .A1(sel[0]), .A2(sel[1]), .ZN(n25) );
  INV_X1 U44 ( .A(m_ready), .ZN(n24) );
  NAND2_X1 U45 ( .A1(m_valid), .A2(n24), .ZN(n46) );
  OAI211_X1 U46 ( .C1(sel[2]), .C2(n25), .A(sel[3]), .B(n46), .ZN(N27) );
  NAND2_X1 U47 ( .A1(clear_acc_delay), .A2(n244), .ZN(n26) );
  MUX2_X1 U48 ( .A(n27), .B(N44), .S(n44), .Z(n228) );
  MUX2_X1 U49 ( .A(n27), .B(N44), .S(n244), .Z(n207) );
  MUX2_X1 U50 ( .A(n28), .B(N43), .S(n44), .Z(n229) );
  MUX2_X1 U51 ( .A(n28), .B(N43), .S(n244), .Z(n206) );
  MUX2_X1 U52 ( .A(n29), .B(n20), .S(n44), .Z(n230) );
  MUX2_X1 U53 ( .A(n32), .B(N41), .S(n44), .Z(n231) );
  MUX2_X1 U54 ( .A(n33), .B(N40), .S(n44), .Z(n232) );
  MUX2_X1 U55 ( .A(n34), .B(N39), .S(n44), .Z(n233) );
  MUX2_X1 U56 ( .A(n35), .B(N38), .S(n44), .Z(n234) );
  MUX2_X1 U57 ( .A(n36), .B(N37), .S(n44), .Z(n235) );
  MUX2_X1 U58 ( .A(n37), .B(N36), .S(n44), .Z(n236) );
  MUX2_X1 U59 ( .A(n37), .B(N36), .S(n244), .Z(n214) );
  MUX2_X1 U60 ( .A(n38), .B(N35), .S(n44), .Z(n237) );
  MUX2_X1 U61 ( .A(n38), .B(N35), .S(n244), .Z(n213) );
  MUX2_X1 U62 ( .A(n39), .B(N34), .S(n44), .Z(n238) );
  MUX2_X1 U63 ( .A(n39), .B(N34), .S(n244), .Z(n212) );
  MUX2_X1 U64 ( .A(n40), .B(N33), .S(n44), .Z(n239) );
  MUX2_X1 U65 ( .A(n40), .B(N33), .S(n244), .Z(n211) );
  MUX2_X1 U66 ( .A(n41), .B(N32), .S(n44), .Z(n240) );
  MUX2_X1 U67 ( .A(n42), .B(N31), .S(n44), .Z(n241) );
  MUX2_X1 U68 ( .A(n42), .B(N31), .S(n244), .Z(n209) );
  MUX2_X1 U69 ( .A(n43), .B(N30), .S(n44), .Z(n242) );
  MUX2_X1 U70 ( .A(n43), .B(N30), .S(n244), .Z(n208) );
  MUX2_X1 U71 ( .A(n45), .B(N29), .S(n44), .Z(n243) );
  MUX2_X1 U72 ( .A(n45), .B(N29), .S(n244), .Z(n201) );
  INV_X1 U73 ( .A(n46), .ZN(n47) );
  OAI21_X1 U74 ( .B1(n47), .B2(n2), .A(n23), .ZN(n48) );
  AOI222_X1 U75 ( .A1(data_out_b[11]), .A2(n22), .B1(adder[11]), .B2(n19), 
        .C1(n68), .C2(n52), .ZN(n53) );
  INV_X1 U76 ( .A(n53), .ZN(n81) );
  AOI222_X1 U77 ( .A1(data_out_b[10]), .A2(n22), .B1(adder[10]), .B2(n19), 
        .C1(n68), .C2(n54), .ZN(n55) );
  INV_X1 U78 ( .A(n55), .ZN(n82) );
  AOI222_X1 U79 ( .A1(data_out_b[8]), .A2(n22), .B1(adder[8]), .B2(n19), .C1(
        n68), .C2(f[8]), .ZN(n56) );
  INV_X1 U80 ( .A(n56), .ZN(n84) );
  AOI222_X1 U81 ( .A1(data_out_b[7]), .A2(n22), .B1(adder[7]), .B2(n19), .C1(
        n68), .C2(f[7]), .ZN(n57) );
  INV_X1 U82 ( .A(n57), .ZN(n85) );
  AOI222_X1 U83 ( .A1(data_out_b[6]), .A2(n22), .B1(adder[6]), .B2(n19), .C1(
        n68), .C2(f[6]), .ZN(n58) );
  INV_X1 U84 ( .A(n58), .ZN(n87) );
  AOI222_X1 U85 ( .A1(data_out_b[5]), .A2(n22), .B1(adder[5]), .B2(n19), .C1(
        n68), .C2(f[5]), .ZN(n59) );
  INV_X1 U86 ( .A(n59), .ZN(n104) );
  AOI222_X1 U87 ( .A1(data_out_b[4]), .A2(n22), .B1(adder[4]), .B2(n19), .C1(
        n68), .C2(f[4]), .ZN(n60) );
  INV_X1 U88 ( .A(n60), .ZN(n113) );
  AOI222_X1 U89 ( .A1(data_out_b[3]), .A2(n22), .B1(adder[3]), .B2(n19), .C1(
        n68), .C2(f[3]), .ZN(n61) );
  INV_X1 U90 ( .A(n61), .ZN(n114) );
  AOI222_X1 U91 ( .A1(data_out_b[2]), .A2(n22), .B1(adder[2]), .B2(n19), .C1(
        n68), .C2(n62), .ZN(n63) );
  INV_X1 U92 ( .A(n63), .ZN(n115) );
  AOI222_X1 U93 ( .A1(data_out_b[1]), .A2(n22), .B1(adder[1]), .B2(n19), .C1(
        n68), .C2(n64), .ZN(n65) );
  INV_X1 U94 ( .A(n65), .ZN(n116) );
  AOI222_X1 U95 ( .A1(data_out_b[0]), .A2(n22), .B1(adder[0]), .B2(n19), .C1(
        n68), .C2(n66), .ZN(n67) );
  INV_X1 U96 ( .A(n67), .ZN(n168) );
  AOI222_X1 U97 ( .A1(data_out_b[9]), .A2(n22), .B1(adder[9]), .B2(n19), .C1(
        n68), .C2(f[9]), .ZN(n69) );
  INV_X1 U98 ( .A(n69), .ZN(n83) );
  NOR4_X1 U99 ( .A1(n52), .A2(n51), .A3(n50), .A4(n49), .ZN(n77) );
  NOR4_X1 U100 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n54), .ZN(n76) );
  NAND4_X1 U101 ( .A1(n73), .A2(n72), .A3(n71), .A4(n70), .ZN(n74) );
  NOR4_X1 U102 ( .A1(n74), .A2(n66), .A3(n64), .A4(n62), .ZN(n75) );
  NAND3_X1 U103 ( .A1(n77), .A2(n76), .A3(n75), .ZN(n79) );
  NAND3_X1 U104 ( .A1(wr_en_y), .A2(n79), .A3(n78), .ZN(n245) );
  OAI22_X1 U105 ( .A1(n185), .A2(n246), .B1(n217), .B2(n245), .ZN(n184) );
  OAI22_X1 U106 ( .A1(n186), .A2(n246), .B1(n218), .B2(n245), .ZN(n183) );
  OAI22_X1 U107 ( .A1(n187), .A2(n246), .B1(n219), .B2(n245), .ZN(n182) );
  OAI22_X1 U108 ( .A1(n195), .A2(n246), .B1(n223), .B2(n245), .ZN(n174) );
  OAI22_X1 U109 ( .A1(n196), .A2(n246), .B1(n224), .B2(n245), .ZN(n173) );
  OAI22_X1 U110 ( .A1(n197), .A2(n246), .B1(n225), .B2(n245), .ZN(n172) );
  OAI22_X1 U111 ( .A1(n198), .A2(n246), .B1(n226), .B2(n245), .ZN(n171) );
  OAI22_X1 U112 ( .A1(n199), .A2(n246), .B1(n227), .B2(n245), .ZN(n170) );
  OAI22_X1 U113 ( .A1(n200), .A2(n246), .B1(n78), .B2(n245), .ZN(n169) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_9_DW_mult_tc_1 ( a, b, 
        product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n9, n12, n13, n16, n18, n19, n21, n25, n27, n29, n31, n32,
         n34, n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n62, n63, n64, n65, n67, n69,
         n70, n72, n73, n74, n75, n76, n77, n78, n79, n80, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n93, n95, n96, n97, n98, n99, n101,
         n103, n104, n105, n106, n107, n109, n111, n112, n113, n114, n115,
         n117, n119, n120, n122, n125, n127, n135, n139, n141, n142, n143,
         n144, n145, n147, n148, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n237, n247, n249, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n418, n419,
         n420, n421, n422, n423, n424, n426, n427, n428, n433, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U148 ( .A(n265), .B(n144), .Z(n145) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U161 ( .A(n177), .B(n168), .CI(n166), .CO(n163), .S(n164) );
  FA_X1 U162 ( .A(n170), .B(n172), .CI(n179), .CO(n165), .S(n166) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n263), .CI(n291), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n317), .B(n252), .CO(n173), .S(n174) );
  FA_X1 U167 ( .A(n180), .B(n187), .CI(n178), .CO(n175), .S(n176) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U170 ( .A(n268), .B(n292), .CI(n274), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U174 ( .A(n275), .B(n293), .CI(n194), .CO(n189), .S(n190) );
  HA_X1 U176 ( .A(n269), .B(n319), .CO(n193), .S(n194) );
  FA_X1 U177 ( .A(n205), .B(n200), .CI(n198), .CO(n195), .S(n196) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U179 ( .A(n276), .B(n284), .CI(n294), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n306), .B(n270), .CI(n320), .CO(n201), .S(n202) );
  FA_X1 U181 ( .A(n208), .B(n213), .CI(n206), .CO(n203), .S(n204) );
  FA_X1 U182 ( .A(n210), .B(n307), .CI(n215), .CO(n205), .S(n206) );
  FA_X1 U183 ( .A(n295), .B(n285), .CI(n254), .CO(n207), .S(n208) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U185 ( .A(n216), .B(n219), .CI(n214), .CO(n211), .S(n212) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n322), .B(n278), .CI(n308), .CO(n215), .S(n216) );
  FA_X1 U188 ( .A(n225), .B(n222), .CI(n220), .CO(n217), .S(n218) );
  FA_X1 U189 ( .A(n255), .B(n309), .CI(n297), .CO(n219), .S(n220) );
  HA_X1 U190 ( .A(n287), .B(n323), .CO(n221), .S(n222) );
  FA_X1 U192 ( .A(n324), .B(n288), .CI(n310), .CO(n225), .S(n226) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  HA_X1 U194 ( .A(n325), .B(n311), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n326), .B(n300), .CI(n312), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  OR2_X1 U414 ( .A1(n196), .A2(n203), .ZN(n490) );
  OR2_X1 U415 ( .A1(n218), .A2(n223), .ZN(n491) );
  BUF_X1 U416 ( .A(n1), .Z(n492) );
  OR2_X1 U417 ( .A1(n176), .A2(n185), .ZN(n493) );
  INV_X1 U418 ( .A(n493), .ZN(n494) );
  NOR2_X1 U419 ( .A1(n176), .A2(n185), .ZN(n78) );
  XNOR2_X1 U420 ( .A(n599), .B(a[12]), .ZN(n37) );
  INV_X1 U421 ( .A(n531), .ZN(n73) );
  OR2_X1 U422 ( .A1(n329), .A2(n258), .ZN(n495) );
  BUF_X1 U423 ( .A(n104), .Z(n540) );
  BUF_X1 U424 ( .A(n96), .Z(n550) );
  OR2_X1 U425 ( .A1(n228), .A2(n231), .ZN(n496) );
  XOR2_X1 U426 ( .A(n602), .B(a[14]), .Z(n41) );
  XNOR2_X1 U427 ( .A(n602), .B(a[12]), .ZN(n427) );
  INV_X1 U428 ( .A(n602), .ZN(n601) );
  INV_X2 U429 ( .A(n591), .ZN(n589) );
  BUF_X2 U430 ( .A(n12), .Z(n528) );
  OR2_X2 U431 ( .A1(n554), .A2(n570), .ZN(n500) );
  XNOR2_X1 U432 ( .A(n591), .B(a[4]), .ZN(n556) );
  XNOR2_X1 U433 ( .A(n594), .B(a[6]), .ZN(n497) );
  INV_X1 U434 ( .A(n497), .ZN(n498) );
  INV_X1 U435 ( .A(n497), .ZN(n21) );
  OR2_X1 U436 ( .A1(n75), .A2(n78), .ZN(n531) );
  OR2_X2 U437 ( .A1(n499), .A2(n557), .ZN(n29) );
  XOR2_X1 U438 ( .A(n598), .B(a[8]), .Z(n499) );
  OR2_X1 U439 ( .A1(n554), .A2(n570), .ZN(n526) );
  BUF_X1 U440 ( .A(n12), .Z(n527) );
  BUF_X4 U441 ( .A(n9), .Z(n582) );
  XNOR2_X1 U442 ( .A(n226), .B(n501), .ZN(n224) );
  XNOR2_X1 U443 ( .A(n229), .B(n298), .ZN(n501) );
  INV_X1 U444 ( .A(n556), .ZN(n502) );
  XOR2_X1 U445 ( .A(n594), .B(a[4]), .Z(n541) );
  INV_X1 U446 ( .A(n594), .ZN(n592) );
  XNOR2_X1 U447 ( .A(n503), .B(n147), .ZN(n144) );
  XNOR2_X1 U448 ( .A(n301), .B(n148), .ZN(n503) );
  INV_X1 U449 ( .A(n591), .ZN(n590) );
  OR2_X1 U450 ( .A1(n541), .A2(n556), .ZN(n522) );
  XOR2_X1 U451 ( .A(n199), .B(n201), .Z(n504) );
  XOR2_X1 U452 ( .A(n504), .B(n192), .Z(n188) );
  XOR2_X1 U453 ( .A(n197), .B(n190), .Z(n505) );
  XOR2_X1 U454 ( .A(n505), .B(n188), .Z(n186) );
  NAND2_X1 U455 ( .A1(n199), .A2(n201), .ZN(n506) );
  NAND2_X1 U456 ( .A1(n199), .A2(n192), .ZN(n507) );
  NAND2_X1 U457 ( .A1(n201), .A2(n192), .ZN(n508) );
  NAND3_X1 U458 ( .A1(n506), .A2(n507), .A3(n508), .ZN(n187) );
  NAND2_X1 U459 ( .A1(n197), .A2(n190), .ZN(n509) );
  NAND2_X1 U460 ( .A1(n197), .A2(n188), .ZN(n510) );
  NAND2_X1 U461 ( .A1(n190), .A2(n188), .ZN(n511) );
  NAND3_X1 U462 ( .A1(n509), .A2(n510), .A3(n511), .ZN(n185) );
  XOR2_X1 U463 ( .A(n283), .B(n253), .Z(n512) );
  XOR2_X1 U464 ( .A(n305), .B(n512), .Z(n192) );
  NAND2_X1 U465 ( .A1(n305), .A2(n283), .ZN(n513) );
  NAND2_X1 U466 ( .A1(n305), .A2(n253), .ZN(n514) );
  NAND2_X1 U467 ( .A1(n283), .A2(n253), .ZN(n515) );
  NAND3_X1 U468 ( .A1(n513), .A2(n514), .A3(n515), .ZN(n191) );
  XNOR2_X1 U469 ( .A(n492), .B(a[2]), .ZN(n9) );
  XOR2_X1 U470 ( .A(n193), .B(n282), .Z(n516) );
  XOR2_X1 U471 ( .A(n191), .B(n516), .Z(n180) );
  NAND2_X1 U472 ( .A1(n191), .A2(n193), .ZN(n517) );
  NAND2_X1 U473 ( .A1(n191), .A2(n282), .ZN(n518) );
  NAND2_X1 U474 ( .A1(n193), .A2(n282), .ZN(n519) );
  NAND3_X1 U475 ( .A1(n517), .A2(n518), .A3(n519), .ZN(n179) );
  NAND2_X1 U476 ( .A1(n428), .A2(n32), .ZN(n34) );
  BUF_X1 U477 ( .A(n586), .Z(n520) );
  INV_X1 U478 ( .A(n598), .ZN(n521) );
  INV_X1 U479 ( .A(n598), .ZN(n597) );
  XNOR2_X1 U480 ( .A(n591), .B(a[2]), .ZN(n571) );
  OR2_X2 U481 ( .A1(n541), .A2(n556), .ZN(n523) );
  OR2_X1 U482 ( .A1(n541), .A2(n556), .ZN(n18) );
  XNOR2_X1 U483 ( .A(n271), .B(n524), .ZN(n147) );
  XNOR2_X1 U484 ( .A(n289), .B(n279), .ZN(n524) );
  INV_X1 U485 ( .A(n589), .ZN(n525) );
  XNOR2_X1 U486 ( .A(n600), .B(a[10]), .ZN(n428) );
  BUF_X2 U487 ( .A(n12), .Z(n529) );
  NAND2_X1 U488 ( .A1(n571), .A2(n9), .ZN(n12) );
  XOR2_X1 U489 ( .A(n586), .B(n249), .Z(n530) );
  BUF_X2 U490 ( .A(n32), .Z(n532) );
  INV_X1 U491 ( .A(n559), .ZN(n32) );
  INV_X1 U492 ( .A(n543), .ZN(n533) );
  INV_X2 U493 ( .A(n596), .ZN(n543) );
  OR2_X1 U494 ( .A1(n204), .A2(n211), .ZN(n534) );
  BUF_X2 U495 ( .A(n585), .Z(n535) );
  INV_X1 U496 ( .A(n249), .ZN(n585) );
  NOR2_X1 U497 ( .A1(n186), .A2(n195), .ZN(n536) );
  NOR2_X1 U498 ( .A1(n186), .A2(n195), .ZN(n82) );
  INV_X1 U499 ( .A(n587), .ZN(n537) );
  CLKBUF_X1 U500 ( .A(n569), .Z(n551) );
  CLKBUF_X1 U501 ( .A(n74), .Z(n538) );
  BUF_X1 U502 ( .A(n568), .Z(n539) );
  INV_X1 U503 ( .A(n556), .ZN(n16) );
  AOI21_X1 U504 ( .B1(n96), .B2(n573), .A(n93), .ZN(n542) );
  INV_X1 U505 ( .A(n596), .ZN(n544) );
  INV_X1 U506 ( .A(n596), .ZN(n595) );
  CLKBUF_X1 U507 ( .A(n539), .Z(n545) );
  NOR2_X1 U508 ( .A1(n164), .A2(n175), .ZN(n546) );
  NAND2_X1 U509 ( .A1(n427), .A2(n37), .ZN(n547) );
  INV_X1 U510 ( .A(n600), .ZN(n548) );
  INV_X1 U511 ( .A(n600), .ZN(n549) );
  NOR2_X1 U512 ( .A1(n164), .A2(n175), .ZN(n75) );
  INV_X1 U513 ( .A(n600), .ZN(n599) );
  OAI21_X1 U514 ( .B1(n91), .B2(n89), .A(n90), .ZN(n552) );
  OAI21_X1 U515 ( .B1(n542), .B2(n89), .A(n90), .ZN(n88) );
  CLKBUF_X1 U516 ( .A(n107), .Z(n553) );
  XNOR2_X1 U517 ( .A(n595), .B(a[6]), .ZN(n554) );
  OAI21_X1 U518 ( .B1(n82), .B2(n86), .A(n83), .ZN(n555) );
  INV_X1 U519 ( .A(n557), .ZN(n27) );
  XNOR2_X1 U520 ( .A(n596), .B(a[8]), .ZN(n557) );
  XNOR2_X1 U521 ( .A(n558), .B(n45), .ZN(product[12]) );
  AND2_X1 U522 ( .A1(n493), .A2(n79), .ZN(n558) );
  INV_X1 U523 ( .A(n588), .ZN(n586) );
  INV_X2 U524 ( .A(n588), .ZN(n587) );
  XNOR2_X1 U525 ( .A(n598), .B(a[10]), .ZN(n559) );
  OAI21_X1 U526 ( .B1(n113), .B2(n115), .A(n114), .ZN(n560) );
  AOI21_X1 U527 ( .B1(n578), .B2(n540), .A(n101), .ZN(n561) );
  XNOR2_X1 U528 ( .A(n552), .B(n51), .ZN(product[10]) );
  NAND2_X1 U529 ( .A1(n226), .A2(n229), .ZN(n562) );
  NAND2_X1 U530 ( .A1(n226), .A2(n298), .ZN(n563) );
  NAND2_X1 U531 ( .A1(n229), .A2(n298), .ZN(n564) );
  NAND3_X1 U532 ( .A1(n562), .A2(n563), .A3(n564), .ZN(n223) );
  NOR2_X1 U533 ( .A1(n567), .A2(n403), .ZN(n565) );
  NOR2_X1 U534 ( .A1(n402), .A2(n585), .ZN(n566) );
  OR2_X1 U535 ( .A1(n565), .A2(n566), .ZN(n324) );
  NAND2_X1 U536 ( .A1(n433), .A2(n585), .ZN(n567) );
  NAND2_X1 U537 ( .A1(n530), .A2(n585), .ZN(n568) );
  AOI21_X1 U538 ( .B1(n80), .B2(n88), .A(n555), .ZN(n569) );
  XNOR2_X1 U539 ( .A(n594), .B(a[6]), .ZN(n570) );
  BUF_X1 U540 ( .A(n43), .Z(n583) );
  NAND2_X1 U541 ( .A1(n572), .A2(n69), .ZN(n47) );
  INV_X1 U542 ( .A(n69), .ZN(n67) );
  NAND2_X1 U543 ( .A1(n73), .A2(n572), .ZN(n64) );
  INV_X1 U544 ( .A(n74), .ZN(n72) );
  AOI21_X1 U545 ( .B1(n96), .B2(n573), .A(n93), .ZN(n91) );
  INV_X1 U546 ( .A(n95), .ZN(n93) );
  NAND2_X1 U547 ( .A1(n127), .A2(n83), .ZN(n50) );
  INV_X1 U548 ( .A(n536), .ZN(n127) );
  NAND2_X1 U549 ( .A1(n490), .A2(n86), .ZN(n51) );
  OR2_X1 U550 ( .A1(n152), .A2(n163), .ZN(n572) );
  NAND2_X1 U551 ( .A1(n573), .A2(n95), .ZN(n53) );
  NAND2_X1 U552 ( .A1(n125), .A2(n76), .ZN(n48) );
  INV_X1 U553 ( .A(n75), .ZN(n125) );
  OAI21_X1 U554 ( .B1(n546), .B2(n79), .A(n76), .ZN(n74) );
  AOI21_X1 U555 ( .B1(n80), .B2(n552), .A(n555), .ZN(n45) );
  NOR2_X1 U556 ( .A1(n536), .A2(n85), .ZN(n80) );
  NAND2_X1 U557 ( .A1(n152), .A2(n163), .ZN(n69) );
  NAND2_X1 U558 ( .A1(n534), .A2(n90), .ZN(n52) );
  OAI21_X1 U559 ( .B1(n115), .B2(n113), .A(n114), .ZN(n112) );
  NAND2_X1 U560 ( .A1(n496), .A2(n106), .ZN(n56) );
  NAND2_X1 U561 ( .A1(n135), .A2(n114), .ZN(n58) );
  NAND2_X1 U562 ( .A1(n491), .A2(n98), .ZN(n54) );
  AOI21_X1 U563 ( .B1(n577), .B2(n112), .A(n109), .ZN(n107) );
  INV_X1 U564 ( .A(n111), .ZN(n109) );
  NOR2_X1 U565 ( .A1(n196), .A2(n203), .ZN(n85) );
  NAND2_X1 U566 ( .A1(n576), .A2(n62), .ZN(n46) );
  AOI21_X1 U567 ( .B1(n538), .B2(n572), .A(n67), .ZN(n65) );
  AOI21_X1 U568 ( .B1(n575), .B2(n120), .A(n117), .ZN(n115) );
  INV_X1 U569 ( .A(n119), .ZN(n117) );
  INV_X1 U570 ( .A(n122), .ZN(n120) );
  NOR2_X1 U571 ( .A1(n204), .A2(n211), .ZN(n89) );
  XNOR2_X1 U572 ( .A(n55), .B(n540), .ZN(product[6]) );
  XNOR2_X1 U573 ( .A(n57), .B(n560), .ZN(product[4]) );
  NAND2_X1 U574 ( .A1(n577), .A2(n111), .ZN(n57) );
  NAND2_X1 U575 ( .A1(n176), .A2(n185), .ZN(n79) );
  NAND2_X1 U576 ( .A1(n196), .A2(n203), .ZN(n86) );
  NAND2_X1 U577 ( .A1(n164), .A2(n175), .ZN(n76) );
  NAND2_X1 U578 ( .A1(n186), .A2(n195), .ZN(n83) );
  OR2_X1 U579 ( .A1(n212), .A2(n217), .ZN(n573) );
  NAND2_X1 U580 ( .A1(n204), .A2(n211), .ZN(n90) );
  NAND2_X1 U581 ( .A1(n212), .A2(n217), .ZN(n95) );
  XNOR2_X1 U582 ( .A(n59), .B(n120), .ZN(product[2]) );
  NAND2_X1 U583 ( .A1(n575), .A2(n119), .ZN(n59) );
  AND2_X1 U584 ( .A1(n495), .A2(n122), .ZN(product[1]) );
  OR2_X1 U585 ( .A1(n328), .A2(n314), .ZN(n575) );
  OR2_X1 U586 ( .A1(n151), .A2(n139), .ZN(n576) );
  NOR2_X1 U587 ( .A1(n218), .A2(n223), .ZN(n97) );
  NAND2_X1 U588 ( .A1(n218), .A2(n223), .ZN(n98) );
  OR2_X1 U589 ( .A1(n232), .A2(n233), .ZN(n577) );
  INV_X1 U590 ( .A(n37), .ZN(n237) );
  OR2_X1 U591 ( .A1(n224), .A2(n227), .ZN(n578) );
  INV_X1 U592 ( .A(n41), .ZN(n235) );
  OR2_X1 U593 ( .A1(n583), .A2(n525), .ZN(n392) );
  AND2_X1 U594 ( .A1(n584), .A2(n559), .ZN(n270) );
  XNOR2_X1 U595 ( .A(n521), .B(n583), .ZN(n352) );
  XNOR2_X1 U596 ( .A(n589), .B(n583), .ZN(n391) );
  XNOR2_X1 U597 ( .A(n155), .B(n579), .ZN(n139) );
  XNOR2_X1 U598 ( .A(n153), .B(n141), .ZN(n579) );
  XNOR2_X1 U599 ( .A(n157), .B(n580), .ZN(n141) );
  XNOR2_X1 U600 ( .A(n145), .B(n143), .ZN(n580) );
  OAI22_X1 U601 ( .A1(n547), .A2(n602), .B1(n337), .B2(n37), .ZN(n252) );
  OR2_X1 U602 ( .A1(n583), .A2(n602), .ZN(n337) );
  NAND2_X1 U603 ( .A1(n433), .A2(n585), .ZN(n6) );
  OAI22_X1 U604 ( .A1(n42), .A2(n604), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U605 ( .A1(n583), .A2(n604), .ZN(n332) );
  XNOR2_X1 U606 ( .A(n549), .B(n583), .ZN(n343) );
  AND2_X1 U607 ( .A1(n584), .A2(n556), .ZN(n300) );
  XNOR2_X1 U608 ( .A(n159), .B(n581), .ZN(n142) );
  XNOR2_X1 U609 ( .A(n315), .B(n261), .ZN(n581) );
  XNOR2_X1 U610 ( .A(n601), .B(n583), .ZN(n336) );
  NAND2_X1 U611 ( .A1(n427), .A2(n37), .ZN(n39) );
  OAI22_X1 U612 ( .A1(n39), .A2(n336), .B1(n37), .B2(n335), .ZN(n263) );
  XNOR2_X1 U613 ( .A(n593), .B(n583), .ZN(n376) );
  AND2_X1 U614 ( .A1(n584), .A2(n237), .ZN(n264) );
  AND2_X1 U615 ( .A1(n584), .A2(n497), .ZN(n288) );
  AND2_X1 U616 ( .A1(n584), .A2(n235), .ZN(n260) );
  OAI22_X1 U617 ( .A1(n39), .A2(n335), .B1(n37), .B2(n334), .ZN(n262) );
  INV_X1 U618 ( .A(n25), .ZN(n598) );
  AND2_X1 U619 ( .A1(n584), .A2(n557), .ZN(n278) );
  NAND2_X1 U620 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U621 ( .A(n603), .B(a[14]), .Z(n426) );
  INV_X1 U622 ( .A(n13), .ZN(n594) );
  AND2_X1 U623 ( .A1(n584), .A2(n247), .ZN(n314) );
  AND2_X1 U624 ( .A1(n584), .A2(n249), .ZN(product[0]) );
  OR2_X1 U625 ( .A1(n583), .A2(n600), .ZN(n344) );
  OR2_X1 U626 ( .A1(n583), .A2(n598), .ZN(n353) );
  OR2_X1 U627 ( .A1(n583), .A2(n533), .ZN(n364) );
  OR2_X1 U628 ( .A1(n583), .A2(n594), .ZN(n377) );
  OAI22_X1 U629 ( .A1(n547), .A2(n334), .B1(n37), .B2(n333), .ZN(n261) );
  XNOR2_X1 U630 ( .A(n601), .B(n422), .ZN(n333) );
  XNOR2_X1 U631 ( .A(n593), .B(b[11]), .ZN(n365) );
  XNOR2_X1 U632 ( .A(n601), .B(n424), .ZN(n335) );
  XNOR2_X1 U633 ( .A(n601), .B(n423), .ZN(n334) );
  OAI22_X1 U634 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U635 ( .A(n603), .B(n424), .ZN(n330) );
  XNOR2_X1 U636 ( .A(n603), .B(n583), .ZN(n331) );
  XNOR2_X1 U637 ( .A(n521), .B(n418), .ZN(n345) );
  XNOR2_X1 U638 ( .A(n548), .B(n420), .ZN(n338) );
  XNOR2_X1 U639 ( .A(n589), .B(b[13]), .ZN(n378) );
  XNOR2_X1 U640 ( .A(n589), .B(n424), .ZN(n390) );
  XNOR2_X1 U641 ( .A(n597), .B(n424), .ZN(n351) );
  XNOR2_X1 U642 ( .A(n549), .B(n424), .ZN(n342) );
  XNOR2_X1 U643 ( .A(n548), .B(n423), .ZN(n341) );
  XNOR2_X1 U644 ( .A(n548), .B(n422), .ZN(n340) );
  XNOR2_X1 U645 ( .A(n549), .B(n421), .ZN(n339) );
  XNOR2_X1 U646 ( .A(n590), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U647 ( .A(n590), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U648 ( .A(n589), .B(n419), .ZN(n385) );
  XNOR2_X1 U649 ( .A(n590), .B(n418), .ZN(n384) );
  XNOR2_X1 U650 ( .A(n589), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U651 ( .A(n589), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U652 ( .A(n589), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U653 ( .A(n593), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U654 ( .A(n593), .B(n418), .ZN(n369) );
  XNOR2_X1 U655 ( .A(n593), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U656 ( .A(n593), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U657 ( .A(n590), .B(n423), .ZN(n389) );
  XNOR2_X1 U658 ( .A(n597), .B(n423), .ZN(n350) );
  XNOR2_X1 U659 ( .A(n590), .B(n422), .ZN(n388) );
  XNOR2_X1 U660 ( .A(n521), .B(n422), .ZN(n349) );
  XNOR2_X1 U661 ( .A(n587), .B(b[11]), .ZN(n397) );
  XNOR2_X1 U662 ( .A(n587), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U663 ( .A(n587), .B(b[13]), .ZN(n395) );
  XNOR2_X1 U664 ( .A(n587), .B(b[14]), .ZN(n394) );
  XNOR2_X1 U665 ( .A(n589), .B(n420), .ZN(n386) );
  XNOR2_X1 U666 ( .A(n597), .B(n421), .ZN(n348) );
  XNOR2_X1 U667 ( .A(n589), .B(n421), .ZN(n387) );
  XNOR2_X1 U668 ( .A(n521), .B(n420), .ZN(n347) );
  XNOR2_X1 U669 ( .A(n521), .B(n419), .ZN(n346) );
  XNOR2_X1 U670 ( .A(n587), .B(b[15]), .ZN(n393) );
  BUF_X1 U671 ( .A(n43), .Z(n584) );
  OAI22_X1 U672 ( .A1(n34), .A2(n339), .B1(n338), .B2(n532), .ZN(n265) );
  OAI22_X1 U673 ( .A1(n34), .A2(n341), .B1(n340), .B2(n532), .ZN(n267) );
  OAI22_X1 U674 ( .A1(n34), .A2(n340), .B1(n339), .B2(n532), .ZN(n266) );
  OAI22_X1 U675 ( .A1(n34), .A2(n342), .B1(n341), .B2(n532), .ZN(n268) );
  OAI22_X1 U676 ( .A1(n34), .A2(n343), .B1(n342), .B2(n532), .ZN(n269) );
  OAI22_X1 U677 ( .A1(n34), .A2(n600), .B1(n344), .B2(n532), .ZN(n253) );
  NAND2_X1 U678 ( .A1(n328), .A2(n314), .ZN(n119) );
  OAI22_X1 U679 ( .A1(n29), .A2(n350), .B1(n349), .B2(n27), .ZN(n275) );
  OAI22_X1 U680 ( .A1(n29), .A2(n346), .B1(n345), .B2(n27), .ZN(n271) );
  OAI22_X1 U681 ( .A1(n29), .A2(n347), .B1(n346), .B2(n27), .ZN(n272) );
  OAI22_X1 U682 ( .A1(n29), .A2(n348), .B1(n347), .B2(n27), .ZN(n273) );
  OAI22_X1 U683 ( .A1(n29), .A2(n349), .B1(n348), .B2(n27), .ZN(n274) );
  OAI22_X1 U684 ( .A1(n29), .A2(n351), .B1(n350), .B2(n27), .ZN(n276) );
  OAI22_X1 U685 ( .A1(n29), .A2(n598), .B1(n353), .B2(n27), .ZN(n254) );
  OAI22_X1 U686 ( .A1(n29), .A2(n352), .B1(n351), .B2(n27), .ZN(n277) );
  NAND2_X1 U687 ( .A1(n228), .A2(n231), .ZN(n106) );
  NOR2_X1 U688 ( .A1(n228), .A2(n231), .ZN(n105) );
  NAND2_X1 U689 ( .A1(n232), .A2(n233), .ZN(n111) );
  INV_X1 U690 ( .A(n103), .ZN(n101) );
  NAND2_X1 U691 ( .A1(n224), .A2(n227), .ZN(n103) );
  XNOR2_X1 U692 ( .A(n543), .B(n419), .ZN(n357) );
  XNOR2_X1 U693 ( .A(n544), .B(n418), .ZN(n356) );
  XNOR2_X1 U694 ( .A(n544), .B(n422), .ZN(n360) );
  XNOR2_X1 U695 ( .A(n543), .B(b[9]), .ZN(n354) );
  XNOR2_X1 U696 ( .A(n543), .B(n421), .ZN(n359) );
  XNOR2_X1 U697 ( .A(n543), .B(n423), .ZN(n361) );
  XNOR2_X1 U698 ( .A(n544), .B(b[8]), .ZN(n355) );
  INV_X1 U699 ( .A(n19), .ZN(n596) );
  INV_X1 U700 ( .A(n113), .ZN(n135) );
  XNOR2_X1 U701 ( .A(n84), .B(n50), .ZN(product[11]) );
  XNOR2_X1 U702 ( .A(n544), .B(n424), .ZN(n362) );
  XNOR2_X1 U703 ( .A(n543), .B(n583), .ZN(n363) );
  XNOR2_X1 U704 ( .A(n544), .B(n420), .ZN(n358) );
  OAI21_X1 U705 ( .B1(n99), .B2(n97), .A(n98), .ZN(n96) );
  AOI21_X1 U706 ( .B1(n578), .B2(n104), .A(n101), .ZN(n99) );
  XNOR2_X1 U707 ( .A(n63), .B(n46), .ZN(product[15]) );
  INV_X1 U708 ( .A(n7), .ZN(n591) );
  XNOR2_X1 U709 ( .A(n77), .B(n48), .ZN(product[13]) );
  NAND2_X1 U710 ( .A1(n578), .A2(n103), .ZN(n55) );
  XOR2_X1 U711 ( .A(n561), .B(n54), .Z(product[7]) );
  INV_X1 U712 ( .A(n1), .ZN(n588) );
  OR2_X1 U713 ( .A1(n583), .A2(n537), .ZN(n409) );
  OAI22_X1 U714 ( .A1(n500), .A2(n358), .B1(n357), .B2(n498), .ZN(n282) );
  OAI22_X1 U715 ( .A1(n500), .A2(n356), .B1(n355), .B2(n498), .ZN(n280) );
  OAI22_X1 U716 ( .A1(n500), .A2(n362), .B1(n361), .B2(n498), .ZN(n286) );
  OAI22_X1 U717 ( .A1(n500), .A2(n360), .B1(n359), .B2(n498), .ZN(n284) );
  OAI22_X1 U718 ( .A1(n526), .A2(n361), .B1(n360), .B2(n498), .ZN(n285) );
  OAI22_X1 U719 ( .A1(n500), .A2(n357), .B1(n356), .B2(n498), .ZN(n281) );
  OAI22_X1 U720 ( .A1(n500), .A2(n533), .B1(n364), .B2(n21), .ZN(n255) );
  OAI22_X1 U721 ( .A1(n500), .A2(n355), .B1(n354), .B2(n498), .ZN(n279) );
  OAI22_X1 U722 ( .A1(n526), .A2(n363), .B1(n362), .B2(n21), .ZN(n287) );
  OAI22_X1 U723 ( .A1(n526), .A2(n359), .B1(n358), .B2(n21), .ZN(n283) );
  XNOR2_X1 U724 ( .A(n592), .B(n423), .ZN(n374) );
  XNOR2_X1 U725 ( .A(n592), .B(n421), .ZN(n372) );
  XNOR2_X1 U726 ( .A(n592), .B(n422), .ZN(n373) );
  XNOR2_X1 U727 ( .A(n592), .B(n419), .ZN(n370) );
  XNOR2_X1 U728 ( .A(n592), .B(n420), .ZN(n371) );
  XNOR2_X1 U729 ( .A(n592), .B(n424), .ZN(n375) );
  OAI21_X1 U730 ( .B1(n87), .B2(n85), .A(n86), .ZN(n84) );
  XNOR2_X1 U731 ( .A(n550), .B(n53), .ZN(product[8]) );
  XNOR2_X1 U732 ( .A(n587), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U733 ( .A(n587), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U734 ( .A(n587), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U735 ( .A(n587), .B(n418), .ZN(n401) );
  XNOR2_X1 U736 ( .A(n520), .B(n420), .ZN(n403) );
  XNOR2_X1 U737 ( .A(n520), .B(n419), .ZN(n402) );
  XNOR2_X1 U738 ( .A(n587), .B(n583), .ZN(n408) );
  XNOR2_X1 U739 ( .A(n587), .B(n421), .ZN(n404) );
  XNOR2_X1 U740 ( .A(n587), .B(n422), .ZN(n405) );
  XNOR2_X1 U741 ( .A(n587), .B(n424), .ZN(n407) );
  XNOR2_X1 U742 ( .A(n587), .B(n423), .ZN(n406) );
  XOR2_X1 U743 ( .A(n586), .B(n249), .Z(n433) );
  NAND2_X1 U744 ( .A1(n151), .A2(n139), .ZN(n62) );
  OAI22_X1 U745 ( .A1(n523), .A2(n370), .B1(n369), .B2(n502), .ZN(n293) );
  OAI22_X1 U746 ( .A1(n522), .A2(n367), .B1(n366), .B2(n502), .ZN(n290) );
  OAI22_X1 U747 ( .A1(n18), .A2(n368), .B1(n367), .B2(n16), .ZN(n291) );
  OAI22_X1 U748 ( .A1(n522), .A2(n375), .B1(n374), .B2(n502), .ZN(n298) );
  OAI22_X1 U749 ( .A1(n523), .A2(n372), .B1(n371), .B2(n16), .ZN(n295) );
  OAI22_X1 U750 ( .A1(n523), .A2(n373), .B1(n372), .B2(n16), .ZN(n296) );
  OAI22_X1 U751 ( .A1(n18), .A2(n369), .B1(n16), .B2(n368), .ZN(n292) );
  OAI22_X1 U752 ( .A1(n523), .A2(n371), .B1(n370), .B2(n16), .ZN(n294) );
  OAI22_X1 U753 ( .A1(n522), .A2(n374), .B1(n373), .B2(n16), .ZN(n297) );
  OAI22_X1 U754 ( .A1(n522), .A2(n594), .B1(n377), .B2(n502), .ZN(n256) );
  OAI22_X1 U755 ( .A1(n523), .A2(n376), .B1(n375), .B2(n502), .ZN(n299) );
  OAI22_X1 U756 ( .A1(n522), .A2(n366), .B1(n365), .B2(n502), .ZN(n289) );
  OAI21_X1 U757 ( .B1(n64), .B2(n551), .A(n65), .ZN(n63) );
  XNOR2_X1 U758 ( .A(n70), .B(n47), .ZN(product[14]) );
  OAI21_X1 U759 ( .B1(n569), .B2(n494), .A(n79), .ZN(n77) );
  OAI21_X1 U760 ( .B1(n45), .B2(n531), .A(n72), .ZN(n70) );
  XOR2_X1 U761 ( .A(n542), .B(n52), .Z(product[9]) );
  INV_X1 U762 ( .A(n88), .ZN(n87) );
  OAI21_X1 U763 ( .B1(n105), .B2(n107), .A(n106), .ZN(n104) );
  NOR2_X1 U764 ( .A1(n234), .A2(n257), .ZN(n113) );
  XOR2_X1 U765 ( .A(n56), .B(n553), .Z(product[5]) );
  XOR2_X1 U766 ( .A(n58), .B(n115), .Z(product[3]) );
  OAI22_X1 U767 ( .A1(n545), .A2(n395), .B1(n394), .B2(n535), .ZN(n316) );
  OAI22_X1 U768 ( .A1(n545), .A2(n394), .B1(n393), .B2(n535), .ZN(n315) );
  OAI22_X1 U769 ( .A1(n6), .A2(n396), .B1(n395), .B2(n535), .ZN(n317) );
  OAI22_X1 U770 ( .A1(n6), .A2(n397), .B1(n396), .B2(n535), .ZN(n318) );
  OAI22_X1 U771 ( .A1(n568), .A2(n398), .B1(n397), .B2(n535), .ZN(n319) );
  OAI22_X1 U772 ( .A1(n568), .A2(n400), .B1(n399), .B2(n535), .ZN(n321) );
  OAI22_X1 U773 ( .A1(n568), .A2(n399), .B1(n398), .B2(n535), .ZN(n320) );
  OAI22_X1 U774 ( .A1(n6), .A2(n401), .B1(n400), .B2(n535), .ZN(n322) );
  OAI22_X1 U775 ( .A1(n568), .A2(n402), .B1(n401), .B2(n535), .ZN(n323) );
  NAND2_X1 U776 ( .A1(n329), .A2(n258), .ZN(n122) );
  OAI22_X1 U777 ( .A1(n567), .A2(n404), .B1(n403), .B2(n585), .ZN(n325) );
  OAI22_X1 U778 ( .A1(n6), .A2(n406), .B1(n405), .B2(n535), .ZN(n327) );
  OAI22_X1 U779 ( .A1(n567), .A2(n405), .B1(n404), .B2(n585), .ZN(n326) );
  OAI22_X1 U780 ( .A1(n6), .A2(n407), .B1(n406), .B2(n535), .ZN(n328) );
  OAI22_X1 U781 ( .A1(n539), .A2(n408), .B1(n407), .B2(n535), .ZN(n329) );
  OAI22_X1 U782 ( .A1(n6), .A2(n537), .B1(n409), .B2(n535), .ZN(n258) );
  OAI22_X1 U783 ( .A1(n528), .A2(n379), .B1(n378), .B2(n582), .ZN(n301) );
  OAI22_X1 U784 ( .A1(n529), .A2(n380), .B1(n379), .B2(n582), .ZN(n302) );
  OAI22_X1 U785 ( .A1(n528), .A2(n385), .B1(n384), .B2(n582), .ZN(n307) );
  OAI22_X1 U786 ( .A1(n529), .A2(n382), .B1(n381), .B2(n582), .ZN(n304) );
  OAI22_X1 U787 ( .A1(n528), .A2(n381), .B1(n380), .B2(n582), .ZN(n303) );
  NAND2_X1 U788 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U789 ( .A1(n529), .A2(n383), .B1(n582), .B2(n382), .ZN(n305) );
  OAI22_X1 U790 ( .A1(n527), .A2(n384), .B1(n383), .B2(n582), .ZN(n306) );
  OAI22_X1 U791 ( .A1(n528), .A2(n386), .B1(n385), .B2(n582), .ZN(n308) );
  OAI22_X1 U792 ( .A1(n528), .A2(n387), .B1(n386), .B2(n582), .ZN(n309) );
  OAI22_X1 U793 ( .A1(n529), .A2(n525), .B1(n392), .B2(n582), .ZN(n257) );
  OAI22_X1 U794 ( .A1(n527), .A2(n389), .B1(n388), .B2(n582), .ZN(n311) );
  OAI22_X1 U795 ( .A1(n529), .A2(n388), .B1(n387), .B2(n582), .ZN(n310) );
  OAI22_X1 U796 ( .A1(n528), .A2(n390), .B1(n389), .B2(n582), .ZN(n312) );
  INV_X1 U797 ( .A(n582), .ZN(n247) );
  OAI22_X1 U798 ( .A1(n529), .A2(n391), .B1(n390), .B2(n582), .ZN(n313) );
  INV_X1 U799 ( .A(n594), .ZN(n593) );
  INV_X1 U800 ( .A(n31), .ZN(n600) );
  INV_X1 U801 ( .A(n36), .ZN(n602) );
  INV_X1 U802 ( .A(n604), .ZN(n603) );
  INV_X1 U803 ( .A(n40), .ZN(n604) );
  XOR2_X1 U804 ( .A(n259), .B(n251), .Z(n148) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_9_DW01_add_2 ( A, B, CI, SUM, 
        CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n4, n7, n8, n9, n10, n11, n12, n13, n14, n15, n18, n19, n20,
         n21, n25, n26, n27, n28, n30, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n48, n49, n51, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n69, n71, n72, n73, n74, n75,
         n77, n79, n80, n81, n82, n83, n85, n87, n88, n90, n94, n99, n100,
         n102, n104, n161, n162, n163, n164, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189;

  OR2_X1 U126 ( .A1(A[14]), .A2(B[14]), .ZN(n161) );
  OR2_X1 U127 ( .A1(A[14]), .A2(B[14]), .ZN(n162) );
  OR2_X1 U128 ( .A1(A[14]), .A2(B[14]), .ZN(n187) );
  BUF_X1 U129 ( .A(n40), .Z(n163) );
  OR2_X1 U130 ( .A1(A[8]), .A2(B[8]), .ZN(n164) );
  AND2_X1 U131 ( .A1(n182), .A2(n90), .ZN(SUM[0]) );
  OR2_X1 U132 ( .A1(A[15]), .A2(B[15]), .ZN(n166) );
  NOR2_X1 U133 ( .A1(A[8]), .A2(B[8]), .ZN(n167) );
  NOR2_X1 U134 ( .A1(A[8]), .A2(B[8]), .ZN(n58) );
  XNOR2_X1 U135 ( .A(n49), .B(n168), .ZN(SUM[10]) );
  AND2_X1 U136 ( .A1(n188), .A2(n48), .ZN(n168) );
  OR2_X2 U137 ( .A1(A[10]), .A2(B[10]), .ZN(n188) );
  XNOR2_X1 U138 ( .A(n169), .B(n41), .ZN(SUM[11]) );
  AND2_X1 U139 ( .A1(n178), .A2(n40), .ZN(n169) );
  AND2_X1 U140 ( .A1(A[14]), .A2(B[14]), .ZN(n170) );
  OR2_X1 U141 ( .A1(A[13]), .A2(B[13]), .ZN(n171) );
  BUF_X1 U142 ( .A(n179), .Z(n172) );
  AOI21_X1 U143 ( .B1(n56), .B2(n64), .A(n57), .ZN(n173) );
  AOI21_X1 U144 ( .B1(n56), .B2(n64), .A(n57), .ZN(n174) );
  AOI21_X1 U145 ( .B1(n188), .B2(n51), .A(n189), .ZN(n175) );
  OAI21_X1 U146 ( .B1(n43), .B2(n55), .A(n175), .ZN(n176) );
  XNOR2_X1 U147 ( .A(n33), .B(n177), .ZN(SUM[13]) );
  AND2_X1 U148 ( .A1(n171), .A2(n28), .ZN(n177) );
  AOI21_X1 U149 ( .B1(n187), .B2(n30), .A(n170), .ZN(n21) );
  OR2_X1 U150 ( .A1(A[11]), .A2(B[11]), .ZN(n178) );
  NOR2_X1 U151 ( .A1(A[12]), .A2(B[12]), .ZN(n179) );
  NOR2_X1 U152 ( .A1(A[12]), .A2(B[12]), .ZN(n36) );
  OAI21_X1 U153 ( .B1(n179), .B2(n40), .A(n37), .ZN(n180) );
  AOI21_X1 U154 ( .B1(n176), .B2(n34), .A(n35), .ZN(n181) );
  OR2_X1 U155 ( .A1(A[0]), .A2(B[0]), .ZN(n182) );
  INV_X1 U156 ( .A(n64), .ZN(n63) );
  INV_X1 U157 ( .A(n174), .ZN(n54) );
  OAI21_X1 U158 ( .B1(n67), .B2(n65), .A(n66), .ZN(n64) );
  AOI21_X1 U159 ( .B1(n186), .B2(n80), .A(n77), .ZN(n75) );
  INV_X1 U160 ( .A(n79), .ZN(n77) );
  AOI21_X1 U161 ( .B1(n176), .B2(n34), .A(n180), .ZN(n33) );
  AOI21_X1 U162 ( .B1(n185), .B2(n72), .A(n69), .ZN(n67) );
  INV_X1 U163 ( .A(n71), .ZN(n69) );
  AOI21_X1 U164 ( .B1(n184), .B2(n88), .A(n85), .ZN(n83) );
  INV_X1 U165 ( .A(n87), .ZN(n85) );
  OAI21_X1 U166 ( .B1(n83), .B2(n81), .A(n82), .ZN(n80) );
  AOI21_X1 U167 ( .B1(n56), .B2(n64), .A(n57), .ZN(n55) );
  AOI21_X1 U168 ( .B1(n54), .B2(n183), .A(n51), .ZN(n49) );
  NAND2_X1 U169 ( .A1(n164), .A2(n59), .ZN(n8) );
  INV_X1 U170 ( .A(n90), .ZN(n88) );
  OAI21_X1 U171 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  INV_X1 U172 ( .A(n53), .ZN(n51) );
  INV_X1 U173 ( .A(n172), .ZN(n94) );
  NAND2_X1 U174 ( .A1(n99), .A2(n62), .ZN(n9) );
  INV_X1 U175 ( .A(n61), .ZN(n99) );
  NAND2_X1 U176 ( .A1(n183), .A2(n53), .ZN(n7) );
  NAND2_X1 U177 ( .A1(n104), .A2(n82), .ZN(n14) );
  INV_X1 U178 ( .A(n81), .ZN(n104) );
  NAND2_X1 U179 ( .A1(n102), .A2(n74), .ZN(n12) );
  INV_X1 U180 ( .A(n73), .ZN(n102) );
  NAND2_X1 U181 ( .A1(n185), .A2(n71), .ZN(n11) );
  NAND2_X1 U182 ( .A1(n186), .A2(n79), .ZN(n13) );
  NAND2_X1 U183 ( .A1(n184), .A2(n87), .ZN(n15) );
  NAND2_X1 U184 ( .A1(n100), .A2(n66), .ZN(n10) );
  INV_X1 U185 ( .A(n65), .ZN(n100) );
  INV_X1 U186 ( .A(n28), .ZN(n30) );
  XOR2_X1 U187 ( .A(n14), .B(n83), .Z(SUM[2]) );
  XNOR2_X1 U188 ( .A(n15), .B(n88), .ZN(SUM[1]) );
  NOR2_X1 U189 ( .A1(A[7]), .A2(B[7]), .ZN(n61) );
  OR2_X1 U190 ( .A1(A[9]), .A2(B[9]), .ZN(n183) );
  NOR2_X1 U191 ( .A1(A[2]), .A2(B[2]), .ZN(n81) );
  NAND2_X1 U192 ( .A1(n94), .A2(n37), .ZN(n4) );
  NAND2_X1 U193 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  OR2_X1 U194 ( .A1(A[1]), .A2(B[1]), .ZN(n184) );
  NOR2_X1 U195 ( .A1(A[6]), .A2(B[6]), .ZN(n65) );
  NOR2_X1 U196 ( .A1(A[11]), .A2(B[11]), .ZN(n39) );
  XNOR2_X1 U197 ( .A(n60), .B(n8), .ZN(SUM[8]) );
  XNOR2_X1 U198 ( .A(n54), .B(n7), .ZN(SUM[9]) );
  NOR2_X1 U199 ( .A1(A[4]), .A2(B[4]), .ZN(n73) );
  NAND2_X1 U200 ( .A1(A[7]), .A2(B[7]), .ZN(n62) );
  OR2_X1 U201 ( .A1(A[5]), .A2(B[5]), .ZN(n185) );
  OR2_X1 U202 ( .A1(A[3]), .A2(B[3]), .ZN(n186) );
  NAND2_X1 U203 ( .A1(A[2]), .A2(B[2]), .ZN(n82) );
  NAND2_X1 U204 ( .A1(A[15]), .A2(B[15]), .ZN(n18) );
  NAND2_X1 U205 ( .A1(A[9]), .A2(B[9]), .ZN(n53) );
  NAND2_X1 U206 ( .A1(A[5]), .A2(B[5]), .ZN(n71) );
  NAND2_X1 U207 ( .A1(A[3]), .A2(B[3]), .ZN(n79) );
  NAND2_X1 U208 ( .A1(A[1]), .A2(B[1]), .ZN(n87) );
  NAND2_X1 U209 ( .A1(A[0]), .A2(B[0]), .ZN(n90) );
  NAND2_X1 U210 ( .A1(A[6]), .A2(B[6]), .ZN(n66) );
  NAND2_X1 U211 ( .A1(A[4]), .A2(B[4]), .ZN(n74) );
  NAND2_X1 U212 ( .A1(A[12]), .A2(B[12]), .ZN(n37) );
  XOR2_X1 U213 ( .A(n63), .B(n9), .Z(SUM[7]) );
  XNOR2_X1 U214 ( .A(n11), .B(n72), .ZN(SUM[5]) );
  XOR2_X1 U215 ( .A(n12), .B(n75), .Z(SUM[4]) );
  XNOR2_X1 U216 ( .A(n13), .B(n80), .ZN(SUM[3]) );
  INV_X1 U217 ( .A(n189), .ZN(n48) );
  NOR2_X1 U218 ( .A1(n167), .A2(n61), .ZN(n56) );
  OAI21_X1 U219 ( .B1(n58), .B2(n62), .A(n59), .ZN(n57) );
  NAND2_X1 U220 ( .A1(A[8]), .A2(B[8]), .ZN(n59) );
  XOR2_X1 U221 ( .A(n10), .B(n67), .Z(SUM[6]) );
  AND2_X1 U222 ( .A1(A[10]), .A2(B[10]), .ZN(n189) );
  OAI21_X1 U223 ( .B1(n75), .B2(n73), .A(n74), .ZN(n72) );
  NAND2_X1 U224 ( .A1(A[11]), .A2(B[11]), .ZN(n40) );
  NAND2_X1 U225 ( .A1(n166), .A2(n18), .ZN(n1) );
  NOR2_X1 U226 ( .A1(A[13]), .A2(B[13]), .ZN(n27) );
  OAI21_X1 U227 ( .B1(n41), .B2(n39), .A(n163), .ZN(n38) );
  NAND2_X1 U228 ( .A1(n162), .A2(n25), .ZN(n2) );
  NAND2_X1 U229 ( .A1(n161), .A2(n171), .ZN(n20) );
  NAND2_X1 U230 ( .A1(A[14]), .A2(B[14]), .ZN(n25) );
  INV_X1 U231 ( .A(n42), .ZN(n41) );
  NOR2_X1 U232 ( .A1(n36), .A2(n39), .ZN(n34) );
  OAI21_X1 U233 ( .B1(n36), .B2(n40), .A(n37), .ZN(n35) );
  XNOR2_X1 U234 ( .A(n19), .B(n1), .ZN(SUM[15]) );
  OAI21_X1 U235 ( .B1(n43), .B2(n173), .A(n44), .ZN(n42) );
  NAND2_X1 U236 ( .A1(n188), .A2(n183), .ZN(n43) );
  AOI21_X1 U237 ( .B1(n188), .B2(n51), .A(n189), .ZN(n44) );
  XNOR2_X1 U238 ( .A(n38), .B(n4), .ZN(SUM[12]) );
  XNOR2_X1 U239 ( .A(n26), .B(n2), .ZN(SUM[14]) );
  OAI21_X1 U240 ( .B1(n33), .B2(n27), .A(n28), .ZN(n26) );
  OAI21_X1 U241 ( .B1(n181), .B2(n20), .A(n21), .ZN(n19) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_9 ( clk, clear_acc, 
        data_out_x, data_out, data_out_w, data_out_b, wr_en_y, m_valid, 
        m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [3:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N27, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, n1, n2, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n87, n104, n113, n114, n115, n116, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n18), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n219), .CK(clk), .Q(n22) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n220), .CK(clk), .Q(n23) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n221), .CK(clk), .Q(n24) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n222), .CK(clk), .Q(n25) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n223), .CK(clk), .Q(n26) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n224), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n225), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n226), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n227), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n228), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n229), .CK(clk), .Q(n34) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n230), .CK(clk), .Q(n35) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n231), .CK(clk), .Q(n36) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n232), .CK(clk), .Q(n37) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n233), .CK(clk), .Q(n38) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n234), .CK(clk), .Q(n39) );
  DFF_X1 \f_reg[7]  ( .D(n80), .CK(clk), .Q(f[7]), .QN(n211) );
  DFF_X1 \f_reg[8]  ( .D(n79), .CK(clk), .Q(f[8]), .QN(n212) );
  DFF_X1 \f_reg[9]  ( .D(n78), .CK(clk), .Q(f[9]), .QN(n213) );
  DFF_X1 \f_reg[10]  ( .D(n77), .CK(clk), .Q(n49), .QN(n214) );
  DFF_X1 \f_reg[11]  ( .D(n76), .CK(clk), .Q(n47), .QN(n215) );
  DFF_X1 \f_reg[12]  ( .D(n2), .CK(clk), .Q(n46), .QN(n216) );
  DFF_X1 \f_reg[13]  ( .D(n75), .CK(clk), .Q(n44), .QN(n217) );
  DFF_X1 \f_reg[14]  ( .D(n8), .CK(clk), .Q(n43), .QN(n218) );
  DFF_X1 \f_reg[15]  ( .D(n7), .CK(clk), .Q(f[15]), .QN(n73) );
  DFF_X1 \data_out_reg[15]  ( .D(n113), .CK(clk), .Q(data_out[15]), .QN(n191)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n114), .CK(clk), .Q(data_out[14]), .QN(n190)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n115), .CK(clk), .Q(data_out[13]), .QN(n189)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n116), .CK(clk), .Q(data_out[12]), .QN(n188)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n164), .CK(clk), .Q(data_out[11]), .QN(n187)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n165), .CK(clk), .Q(data_out[10]), .QN(n186)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n166), .CK(clk), .Q(data_out[9]), .QN(n185) );
  DFF_X1 \data_out_reg[8]  ( .D(n167), .CK(clk), .Q(data_out[8]), .QN(n184) );
  DFF_X1 \data_out_reg[7]  ( .D(n168), .CK(clk), .Q(data_out[7]), .QN(n183) );
  DFF_X1 \data_out_reg[6]  ( .D(n169), .CK(clk), .Q(data_out[6]), .QN(n182) );
  DFF_X1 \data_out_reg[5]  ( .D(n170), .CK(clk), .Q(data_out[5]), .QN(n181) );
  DFF_X1 \data_out_reg[4]  ( .D(n171), .CK(clk), .Q(data_out[4]), .QN(n180) );
  DFF_X1 \data_out_reg[3]  ( .D(n172), .CK(clk), .Q(data_out[3]), .QN(n179) );
  DFF_X1 \data_out_reg[2]  ( .D(n173), .CK(clk), .Q(data_out[2]), .QN(n178) );
  DFF_X1 \data_out_reg[1]  ( .D(n174), .CK(clk), .Q(data_out[1]), .QN(n177) );
  DFF_X1 \data_out_reg[0]  ( .D(n175), .CK(clk), .Q(data_out[0]), .QN(n176) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_9_DW_mult_tc_1 mult_960 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_9_DW01_add_2 add_961 ( .A({n198, 
        n197, n196, n195, n194, n193, n207, n206, n205, n204, n203, n202, n201, 
        n200, n199, n192}), .B({f[15], n43, n44, n46, n47, n49, f[9:3], n57, 
        n59, n61}), .CI(1'b0), .SUM(adder) );
  DFF_X2 delay_reg ( .D(N27), .CK(clk), .Q(n12), .QN(n235) );
  DFF_X1 \f_reg[3]  ( .D(n84), .CK(clk), .Q(f[3]), .QN(n65) );
  DFF_X1 \f_reg[0]  ( .D(n104), .CK(clk), .Q(n61), .QN(n208) );
  DFF_X1 \f_reg[2]  ( .D(n85), .CK(clk), .Q(n57), .QN(n210) );
  DFF_X1 \f_reg[1]  ( .D(n87), .CK(clk), .Q(n59), .QN(n209) );
  DFF_X1 \f_reg[4]  ( .D(n83), .CK(clk), .Q(f[4]), .QN(n66) );
  DFF_X1 \f_reg[5]  ( .D(n82), .CK(clk), .Q(f[5]), .QN(n67) );
  DFF_X1 \f_reg[6]  ( .D(n81), .CK(clk), .Q(f[6]), .QN(n68) );
  AND2_X1 U3 ( .A1(clear_acc_delay), .A2(n235), .ZN(n1) );
  AND2_X2 U4 ( .A1(n42), .A2(n19), .ZN(n16) );
  NAND3_X1 U5 ( .A1(n5), .A2(n4), .A3(n6), .ZN(n2) );
  MUX2_X2 U6 ( .A(n29), .B(N37), .S(n235), .Z(n206) );
  MUX2_X2 U8 ( .A(n24), .B(N42), .S(n235), .Z(n196) );
  NAND2_X1 U9 ( .A1(data_out_b[12]), .A2(n18), .ZN(n4) );
  NAND2_X1 U10 ( .A1(adder[12]), .A2(n16), .ZN(n5) );
  NAND2_X1 U11 ( .A1(n63), .A2(n46), .ZN(n6) );
  NAND3_X1 U12 ( .A1(n10), .A2(n9), .A3(n11), .ZN(n7) );
  MUX2_X2 U13 ( .A(N43), .B(n23), .S(n12), .Z(n197) );
  MUX2_X2 U14 ( .A(n26), .B(N40), .S(n235), .Z(n194) );
  MUX2_X2 U15 ( .A(n25), .B(N41), .S(n235), .Z(n195) );
  NAND3_X1 U16 ( .A1(n14), .A2(n13), .A3(n15), .ZN(n8) );
  NAND2_X1 U17 ( .A1(data_out_b[15]), .A2(n18), .ZN(n9) );
  NAND2_X1 U18 ( .A1(adder[15]), .A2(n16), .ZN(n10) );
  NAND2_X1 U19 ( .A1(n63), .A2(f[15]), .ZN(n11) );
  NAND2_X1 U20 ( .A1(data_out_b[14]), .A2(n18), .ZN(n13) );
  NAND2_X1 U21 ( .A1(adder[14]), .A2(n16), .ZN(n14) );
  NAND2_X1 U22 ( .A1(n63), .A2(n43), .ZN(n15) );
  INV_X2 U23 ( .A(n42), .ZN(n63) );
  INV_X1 U24 ( .A(n19), .ZN(n18) );
  INV_X1 U25 ( .A(clear_acc), .ZN(n19) );
  NAND2_X1 U26 ( .A1(n17), .A2(N27), .ZN(n237) );
  OAI22_X1 U27 ( .A1(n179), .A2(n237), .B1(n65), .B2(n236), .ZN(n172) );
  OAI22_X1 U28 ( .A1(n180), .A2(n237), .B1(n66), .B2(n236), .ZN(n171) );
  OAI22_X1 U29 ( .A1(n181), .A2(n237), .B1(n67), .B2(n236), .ZN(n170) );
  OAI22_X1 U30 ( .A1(n182), .A2(n237), .B1(n68), .B2(n236), .ZN(n169) );
  OAI22_X1 U31 ( .A1(n183), .A2(n237), .B1(n211), .B2(n236), .ZN(n168) );
  OAI22_X1 U32 ( .A1(n184), .A2(n237), .B1(n212), .B2(n236), .ZN(n167) );
  OAI22_X1 U33 ( .A1(n185), .A2(n237), .B1(n213), .B2(n236), .ZN(n166) );
  INV_X1 U34 ( .A(wr_en_y), .ZN(n17) );
  AND2_X1 U35 ( .A1(sel[0]), .A2(sel[1]), .ZN(n21) );
  INV_X1 U36 ( .A(m_ready), .ZN(n20) );
  NAND2_X1 U37 ( .A1(m_valid), .A2(n20), .ZN(n40) );
  OAI211_X1 U38 ( .C1(sel[2]), .C2(n21), .A(sel[3]), .B(n40), .ZN(N27) );
  MUX2_X1 U39 ( .A(n22), .B(N44), .S(n1), .Z(n219) );
  MUX2_X1 U40 ( .A(n22), .B(N44), .S(n235), .Z(n198) );
  MUX2_X1 U41 ( .A(n23), .B(N43), .S(n1), .Z(n220) );
  MUX2_X1 U42 ( .A(n24), .B(N42), .S(n1), .Z(n221) );
  MUX2_X1 U43 ( .A(n25), .B(N41), .S(n1), .Z(n222) );
  MUX2_X1 U44 ( .A(n26), .B(N40), .S(n1), .Z(n223) );
  MUX2_X1 U45 ( .A(n27), .B(N39), .S(n1), .Z(n224) );
  MUX2_X1 U46 ( .A(n27), .B(N39), .S(n235), .Z(n193) );
  MUX2_X1 U47 ( .A(n28), .B(N38), .S(n1), .Z(n225) );
  MUX2_X1 U48 ( .A(n28), .B(N38), .S(n235), .Z(n207) );
  MUX2_X1 U49 ( .A(n29), .B(N37), .S(n1), .Z(n226) );
  MUX2_X1 U50 ( .A(n32), .B(N36), .S(n1), .Z(n227) );
  MUX2_X1 U51 ( .A(n32), .B(N36), .S(n235), .Z(n205) );
  MUX2_X1 U52 ( .A(n33), .B(N35), .S(n1), .Z(n228) );
  MUX2_X1 U53 ( .A(n33), .B(N35), .S(n235), .Z(n204) );
  MUX2_X1 U54 ( .A(n34), .B(N34), .S(n1), .Z(n229) );
  MUX2_X1 U55 ( .A(n34), .B(N34), .S(n235), .Z(n203) );
  MUX2_X1 U56 ( .A(n35), .B(N33), .S(n1), .Z(n230) );
  MUX2_X1 U57 ( .A(n35), .B(N33), .S(n235), .Z(n202) );
  MUX2_X1 U58 ( .A(n36), .B(N32), .S(n1), .Z(n231) );
  MUX2_X1 U59 ( .A(n36), .B(N32), .S(n235), .Z(n201) );
  MUX2_X1 U60 ( .A(n37), .B(N31), .S(n1), .Z(n232) );
  MUX2_X1 U61 ( .A(n37), .B(N31), .S(n235), .Z(n200) );
  MUX2_X1 U62 ( .A(n38), .B(N30), .S(n1), .Z(n233) );
  MUX2_X1 U63 ( .A(n38), .B(N30), .S(n235), .Z(n199) );
  MUX2_X1 U64 ( .A(n39), .B(N29), .S(n1), .Z(n234) );
  MUX2_X1 U65 ( .A(n39), .B(N29), .S(n235), .Z(n192) );
  INV_X1 U66 ( .A(n40), .ZN(n41) );
  OAI21_X1 U67 ( .B1(n41), .B2(n12), .A(n19), .ZN(n42) );
  AOI222_X1 U68 ( .A1(data_out_b[13]), .A2(n18), .B1(adder[13]), .B2(n16), 
        .C1(n63), .C2(n44), .ZN(n45) );
  INV_X1 U69 ( .A(n45), .ZN(n75) );
  AOI222_X1 U70 ( .A1(data_out_b[11]), .A2(n18), .B1(adder[11]), .B2(n16), 
        .C1(n63), .C2(n47), .ZN(n48) );
  INV_X1 U71 ( .A(n48), .ZN(n76) );
  AOI222_X1 U72 ( .A1(data_out_b[10]), .A2(n18), .B1(adder[10]), .B2(n16), 
        .C1(n63), .C2(n49), .ZN(n50) );
  INV_X1 U73 ( .A(n50), .ZN(n77) );
  AOI222_X1 U74 ( .A1(data_out_b[8]), .A2(n18), .B1(adder[8]), .B2(n16), .C1(
        n63), .C2(f[8]), .ZN(n51) );
  INV_X1 U75 ( .A(n51), .ZN(n79) );
  AOI222_X1 U76 ( .A1(data_out_b[7]), .A2(n18), .B1(adder[7]), .B2(n16), .C1(
        n63), .C2(f[7]), .ZN(n52) );
  INV_X1 U77 ( .A(n52), .ZN(n80) );
  AOI222_X1 U78 ( .A1(data_out_b[6]), .A2(n18), .B1(adder[6]), .B2(n16), .C1(
        n63), .C2(f[6]), .ZN(n53) );
  INV_X1 U79 ( .A(n53), .ZN(n81) );
  AOI222_X1 U80 ( .A1(data_out_b[5]), .A2(n18), .B1(adder[5]), .B2(n16), .C1(
        n63), .C2(f[5]), .ZN(n54) );
  INV_X1 U81 ( .A(n54), .ZN(n82) );
  AOI222_X1 U82 ( .A1(data_out_b[4]), .A2(n18), .B1(adder[4]), .B2(n16), .C1(
        n63), .C2(f[4]), .ZN(n55) );
  INV_X1 U83 ( .A(n55), .ZN(n83) );
  AOI222_X1 U84 ( .A1(data_out_b[3]), .A2(n18), .B1(adder[3]), .B2(n16), .C1(
        n63), .C2(f[3]), .ZN(n56) );
  INV_X1 U85 ( .A(n56), .ZN(n84) );
  AOI222_X1 U86 ( .A1(data_out_b[2]), .A2(n18), .B1(adder[2]), .B2(n16), .C1(
        n63), .C2(n57), .ZN(n58) );
  INV_X1 U87 ( .A(n58), .ZN(n85) );
  AOI222_X1 U88 ( .A1(data_out_b[1]), .A2(n18), .B1(adder[1]), .B2(n16), .C1(
        n63), .C2(n59), .ZN(n60) );
  INV_X1 U89 ( .A(n60), .ZN(n87) );
  AOI222_X1 U90 ( .A1(data_out_b[0]), .A2(n18), .B1(adder[0]), .B2(n16), .C1(
        n63), .C2(n61), .ZN(n62) );
  INV_X1 U91 ( .A(n62), .ZN(n104) );
  AOI222_X1 U92 ( .A1(data_out_b[9]), .A2(n18), .B1(adder[9]), .B2(n16), .C1(
        n63), .C2(f[9]), .ZN(n64) );
  INV_X1 U93 ( .A(n64), .ZN(n78) );
  NOR4_X1 U94 ( .A1(n47), .A2(n46), .A3(n44), .A4(n43), .ZN(n72) );
  NOR4_X1 U95 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n49), .ZN(n71) );
  NAND4_X1 U96 ( .A1(n68), .A2(n67), .A3(n66), .A4(n65), .ZN(n69) );
  NOR4_X1 U97 ( .A1(n69), .A2(n61), .A3(n59), .A4(n57), .ZN(n70) );
  NAND3_X1 U98 ( .A1(n72), .A2(n71), .A3(n70), .ZN(n74) );
  NAND3_X1 U99 ( .A1(wr_en_y), .A2(n74), .A3(n73), .ZN(n236) );
  OAI22_X1 U100 ( .A1(n176), .A2(n237), .B1(n208), .B2(n236), .ZN(n175) );
  OAI22_X1 U101 ( .A1(n177), .A2(n237), .B1(n209), .B2(n236), .ZN(n174) );
  OAI22_X1 U102 ( .A1(n178), .A2(n237), .B1(n210), .B2(n236), .ZN(n173) );
  OAI22_X1 U103 ( .A1(n186), .A2(n237), .B1(n214), .B2(n236), .ZN(n165) );
  OAI22_X1 U104 ( .A1(n187), .A2(n237), .B1(n215), .B2(n236), .ZN(n164) );
  OAI22_X1 U105 ( .A1(n188), .A2(n237), .B1(n216), .B2(n236), .ZN(n116) );
  OAI22_X1 U106 ( .A1(n189), .A2(n237), .B1(n217), .B2(n236), .ZN(n115) );
  OAI22_X1 U107 ( .A1(n190), .A2(n237), .B1(n218), .B2(n236), .ZN(n114) );
  OAI22_X1 U108 ( .A1(n191), .A2(n237), .B1(n73), .B2(n236), .ZN(n113) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_8_DW_mult_tc_1 ( a, b, 
        product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n9, n13, n16, n18, n19, n21, n23, n25, n29, n31, n32, n34,
         n36, n37, n39, n40, n41, n42, n43, n46, n47, n48, n50, n53, n54, n55,
         n56, n57, n58, n59, n62, n63, n64, n65, n67, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n93, n95, n96, n97, n98, n99, n103, n104, n105,
         n106, n107, n109, n111, n112, n113, n114, n115, n117, n119, n120,
         n122, n125, n126, n129, n131, n135, n139, n141, n142, n143, n144,
         n145, n146, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n237, n245, n247, n249, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n418, n419, n420, n421, n422, n423, n424, n426, n427, n428, n429,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U148 ( .A(n265), .B(n144), .Z(n145) );
  XOR2_X1 U152 ( .A(n301), .B(n148), .Z(n149) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U161 ( .A(n177), .B(n168), .CI(n166), .CO(n163), .S(n164) );
  FA_X1 U162 ( .A(n172), .B(n170), .CI(n179), .CO(n165), .S(n166) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n291), .CI(n263), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n252), .B(n317), .CO(n173), .S(n174) );
  FA_X1 U167 ( .A(n180), .B(n187), .CI(n178), .CO(n175), .S(n176) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U169 ( .A(n193), .B(n282), .CI(n191), .CO(n179), .S(n180) );
  FA_X1 U170 ( .A(n274), .B(n268), .CI(n292), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U172 ( .A(n197), .B(n190), .CI(n188), .CO(n185), .S(n186) );
  FA_X1 U173 ( .A(n199), .B(n201), .CI(n192), .CO(n187), .S(n188) );
  FA_X1 U174 ( .A(n194), .B(n275), .CI(n293), .CO(n189), .S(n190) );
  FA_X1 U175 ( .A(n283), .B(n253), .CI(n305), .CO(n191), .S(n192) );
  HA_X1 U176 ( .A(n269), .B(n319), .CO(n193), .S(n194) );
  FA_X1 U177 ( .A(n205), .B(n200), .CI(n198), .CO(n195), .S(n196) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U179 ( .A(n276), .B(n284), .CI(n294), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n320), .B(n270), .CI(n306), .CO(n201), .S(n202) );
  FA_X1 U182 ( .A(n215), .B(n307), .CI(n210), .CO(n205), .S(n206) );
  FA_X1 U183 ( .A(n254), .B(n285), .CI(n295), .CO(n207), .S(n208) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U187 ( .A(n322), .B(n278), .CI(n308), .CO(n215), .S(n216) );
  FA_X1 U188 ( .A(n225), .B(n222), .CI(n220), .CO(n217), .S(n218) );
  FA_X1 U189 ( .A(n255), .B(n309), .CI(n297), .CO(n219), .S(n220) );
  HA_X1 U190 ( .A(n287), .B(n323), .CO(n221), .S(n222) );
  FA_X1 U191 ( .A(n229), .B(n298), .CI(n226), .CO(n223), .S(n224) );
  FA_X1 U192 ( .A(n288), .B(n324), .CI(n310), .CO(n225), .S(n226) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  HA_X1 U194 ( .A(n311), .B(n325), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n326), .B(n312), .CI(n300), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  AND2_X1 U414 ( .A1(n558), .A2(n557), .ZN(n490) );
  AND2_X1 U415 ( .A1(n558), .A2(n557), .ZN(n555) );
  XNOR2_X1 U416 ( .A(n583), .B(a[6]), .ZN(n491) );
  CLKBUF_X1 U417 ( .A(n91), .Z(n549) );
  BUF_X1 U418 ( .A(n16), .Z(n535) );
  NAND2_X1 U419 ( .A1(n561), .A2(n535), .ZN(n503) );
  OR2_X1 U420 ( .A1(n224), .A2(n227), .ZN(n566) );
  OR2_X1 U421 ( .A1(n329), .A2(n258), .ZN(n492) );
  XNOR2_X1 U422 ( .A(n549), .B(n493), .ZN(product[9]) );
  AND2_X1 U423 ( .A1(n129), .A2(n90), .ZN(n493) );
  OR2_X1 U424 ( .A1(n228), .A2(n231), .ZN(n494) );
  BUF_X2 U425 ( .A(n1), .Z(n527) );
  INV_X1 U426 ( .A(n541), .ZN(n495) );
  INV_X1 U427 ( .A(n541), .ZN(n530) );
  XNOR2_X1 U428 ( .A(n497), .B(n496), .ZN(product[12]) );
  NAND2_X1 U429 ( .A1(n557), .A2(n558), .ZN(n496) );
  NAND2_X1 U430 ( .A1(n126), .A2(n79), .ZN(n497) );
  INV_X1 U431 ( .A(n510), .ZN(n498) );
  INV_X2 U432 ( .A(n585), .ZN(n510) );
  INV_X2 U433 ( .A(n585), .ZN(n584) );
  XNOR2_X1 U434 ( .A(n149), .B(n499), .ZN(n144) );
  XNOR2_X1 U435 ( .A(n271), .B(n146), .ZN(n499) );
  BUF_X2 U436 ( .A(n16), .Z(n571) );
  INV_X1 U437 ( .A(n583), .ZN(n581) );
  AOI21_X1 U438 ( .B1(n567), .B2(n112), .A(n109), .ZN(n500) );
  INV_X2 U439 ( .A(n591), .ZN(n590) );
  NAND2_X1 U440 ( .A1(n561), .A2(n535), .ZN(n18) );
  CLKBUF_X1 U441 ( .A(n548), .Z(n501) );
  INV_X1 U442 ( .A(n573), .ZN(n502) );
  OR2_X1 U443 ( .A1(n196), .A2(n203), .ZN(n504) );
  NAND2_X1 U444 ( .A1(n533), .A2(n429), .ZN(n29) );
  OR2_X1 U445 ( .A1(n538), .A2(n559), .ZN(n531) );
  INV_X1 U446 ( .A(n586), .ZN(n505) );
  BUF_X2 U447 ( .A(n9), .Z(n506) );
  CLKBUF_X1 U448 ( .A(n9), .Z(n572) );
  XNOR2_X1 U449 ( .A(n587), .B(a[8]), .ZN(n429) );
  INV_X1 U450 ( .A(n579), .ZN(n507) );
  INV_X2 U451 ( .A(n580), .ZN(n579) );
  INV_X1 U452 ( .A(n559), .ZN(n508) );
  CLKBUF_X1 U453 ( .A(n546), .Z(n509) );
  INV_X1 U454 ( .A(n548), .ZN(n511) );
  OR2_X1 U455 ( .A1(n186), .A2(n195), .ZN(n512) );
  NOR2_X1 U456 ( .A1(n196), .A2(n203), .ZN(n85) );
  XOR2_X1 U457 ( .A(n286), .B(n296), .Z(n513) );
  XOR2_X1 U458 ( .A(n513), .B(n221), .Z(n214) );
  XOR2_X1 U459 ( .A(n216), .B(n219), .Z(n514) );
  XOR2_X1 U460 ( .A(n514), .B(n214), .Z(n212) );
  NAND2_X1 U461 ( .A1(n286), .A2(n296), .ZN(n515) );
  NAND2_X1 U462 ( .A1(n286), .A2(n221), .ZN(n516) );
  NAND2_X1 U463 ( .A1(n296), .A2(n221), .ZN(n517) );
  NAND3_X1 U464 ( .A1(n515), .A2(n516), .A3(n517), .ZN(n213) );
  NAND2_X1 U465 ( .A1(n216), .A2(n219), .ZN(n518) );
  NAND2_X1 U466 ( .A1(n216), .A2(n214), .ZN(n519) );
  NAND2_X1 U467 ( .A1(n219), .A2(n214), .ZN(n520) );
  NAND3_X1 U468 ( .A1(n518), .A2(n519), .A3(n520), .ZN(n211) );
  CLKBUF_X1 U469 ( .A(n7), .Z(n521) );
  NOR2_X2 U470 ( .A1(n176), .A2(n185), .ZN(n78) );
  CLKBUF_X1 U471 ( .A(n104), .Z(n522) );
  AOI21_X1 U472 ( .B1(n554), .B2(n522), .A(n556), .ZN(n523) );
  XNOR2_X1 U473 ( .A(n88), .B(n524), .ZN(product[10]) );
  NAND2_X1 U474 ( .A1(n504), .A2(n86), .ZN(n524) );
  XNOR2_X1 U475 ( .A(n589), .B(a[10]), .ZN(n428) );
  NOR2_X1 U476 ( .A1(n186), .A2(n195), .ZN(n525) );
  NOR2_X1 U477 ( .A1(n186), .A2(n195), .ZN(n82) );
  INV_X1 U478 ( .A(n587), .ZN(n526) );
  INV_X1 U479 ( .A(n587), .ZN(n586) );
  BUF_X1 U480 ( .A(n37), .Z(n528) );
  XNOR2_X1 U481 ( .A(n583), .B(a[4]), .ZN(n561) );
  XOR2_X1 U482 ( .A(n585), .B(a[6]), .Z(n538) );
  INV_X1 U483 ( .A(n581), .ZN(n529) );
  XNOR2_X1 U484 ( .A(n19), .B(a[8]), .ZN(n533) );
  INV_X1 U485 ( .A(n533), .ZN(n541) );
  NAND2_X1 U486 ( .A1(n32), .A2(n428), .ZN(n532) );
  OAI21_X1 U487 ( .B1(n91), .B2(n89), .A(n90), .ZN(n534) );
  CLKBUF_X1 U488 ( .A(n18), .Z(n536) );
  BUF_X2 U489 ( .A(n577), .Z(n537) );
  INV_X1 U490 ( .A(n577), .ZN(n553) );
  OR2_X2 U491 ( .A1(n538), .A2(n491), .ZN(n23) );
  INV_X1 U492 ( .A(n559), .ZN(n21) );
  INV_X2 U493 ( .A(n589), .ZN(n588) );
  CLKBUF_X1 U494 ( .A(n96), .Z(n539) );
  NOR2_X1 U495 ( .A1(n164), .A2(n175), .ZN(n540) );
  NOR2_X1 U496 ( .A1(n164), .A2(n175), .ZN(n75) );
  INV_X1 U497 ( .A(n548), .ZN(n32) );
  XOR2_X1 U498 ( .A(n208), .B(n213), .Z(n542) );
  XOR2_X1 U499 ( .A(n206), .B(n542), .Z(n204) );
  NAND2_X1 U500 ( .A1(n206), .A2(n208), .ZN(n543) );
  NAND2_X1 U501 ( .A1(n206), .A2(n213), .ZN(n544) );
  NAND2_X1 U502 ( .A1(n208), .A2(n213), .ZN(n545) );
  NAND3_X1 U503 ( .A1(n543), .A2(n544), .A3(n545), .ZN(n203) );
  XNOR2_X1 U504 ( .A(n580), .B(a[2]), .ZN(n560) );
  NAND2_X1 U505 ( .A1(n560), .A2(n9), .ZN(n546) );
  NAND2_X1 U506 ( .A1(n560), .A2(n9), .ZN(n547) );
  XOR2_X1 U507 ( .A(n580), .B(a[4]), .Z(n16) );
  XNOR2_X1 U508 ( .A(n587), .B(a[10]), .ZN(n548) );
  OR2_X1 U509 ( .A1(n550), .A2(n553), .ZN(n6) );
  XNOR2_X1 U510 ( .A(n1), .B(n249), .ZN(n550) );
  OR2_X2 U511 ( .A1(n550), .A2(n553), .ZN(n551) );
  OR2_X2 U512 ( .A1(n550), .A2(n553), .ZN(n552) );
  CLKBUF_X1 U513 ( .A(n566), .Z(n554) );
  AND2_X1 U514 ( .A1(n224), .A2(n227), .ZN(n556) );
  NAND2_X1 U515 ( .A1(n534), .A2(n80), .ZN(n557) );
  INV_X1 U516 ( .A(n81), .ZN(n558) );
  XNOR2_X1 U517 ( .A(n583), .B(a[6]), .ZN(n559) );
  BUF_X1 U518 ( .A(n43), .Z(n575) );
  NAND2_X1 U519 ( .A1(n562), .A2(n69), .ZN(n47) );
  INV_X1 U520 ( .A(n73), .ZN(n71) );
  AOI21_X1 U521 ( .B1(n74), .B2(n562), .A(n67), .ZN(n65) );
  INV_X1 U522 ( .A(n69), .ZN(n67) );
  NAND2_X1 U523 ( .A1(n562), .A2(n73), .ZN(n64) );
  INV_X1 U524 ( .A(n74), .ZN(n72) );
  AOI21_X1 U525 ( .B1(n96), .B2(n563), .A(n93), .ZN(n91) );
  INV_X1 U526 ( .A(n95), .ZN(n93) );
  INV_X1 U527 ( .A(n78), .ZN(n126) );
  OR2_X1 U528 ( .A1(n152), .A2(n163), .ZN(n562) );
  NAND2_X1 U529 ( .A1(n125), .A2(n76), .ZN(n48) );
  INV_X1 U530 ( .A(n75), .ZN(n125) );
  OAI21_X1 U531 ( .B1(n540), .B2(n79), .A(n76), .ZN(n74) );
  INV_X1 U532 ( .A(n89), .ZN(n129) );
  NOR2_X1 U533 ( .A1(n75), .A2(n78), .ZN(n73) );
  XNOR2_X1 U534 ( .A(n84), .B(n50), .ZN(product[11]) );
  NAND2_X1 U535 ( .A1(n512), .A2(n83), .ZN(n50) );
  NAND2_X1 U536 ( .A1(n152), .A2(n163), .ZN(n69) );
  NAND2_X1 U537 ( .A1(n563), .A2(n95), .ZN(n53) );
  INV_X1 U538 ( .A(n111), .ZN(n109) );
  NAND2_X1 U539 ( .A1(n494), .A2(n106), .ZN(n56) );
  NAND2_X1 U540 ( .A1(n131), .A2(n98), .ZN(n54) );
  INV_X1 U541 ( .A(n97), .ZN(n131) );
  OR2_X1 U542 ( .A1(n212), .A2(n217), .ZN(n563) );
  NAND2_X1 U543 ( .A1(n566), .A2(n103), .ZN(n55) );
  AOI21_X1 U544 ( .B1(n564), .B2(n120), .A(n117), .ZN(n115) );
  INV_X1 U545 ( .A(n119), .ZN(n117) );
  XOR2_X1 U546 ( .A(n58), .B(n115), .Z(product[3]) );
  NAND2_X1 U547 ( .A1(n135), .A2(n114), .ZN(n58) );
  XNOR2_X1 U548 ( .A(n57), .B(n112), .ZN(product[4]) );
  NAND2_X1 U549 ( .A1(n567), .A2(n111), .ZN(n57) );
  NAND2_X1 U550 ( .A1(n176), .A2(n185), .ZN(n79) );
  NAND2_X1 U551 ( .A1(n164), .A2(n175), .ZN(n76) );
  NAND2_X1 U552 ( .A1(n212), .A2(n217), .ZN(n95) );
  NAND2_X1 U553 ( .A1(n204), .A2(n211), .ZN(n90) );
  NAND2_X1 U554 ( .A1(n196), .A2(n203), .ZN(n86) );
  XNOR2_X1 U555 ( .A(n59), .B(n120), .ZN(product[2]) );
  NAND2_X1 U556 ( .A1(n564), .A2(n119), .ZN(n59) );
  NAND2_X1 U557 ( .A1(n328), .A2(n314), .ZN(n119) );
  OR2_X1 U558 ( .A1(n328), .A2(n314), .ZN(n564) );
  OR2_X1 U559 ( .A1(n151), .A2(n139), .ZN(n565) );
  NOR2_X1 U560 ( .A1(n228), .A2(n231), .ZN(n105) );
  NOR2_X1 U561 ( .A1(n218), .A2(n223), .ZN(n97) );
  NOR2_X1 U562 ( .A1(n234), .A2(n257), .ZN(n113) );
  NAND2_X1 U563 ( .A1(n218), .A2(n223), .ZN(n98) );
  NAND2_X1 U564 ( .A1(n228), .A2(n231), .ZN(n106) );
  INV_X1 U565 ( .A(n37), .ZN(n237) );
  OR2_X1 U566 ( .A1(n232), .A2(n233), .ZN(n567) );
  INV_X1 U567 ( .A(n41), .ZN(n235) );
  AND2_X1 U568 ( .A1(n492), .A2(n122), .ZN(product[1]) );
  XNOR2_X1 U569 ( .A(n588), .B(a[12]), .ZN(n37) );
  OR2_X1 U570 ( .A1(n575), .A2(n507), .ZN(n392) );
  XNOR2_X1 U571 ( .A(n521), .B(n575), .ZN(n391) );
  XNOR2_X1 U572 ( .A(n590), .B(a[14]), .ZN(n41) );
  INV_X1 U573 ( .A(n249), .ZN(n577) );
  AND2_X1 U574 ( .A1(n576), .A2(n237), .ZN(n264) );
  XNOR2_X1 U575 ( .A(n526), .B(n575), .ZN(n352) );
  AND2_X1 U576 ( .A1(n576), .A2(n501), .ZN(n270) );
  AND2_X1 U577 ( .A1(n576), .A2(n491), .ZN(n288) );
  OAI22_X1 U578 ( .A1(n39), .A2(n336), .B1(n528), .B2(n335), .ZN(n263) );
  XNOR2_X1 U579 ( .A(n582), .B(n575), .ZN(n376) );
  XNOR2_X1 U580 ( .A(n155), .B(n569), .ZN(n139) );
  XNOR2_X1 U581 ( .A(n153), .B(n141), .ZN(n569) );
  XNOR2_X1 U582 ( .A(n157), .B(n570), .ZN(n141) );
  XNOR2_X1 U583 ( .A(n145), .B(n143), .ZN(n570) );
  OAI22_X1 U584 ( .A1(n39), .A2(n591), .B1(n337), .B2(n528), .ZN(n252) );
  OR2_X1 U585 ( .A1(n575), .A2(n591), .ZN(n337) );
  OAI22_X1 U586 ( .A1(n42), .A2(n593), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U587 ( .A1(n575), .A2(n593), .ZN(n332) );
  AND2_X1 U588 ( .A1(n576), .A2(n245), .ZN(n300) );
  XOR2_X1 U589 ( .A(n315), .B(n261), .Z(n150) );
  OAI22_X1 U590 ( .A1(n39), .A2(n334), .B1(n528), .B2(n333), .ZN(n261) );
  XNOR2_X1 U591 ( .A(n590), .B(n575), .ZN(n336) );
  AND2_X1 U592 ( .A1(n576), .A2(n247), .ZN(n314) );
  AND2_X1 U593 ( .A1(n576), .A2(n235), .ZN(n260) );
  OAI22_X1 U594 ( .A1(n39), .A2(n335), .B1(n528), .B2(n334), .ZN(n262) );
  NAND2_X1 U595 ( .A1(n427), .A2(n37), .ZN(n39) );
  XOR2_X1 U596 ( .A(n590), .B(a[12]), .Z(n427) );
  INV_X1 U597 ( .A(n25), .ZN(n587) );
  AND2_X1 U598 ( .A1(n576), .A2(n541), .ZN(n278) );
  NAND2_X1 U599 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U600 ( .A(n592), .B(a[14]), .Z(n426) );
  INV_X1 U601 ( .A(n13), .ZN(n583) );
  XNOR2_X1 U602 ( .A(n510), .B(n575), .ZN(n363) );
  AND2_X1 U603 ( .A1(n576), .A2(n249), .ZN(product[0]) );
  OR2_X1 U604 ( .A1(n575), .A2(n589), .ZN(n344) );
  OR2_X1 U605 ( .A1(n575), .A2(n498), .ZN(n364) );
  OR2_X1 U606 ( .A1(n575), .A2(n529), .ZN(n377) );
  OR2_X1 U607 ( .A1(n575), .A2(n505), .ZN(n353) );
  XNOR2_X1 U608 ( .A(n578), .B(b[15]), .ZN(n393) );
  XNOR2_X1 U609 ( .A(n510), .B(b[9]), .ZN(n354) );
  XNOR2_X1 U610 ( .A(n582), .B(b[11]), .ZN(n365) );
  XNOR2_X1 U611 ( .A(n590), .B(n424), .ZN(n335) );
  XNOR2_X1 U612 ( .A(n590), .B(n423), .ZN(n334) );
  OAI22_X1 U613 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U614 ( .A(n592), .B(n424), .ZN(n330) );
  XNOR2_X1 U615 ( .A(n592), .B(n575), .ZN(n331) );
  XNOR2_X1 U616 ( .A(n526), .B(n418), .ZN(n345) );
  XNOR2_X1 U617 ( .A(n588), .B(n420), .ZN(n338) );
  XNOR2_X1 U618 ( .A(n579), .B(b[13]), .ZN(n378) );
  XNOR2_X1 U619 ( .A(n521), .B(n424), .ZN(n390) );
  XNOR2_X1 U620 ( .A(n586), .B(n424), .ZN(n351) );
  XNOR2_X1 U621 ( .A(n584), .B(n424), .ZN(n362) );
  XNOR2_X1 U622 ( .A(n579), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U623 ( .A(n579), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U624 ( .A(n579), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U625 ( .A(n579), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U626 ( .A(n579), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U627 ( .A(n579), .B(n419), .ZN(n385) );
  XNOR2_X1 U628 ( .A(n579), .B(n418), .ZN(n384) );
  XNOR2_X1 U629 ( .A(n582), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U630 ( .A(n582), .B(n418), .ZN(n369) );
  XNOR2_X1 U631 ( .A(n582), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U632 ( .A(n582), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U633 ( .A(n521), .B(n422), .ZN(n388) );
  XNOR2_X1 U634 ( .A(n521), .B(n423), .ZN(n389) );
  XNOR2_X1 U635 ( .A(n526), .B(n422), .ZN(n349) );
  XNOR2_X1 U636 ( .A(n586), .B(n423), .ZN(n350) );
  XNOR2_X1 U637 ( .A(n584), .B(n422), .ZN(n360) );
  XNOR2_X1 U638 ( .A(n584), .B(n423), .ZN(n361) );
  XNOR2_X1 U639 ( .A(n578), .B(b[11]), .ZN(n397) );
  XNOR2_X1 U640 ( .A(n578), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U641 ( .A(n578), .B(b[13]), .ZN(n395) );
  XNOR2_X1 U642 ( .A(n578), .B(b[14]), .ZN(n394) );
  XNOR2_X1 U643 ( .A(n590), .B(n422), .ZN(n333) );
  XNOR2_X1 U644 ( .A(n584), .B(n421), .ZN(n359) );
  XNOR2_X1 U645 ( .A(n584), .B(n420), .ZN(n358) );
  XNOR2_X1 U646 ( .A(n521), .B(n421), .ZN(n387) );
  XNOR2_X1 U647 ( .A(n586), .B(n421), .ZN(n348) );
  XNOR2_X1 U648 ( .A(n526), .B(n420), .ZN(n347) );
  XNOR2_X1 U649 ( .A(n521), .B(n420), .ZN(n386) );
  XNOR2_X1 U650 ( .A(n588), .B(n421), .ZN(n339) );
  XNOR2_X1 U651 ( .A(n510), .B(n418), .ZN(n356) );
  XNOR2_X1 U652 ( .A(n510), .B(n419), .ZN(n357) );
  XNOR2_X1 U653 ( .A(n526), .B(n419), .ZN(n346) );
  XNOR2_X1 U654 ( .A(n510), .B(b[8]), .ZN(n355) );
  BUF_X1 U655 ( .A(n43), .Z(n576) );
  XNOR2_X1 U656 ( .A(n588), .B(n424), .ZN(n342) );
  XNOR2_X1 U657 ( .A(n588), .B(n423), .ZN(n341) );
  XNOR2_X1 U658 ( .A(n588), .B(n575), .ZN(n343) );
  XNOR2_X1 U659 ( .A(n588), .B(n422), .ZN(n340) );
  OAI22_X1 U660 ( .A1(n551), .A2(n395), .B1(n394), .B2(n537), .ZN(n316) );
  OAI22_X1 U661 ( .A1(n552), .A2(n394), .B1(n393), .B2(n537), .ZN(n315) );
  OAI22_X1 U662 ( .A1(n552), .A2(n399), .B1(n398), .B2(n537), .ZN(n320) );
  OAI22_X1 U663 ( .A1(n551), .A2(n401), .B1(n400), .B2(n537), .ZN(n322) );
  OAI22_X1 U664 ( .A1(n551), .A2(n402), .B1(n401), .B2(n537), .ZN(n323) );
  OAI22_X1 U665 ( .A1(n551), .A2(n400), .B1(n399), .B2(n537), .ZN(n321) );
  OAI22_X1 U666 ( .A1(n6), .A2(n404), .B1(n403), .B2(n537), .ZN(n325) );
  OAI22_X1 U667 ( .A1(n552), .A2(n406), .B1(n405), .B2(n537), .ZN(n327) );
  OAI22_X1 U668 ( .A1(n552), .A2(n397), .B1(n396), .B2(n537), .ZN(n318) );
  OAI22_X1 U669 ( .A1(n552), .A2(n405), .B1(n404), .B2(n537), .ZN(n326) );
  OAI22_X1 U670 ( .A1(n552), .A2(n398), .B1(n397), .B2(n537), .ZN(n319) );
  OAI22_X1 U671 ( .A1(n551), .A2(n396), .B1(n395), .B2(n537), .ZN(n317) );
  OAI22_X1 U672 ( .A1(n6), .A2(n403), .B1(n402), .B2(n537), .ZN(n324) );
  OAI22_X1 U673 ( .A1(n552), .A2(n407), .B1(n406), .B2(n537), .ZN(n328) );
  OAI22_X1 U674 ( .A1(n551), .A2(n408), .B1(n407), .B2(n537), .ZN(n329) );
  OAI22_X1 U675 ( .A1(n34), .A2(n339), .B1(n338), .B2(n511), .ZN(n265) );
  OAI22_X1 U676 ( .A1(n532), .A2(n340), .B1(n339), .B2(n511), .ZN(n266) );
  OAI22_X1 U677 ( .A1(n532), .A2(n341), .B1(n340), .B2(n511), .ZN(n267) );
  OAI22_X1 U678 ( .A1(n532), .A2(n342), .B1(n341), .B2(n511), .ZN(n268) );
  OAI22_X1 U679 ( .A1(n532), .A2(n343), .B1(n342), .B2(n511), .ZN(n269) );
  OAI22_X1 U680 ( .A1(n34), .A2(n589), .B1(n344), .B2(n511), .ZN(n253) );
  NAND2_X1 U681 ( .A1(n428), .A2(n32), .ZN(n34) );
  XNOR2_X1 U682 ( .A(a[2]), .B(n1), .ZN(n9) );
  INV_X1 U683 ( .A(n1), .ZN(n573) );
  INV_X1 U684 ( .A(n578), .ZN(n574) );
  INV_X1 U685 ( .A(n19), .ZN(n585) );
  NOR2_X1 U686 ( .A1(n204), .A2(n211), .ZN(n89) );
  OAI22_X1 U687 ( .A1(n29), .A2(n346), .B1(n345), .B2(n495), .ZN(n271) );
  OAI22_X1 U688 ( .A1(n29), .A2(n350), .B1(n349), .B2(n495), .ZN(n275) );
  OAI22_X1 U689 ( .A1(n29), .A2(n347), .B1(n346), .B2(n530), .ZN(n272) );
  OAI22_X1 U690 ( .A1(n29), .A2(n351), .B1(n350), .B2(n530), .ZN(n276) );
  OAI22_X1 U691 ( .A1(n29), .A2(n505), .B1(n353), .B2(n530), .ZN(n254) );
  OAI22_X1 U692 ( .A1(n29), .A2(n348), .B1(n347), .B2(n495), .ZN(n273) );
  OAI22_X1 U693 ( .A1(n29), .A2(n349), .B1(n348), .B2(n495), .ZN(n274) );
  OAI22_X1 U694 ( .A1(n29), .A2(n352), .B1(n351), .B2(n495), .ZN(n277) );
  NOR2_X1 U695 ( .A1(n525), .A2(n85), .ZN(n80) );
  OAI21_X1 U696 ( .B1(n82), .B2(n86), .A(n83), .ZN(n81) );
  NAND2_X1 U697 ( .A1(n186), .A2(n195), .ZN(n83) );
  XNOR2_X1 U698 ( .A(n63), .B(n46), .ZN(product[15]) );
  NAND2_X1 U699 ( .A1(n565), .A2(n62), .ZN(n46) );
  INV_X1 U700 ( .A(n7), .ZN(n580) );
  OAI21_X1 U701 ( .B1(n87), .B2(n85), .A(n86), .ZN(n84) );
  XNOR2_X1 U702 ( .A(n55), .B(n522), .ZN(product[6]) );
  XOR2_X1 U703 ( .A(n56), .B(n500), .Z(product[5]) );
  INV_X1 U704 ( .A(n573), .ZN(n578) );
  OR2_X1 U705 ( .A1(n575), .A2(n574), .ZN(n409) );
  NAND2_X1 U706 ( .A1(n224), .A2(n227), .ZN(n103) );
  OAI21_X1 U707 ( .B1(n91), .B2(n89), .A(n90), .ZN(n88) );
  INV_X1 U708 ( .A(n88), .ZN(n87) );
  OAI21_X1 U709 ( .B1(n113), .B2(n115), .A(n114), .ZN(n112) );
  INV_X1 U710 ( .A(n113), .ZN(n135) );
  XNOR2_X1 U711 ( .A(n77), .B(n48), .ZN(product[13]) );
  OAI22_X1 U712 ( .A1(n23), .A2(n358), .B1(n357), .B2(n21), .ZN(n282) );
  OAI22_X1 U713 ( .A1(n531), .A2(n356), .B1(n355), .B2(n508), .ZN(n280) );
  OAI22_X1 U714 ( .A1(n531), .A2(n362), .B1(n361), .B2(n508), .ZN(n286) );
  OAI22_X1 U715 ( .A1(n23), .A2(n357), .B1(n356), .B2(n508), .ZN(n281) );
  OAI22_X1 U716 ( .A1(n23), .A2(n360), .B1(n359), .B2(n508), .ZN(n284) );
  OAI22_X1 U717 ( .A1(n531), .A2(n498), .B1(n364), .B2(n508), .ZN(n255) );
  OAI22_X1 U718 ( .A1(n23), .A2(n361), .B1(n360), .B2(n21), .ZN(n285) );
  OAI22_X1 U719 ( .A1(n531), .A2(n355), .B1(n354), .B2(n21), .ZN(n279) );
  XNOR2_X1 U720 ( .A(n581), .B(n424), .ZN(n375) );
  OAI22_X1 U721 ( .A1(n531), .A2(n363), .B1(n362), .B2(n21), .ZN(n287) );
  OAI22_X1 U722 ( .A1(n23), .A2(n359), .B1(n358), .B2(n21), .ZN(n283) );
  XNOR2_X1 U723 ( .A(n581), .B(n423), .ZN(n374) );
  XNOR2_X1 U724 ( .A(n581), .B(n421), .ZN(n372) );
  XNOR2_X1 U725 ( .A(n581), .B(n422), .ZN(n373) );
  XNOR2_X1 U726 ( .A(n581), .B(n419), .ZN(n370) );
  XNOR2_X1 U727 ( .A(n581), .B(n420), .ZN(n371) );
  OAI21_X1 U728 ( .B1(n107), .B2(n105), .A(n106), .ZN(n104) );
  AOI21_X1 U729 ( .B1(n567), .B2(n112), .A(n109), .ZN(n107) );
  NAND2_X1 U730 ( .A1(n232), .A2(n233), .ZN(n111) );
  NAND2_X1 U731 ( .A1(n151), .A2(n139), .ZN(n62) );
  OAI22_X1 U732 ( .A1(n536), .A2(n367), .B1(n366), .B2(n571), .ZN(n290) );
  OAI22_X1 U733 ( .A1(n536), .A2(n370), .B1(n369), .B2(n571), .ZN(n293) );
  OAI22_X1 U734 ( .A1(n503), .A2(n368), .B1(n367), .B2(n571), .ZN(n291) );
  OAI22_X1 U735 ( .A1(n18), .A2(n372), .B1(n371), .B2(n571), .ZN(n295) );
  OAI22_X1 U736 ( .A1(n536), .A2(n375), .B1(n374), .B2(n571), .ZN(n298) );
  OAI22_X1 U737 ( .A1(n18), .A2(n369), .B1(n368), .B2(n571), .ZN(n292) );
  OAI22_X1 U738 ( .A1(n503), .A2(n376), .B1(n375), .B2(n571), .ZN(n299) );
  OAI22_X1 U739 ( .A1(n503), .A2(n529), .B1(n377), .B2(n571), .ZN(n256) );
  OAI22_X1 U740 ( .A1(n503), .A2(n371), .B1(n370), .B2(n571), .ZN(n294) );
  OAI22_X1 U741 ( .A1(n18), .A2(n374), .B1(n373), .B2(n571), .ZN(n297) );
  OAI22_X1 U742 ( .A1(n503), .A2(n373), .B1(n372), .B2(n571), .ZN(n296) );
  OAI22_X1 U743 ( .A1(n503), .A2(n366), .B1(n365), .B2(n571), .ZN(n289) );
  INV_X1 U744 ( .A(n535), .ZN(n245) );
  XNOR2_X1 U745 ( .A(n527), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U746 ( .A(n527), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U747 ( .A(n527), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U748 ( .A(n502), .B(n418), .ZN(n401) );
  XNOR2_X1 U749 ( .A(n527), .B(n419), .ZN(n402) );
  XNOR2_X1 U750 ( .A(n527), .B(n420), .ZN(n403) );
  XNOR2_X1 U751 ( .A(n502), .B(n575), .ZN(n408) );
  XNOR2_X1 U752 ( .A(n527), .B(n422), .ZN(n405) );
  XNOR2_X1 U753 ( .A(n527), .B(n421), .ZN(n404) );
  XNOR2_X1 U754 ( .A(n502), .B(n423), .ZN(n406) );
  XNOR2_X1 U755 ( .A(n502), .B(n424), .ZN(n407) );
  OAI21_X1 U756 ( .B1(n490), .B2(n71), .A(n72), .ZN(n70) );
  OAI21_X1 U757 ( .B1(n555), .B2(n78), .A(n79), .ZN(n77) );
  XNOR2_X1 U758 ( .A(n70), .B(n47), .ZN(product[14]) );
  OAI21_X1 U759 ( .B1(n64), .B2(n490), .A(n65), .ZN(n63) );
  XNOR2_X1 U760 ( .A(n539), .B(n53), .ZN(product[8]) );
  INV_X1 U761 ( .A(n122), .ZN(n120) );
  NAND2_X1 U762 ( .A1(n329), .A2(n258), .ZN(n122) );
  OAI21_X1 U763 ( .B1(n99), .B2(n97), .A(n98), .ZN(n96) );
  AOI21_X1 U764 ( .B1(n566), .B2(n104), .A(n556), .ZN(n99) );
  OAI22_X1 U765 ( .A1(n551), .A2(n574), .B1(n409), .B2(n537), .ZN(n258) );
  XOR2_X1 U766 ( .A(n523), .B(n54), .Z(product[7]) );
  OAI22_X1 U767 ( .A1(n509), .A2(n379), .B1(n378), .B2(n506), .ZN(n301) );
  OAI22_X1 U768 ( .A1(n509), .A2(n380), .B1(n379), .B2(n506), .ZN(n302) );
  OAI22_X1 U769 ( .A1(n547), .A2(n385), .B1(n384), .B2(n506), .ZN(n307) );
  OAI22_X1 U770 ( .A1(n547), .A2(n382), .B1(n381), .B2(n506), .ZN(n304) );
  OAI22_X1 U771 ( .A1(n509), .A2(n381), .B1(n380), .B2(n506), .ZN(n303) );
  NAND2_X1 U772 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U773 ( .A1(n383), .A2(n546), .B1(n382), .B2(n506), .ZN(n305) );
  OAI22_X1 U774 ( .A1(n547), .A2(n384), .B1(n383), .B2(n572), .ZN(n306) );
  OAI22_X1 U775 ( .A1(n546), .A2(n386), .B1(n506), .B2(n385), .ZN(n308) );
  OAI22_X1 U776 ( .A1(n547), .A2(n387), .B1(n386), .B2(n506), .ZN(n309) );
  OAI22_X1 U777 ( .A1(n547), .A2(n507), .B1(n392), .B2(n506), .ZN(n257) );
  OAI22_X1 U778 ( .A1(n546), .A2(n389), .B1(n388), .B2(n572), .ZN(n311) );
  OAI22_X1 U779 ( .A1(n546), .A2(n388), .B1(n572), .B2(n387), .ZN(n310) );
  OAI22_X1 U780 ( .A1(n546), .A2(n390), .B1(n389), .B2(n506), .ZN(n312) );
  INV_X1 U781 ( .A(n506), .ZN(n247) );
  OAI22_X1 U782 ( .A1(n547), .A2(n391), .B1(n390), .B2(n506), .ZN(n313) );
  INV_X1 U783 ( .A(n583), .ZN(n582) );
  INV_X1 U784 ( .A(n31), .ZN(n589) );
  INV_X1 U785 ( .A(n36), .ZN(n591) );
  INV_X1 U786 ( .A(n593), .ZN(n592) );
  INV_X1 U787 ( .A(n40), .ZN(n593) );
  XOR2_X1 U788 ( .A(n259), .B(n251), .Z(n148) );
  XOR2_X1 U789 ( .A(n289), .B(n279), .Z(n146) );
  XOR2_X1 U790 ( .A(n159), .B(n150), .Z(n142) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_8_DW01_add_2 ( A, B, CI, SUM, 
        CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n18,
         n19, n20, n21, n25, n26, n28, n30, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n48, n49, n51, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n71, n72, n73, n74,
         n75, n77, n79, n80, n81, n82, n83, n85, n87, n88, n90, n94, n98, n99,
         n100, n102, n104, n161, n162, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177;

  NAND2_X1 U126 ( .A1(A[11]), .A2(B[11]), .ZN(n161) );
  OR2_X1 U127 ( .A1(A[11]), .A2(B[11]), .ZN(n162) );
  AND2_X1 U128 ( .A1(n167), .A2(n90), .ZN(SUM[0]) );
  OR2_X1 U129 ( .A1(A[15]), .A2(B[15]), .ZN(n164) );
  NOR2_X2 U130 ( .A1(A[8]), .A2(B[8]), .ZN(n58) );
  NOR2_X1 U131 ( .A1(A[11]), .A2(B[11]), .ZN(n39) );
  OR2_X2 U132 ( .A1(A[14]), .A2(B[14]), .ZN(n177) );
  AOI21_X1 U133 ( .B1(n42), .B2(n34), .A(n35), .ZN(n165) );
  AOI21_X1 U134 ( .B1(n42), .B2(n34), .A(n35), .ZN(n33) );
  AND2_X1 U135 ( .A1(A[14]), .A2(B[14]), .ZN(n166) );
  OR2_X2 U136 ( .A1(A[10]), .A2(B[10]), .ZN(n173) );
  OR2_X1 U137 ( .A1(A[0]), .A2(B[0]), .ZN(n167) );
  INV_X1 U138 ( .A(n64), .ZN(n63) );
  INV_X1 U139 ( .A(n55), .ZN(n54) );
  INV_X1 U140 ( .A(n71), .ZN(n69) );
  AOI21_X1 U141 ( .B1(n169), .B2(n88), .A(n85), .ZN(n83) );
  INV_X1 U142 ( .A(n87), .ZN(n85) );
  OAI21_X1 U143 ( .B1(n83), .B2(n81), .A(n82), .ZN(n80) );
  NAND2_X1 U144 ( .A1(n177), .A2(n171), .ZN(n20) );
  AOI21_X1 U145 ( .B1(n177), .B2(n30), .A(n166), .ZN(n21) );
  AOI21_X1 U146 ( .B1(n56), .B2(n64), .A(n57), .ZN(n55) );
  AOI21_X1 U147 ( .B1(n170), .B2(n80), .A(n77), .ZN(n75) );
  INV_X1 U148 ( .A(n79), .ZN(n77) );
  AOI21_X1 U149 ( .B1(n54), .B2(n168), .A(n51), .ZN(n49) );
  INV_X1 U150 ( .A(n90), .ZN(n88) );
  OAI21_X1 U151 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  INV_X1 U152 ( .A(n53), .ZN(n51) );
  INV_X1 U153 ( .A(n174), .ZN(n94) );
  NAND2_X1 U154 ( .A1(n170), .A2(n79), .ZN(n13) );
  NAND2_X1 U155 ( .A1(n99), .A2(n62), .ZN(n9) );
  INV_X1 U156 ( .A(n61), .ZN(n99) );
  NAND2_X1 U157 ( .A1(n168), .A2(n53), .ZN(n7) );
  NAND2_X1 U158 ( .A1(n104), .A2(n82), .ZN(n14) );
  INV_X1 U159 ( .A(n81), .ZN(n104) );
  NAND2_X1 U160 ( .A1(n98), .A2(n59), .ZN(n8) );
  INV_X1 U161 ( .A(n58), .ZN(n98) );
  NAND2_X1 U162 ( .A1(n169), .A2(n87), .ZN(n15) );
  NAND2_X1 U163 ( .A1(n172), .A2(n71), .ZN(n11) );
  NAND2_X1 U164 ( .A1(n100), .A2(n66), .ZN(n10) );
  INV_X1 U165 ( .A(n65), .ZN(n100) );
  NAND2_X1 U166 ( .A1(n102), .A2(n74), .ZN(n12) );
  INV_X1 U167 ( .A(n73), .ZN(n102) );
  INV_X1 U168 ( .A(n175), .ZN(n48) );
  XNOR2_X1 U169 ( .A(n13), .B(n80), .ZN(SUM[3]) );
  NAND2_X1 U170 ( .A1(n37), .A2(n94), .ZN(n4) );
  XOR2_X1 U171 ( .A(n41), .B(n5), .Z(SUM[11]) );
  NOR2_X1 U172 ( .A1(A[7]), .A2(B[7]), .ZN(n61) );
  OR2_X1 U173 ( .A1(A[9]), .A2(B[9]), .ZN(n168) );
  NOR2_X1 U174 ( .A1(A[2]), .A2(B[2]), .ZN(n81) );
  XOR2_X1 U175 ( .A(n49), .B(n6), .Z(SUM[10]) );
  OR2_X1 U176 ( .A1(A[1]), .A2(B[1]), .ZN(n169) );
  OR2_X1 U177 ( .A1(A[3]), .A2(B[3]), .ZN(n170) );
  OR2_X1 U178 ( .A1(A[13]), .A2(B[13]), .ZN(n171) );
  XNOR2_X1 U179 ( .A(n60), .B(n8), .ZN(SUM[8]) );
  XNOR2_X1 U180 ( .A(n54), .B(n7), .ZN(SUM[9]) );
  NOR2_X1 U181 ( .A1(A[6]), .A2(B[6]), .ZN(n65) );
  NOR2_X1 U182 ( .A1(A[4]), .A2(B[4]), .ZN(n73) );
  NAND2_X1 U183 ( .A1(A[7]), .A2(B[7]), .ZN(n62) );
  NAND2_X1 U184 ( .A1(A[2]), .A2(B[2]), .ZN(n82) );
  NAND2_X1 U185 ( .A1(A[9]), .A2(B[9]), .ZN(n53) );
  NAND2_X1 U186 ( .A1(A[5]), .A2(B[5]), .ZN(n71) );
  NAND2_X1 U187 ( .A1(A[1]), .A2(B[1]), .ZN(n87) );
  NAND2_X1 U188 ( .A1(A[0]), .A2(B[0]), .ZN(n90) );
  OR2_X1 U189 ( .A1(A[5]), .A2(B[5]), .ZN(n172) );
  NAND2_X1 U190 ( .A1(A[6]), .A2(B[6]), .ZN(n66) );
  NAND2_X1 U191 ( .A1(A[4]), .A2(B[4]), .ZN(n74) );
  NAND2_X1 U192 ( .A1(A[8]), .A2(B[8]), .ZN(n59) );
  XOR2_X1 U193 ( .A(n63), .B(n9), .Z(SUM[7]) );
  XOR2_X1 U194 ( .A(n14), .B(n83), .Z(SUM[2]) );
  XNOR2_X1 U195 ( .A(n15), .B(n88), .ZN(SUM[1]) );
  NAND2_X1 U196 ( .A1(n164), .A2(n18), .ZN(n1) );
  NAND2_X1 U197 ( .A1(A[15]), .A2(B[15]), .ZN(n18) );
  NOR2_X1 U198 ( .A1(A[12]), .A2(B[12]), .ZN(n174) );
  NOR2_X1 U199 ( .A1(A[12]), .A2(B[12]), .ZN(n36) );
  AND2_X1 U200 ( .A1(A[10]), .A2(B[10]), .ZN(n175) );
  NOR2_X1 U201 ( .A1(n58), .A2(n61), .ZN(n56) );
  OAI21_X1 U202 ( .B1(n58), .B2(n62), .A(n59), .ZN(n57) );
  NAND2_X1 U203 ( .A1(n171), .A2(n28), .ZN(n3) );
  INV_X1 U204 ( .A(n28), .ZN(n30) );
  NAND2_X1 U205 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  INV_X1 U206 ( .A(n171), .ZN(n176) );
  NAND2_X1 U207 ( .A1(n177), .A2(n25), .ZN(n2) );
  XOR2_X1 U208 ( .A(n10), .B(n67), .Z(SUM[6]) );
  OAI21_X1 U209 ( .B1(n67), .B2(n65), .A(n66), .ZN(n64) );
  AOI21_X1 U210 ( .B1(n172), .B2(n72), .A(n69), .ZN(n67) );
  XNOR2_X1 U211 ( .A(n11), .B(n72), .ZN(SUM[5]) );
  OAI21_X1 U212 ( .B1(n75), .B2(n73), .A(n74), .ZN(n72) );
  NAND2_X1 U213 ( .A1(A[12]), .A2(B[12]), .ZN(n37) );
  OAI21_X1 U214 ( .B1(n40), .B2(n36), .A(n37), .ZN(n35) );
  NAND2_X1 U215 ( .A1(n162), .A2(n161), .ZN(n5) );
  NAND2_X1 U216 ( .A1(A[11]), .A2(B[11]), .ZN(n40) );
  NAND2_X1 U217 ( .A1(A[14]), .A2(B[14]), .ZN(n25) );
  XOR2_X1 U218 ( .A(n12), .B(n75), .Z(SUM[4]) );
  INV_X1 U219 ( .A(n42), .ZN(n41) );
  NAND2_X1 U220 ( .A1(A[3]), .A2(B[3]), .ZN(n79) );
  OAI21_X1 U221 ( .B1(n41), .B2(n39), .A(n40), .ZN(n38) );
  NOR2_X1 U222 ( .A1(n174), .A2(n39), .ZN(n34) );
  OAI21_X1 U223 ( .B1(n43), .B2(n55), .A(n44), .ZN(n42) );
  AOI21_X1 U224 ( .B1(n173), .B2(n51), .A(n175), .ZN(n44) );
  XNOR2_X1 U225 ( .A(n38), .B(n4), .ZN(SUM[12]) );
  XNOR2_X1 U226 ( .A(n19), .B(n1), .ZN(SUM[15]) );
  NAND2_X1 U227 ( .A1(n173), .A2(n48), .ZN(n6) );
  NAND2_X1 U228 ( .A1(n173), .A2(n168), .ZN(n43) );
  XNOR2_X1 U229 ( .A(n26), .B(n2), .ZN(SUM[14]) );
  XOR2_X1 U230 ( .A(n165), .B(n3), .Z(SUM[13]) );
  OAI21_X1 U231 ( .B1(n33), .B2(n176), .A(n28), .ZN(n26) );
  OAI21_X1 U232 ( .B1(n165), .B2(n20), .A(n21), .ZN(n19) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_8 ( clk, clear_acc, 
        data_out_x, data_out, data_out_w, data_out_b, wr_en_y, m_valid, 
        m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [3:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N27, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, n1, n2, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n87, n104, n113, n114, n115, n116, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n17), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n221), .CK(clk), .Q(n21) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n222), .CK(clk), .Q(n22) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n223), .CK(clk), .Q(n23) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n224), .CK(clk), .Q(n24) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n225), .CK(clk), .Q(n25) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n226), .CK(clk), .Q(n26) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n227), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n228), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n229), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n230), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n231), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n232), .CK(clk), .Q(n34) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n233), .CK(clk), .Q(n35) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n234), .CK(clk), .Q(n36) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n235), .CK(clk), .Q(n37) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n236), .CK(clk), .Q(n38) );
  DFF_X1 \f_reg[8]  ( .D(n80), .CK(clk), .Q(f[8]), .QN(n214) );
  DFF_X1 \f_reg[9]  ( .D(n79), .CK(clk), .Q(f[9]), .QN(n215) );
  DFF_X1 \f_reg[10]  ( .D(n78), .CK(clk), .Q(n49), .QN(n216) );
  DFF_X1 \f_reg[11]  ( .D(n77), .CK(clk), .Q(n47), .QN(n217) );
  DFF_X1 \f_reg[12]  ( .D(n76), .CK(clk), .Q(n45), .QN(n218) );
  DFF_X1 \f_reg[13]  ( .D(n75), .CK(clk), .Q(n43), .QN(n219) );
  DFF_X1 \f_reg[14]  ( .D(n2), .CK(clk), .Q(n42), .QN(n220) );
  DFF_X1 \f_reg[15]  ( .D(n4), .CK(clk), .Q(f[15]), .QN(n73) );
  DFF_X1 \data_out_reg[15]  ( .D(n114), .CK(clk), .Q(data_out[15]), .QN(n193)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n115), .CK(clk), .Q(data_out[14]), .QN(n192)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n116), .CK(clk), .Q(data_out[13]), .QN(n191)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n165), .CK(clk), .Q(data_out[12]), .QN(n190)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n166), .CK(clk), .Q(data_out[11]), .QN(n189)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n167), .CK(clk), .Q(data_out[10]), .QN(n188)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n168), .CK(clk), .Q(data_out[9]), .QN(n187) );
  DFF_X1 \data_out_reg[8]  ( .D(n169), .CK(clk), .Q(data_out[8]), .QN(n186) );
  DFF_X1 \data_out_reg[7]  ( .D(n170), .CK(clk), .Q(data_out[7]), .QN(n185) );
  DFF_X1 \data_out_reg[6]  ( .D(n171), .CK(clk), .Q(data_out[6]), .QN(n184) );
  DFF_X1 \data_out_reg[5]  ( .D(n172), .CK(clk), .Q(data_out[5]), .QN(n183) );
  DFF_X1 \data_out_reg[4]  ( .D(n173), .CK(clk), .Q(data_out[4]), .QN(n182) );
  DFF_X1 \data_out_reg[3]  ( .D(n174), .CK(clk), .Q(data_out[3]), .QN(n181) );
  DFF_X1 \data_out_reg[2]  ( .D(n175), .CK(clk), .Q(data_out[2]), .QN(n180) );
  DFF_X1 \data_out_reg[1]  ( .D(n176), .CK(clk), .Q(data_out[1]), .QN(n179) );
  DFF_X1 \data_out_reg[0]  ( .D(n177), .CK(clk), .Q(data_out[0]), .QN(n178) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_8_DW_mult_tc_1 mult_960 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_8_DW01_add_2 add_961 ( .A({n200, 
        n199, n198, n197, n196, n195, n209, n208, n207, n206, n205, n204, n203, 
        n202, n201, n194}), .B({f[15], n42, n43, n45, n47, n49, f[9:3], n57, 
        n59, n61}), .CI(1'b0), .SUM(adder) );
  DFF_X2 delay_reg ( .D(N27), .CK(clk), .Q(n10), .QN(n237) );
  DFF_X1 \f_reg[2]  ( .D(n87), .CK(clk), .Q(n57), .QN(n212) );
  DFF_X1 \f_reg[1]  ( .D(n104), .CK(clk), .Q(n59), .QN(n211) );
  DFF_X1 \f_reg[4]  ( .D(n84), .CK(clk), .Q(f[4]), .QN(n66) );
  DFF_X1 \f_reg[3]  ( .D(n85), .CK(clk), .Q(f[3]), .QN(n65) );
  DFF_X1 \f_reg[0]  ( .D(n113), .CK(clk), .Q(n61), .QN(n210) );
  DFF_X1 \f_reg[5]  ( .D(n83), .CK(clk), .Q(f[5]), .QN(n67) );
  DFF_X1 \f_reg[6]  ( .D(n82), .CK(clk), .Q(f[6]), .QN(n68) );
  DFF_X1 \f_reg[7]  ( .D(n81), .CK(clk), .Q(f[7]), .QN(n213) );
  MUX2_X1 U3 ( .A(N39), .B(n26), .S(n10), .Z(n195) );
  AND2_X1 U4 ( .A1(clear_acc_delay), .A2(n237), .ZN(n1) );
  AND2_X2 U5 ( .A1(n41), .A2(n18), .ZN(n14) );
  MUX2_X2 U6 ( .A(n28), .B(N37), .S(n237), .Z(n208) );
  NAND3_X1 U8 ( .A1(n8), .A2(n7), .A3(n9), .ZN(n2) );
  MUX2_X2 U9 ( .A(n25), .B(N40), .S(n237), .Z(n196) );
  NAND3_X1 U10 ( .A1(n12), .A2(n11), .A3(n13), .ZN(n4) );
  NAND2_X1 U11 ( .A1(N41), .A2(n237), .ZN(n5) );
  NAND2_X1 U12 ( .A1(n24), .A2(n10), .ZN(n6) );
  NAND2_X1 U13 ( .A1(n5), .A2(n6), .ZN(n197) );
  NAND2_X1 U14 ( .A1(data_out_b[14]), .A2(n17), .ZN(n7) );
  NAND2_X1 U15 ( .A1(adder[14]), .A2(n14), .ZN(n8) );
  NAND2_X1 U16 ( .A1(n63), .A2(n42), .ZN(n9) );
  NAND2_X1 U17 ( .A1(data_out_b[15]), .A2(n17), .ZN(n11) );
  NAND2_X1 U18 ( .A1(adder[15]), .A2(n14), .ZN(n12) );
  NAND2_X1 U19 ( .A1(n63), .A2(f[15]), .ZN(n13) );
  INV_X2 U20 ( .A(n41), .ZN(n63) );
  INV_X1 U21 ( .A(n18), .ZN(n17) );
  INV_X1 U22 ( .A(clear_acc), .ZN(n18) );
  NAND2_X1 U23 ( .A1(n16), .A2(N27), .ZN(n239) );
  OAI22_X1 U24 ( .A1(n181), .A2(n239), .B1(n65), .B2(n238), .ZN(n174) );
  OAI22_X1 U25 ( .A1(n182), .A2(n239), .B1(n66), .B2(n238), .ZN(n173) );
  OAI22_X1 U26 ( .A1(n183), .A2(n239), .B1(n67), .B2(n238), .ZN(n172) );
  OAI22_X1 U27 ( .A1(n184), .A2(n239), .B1(n68), .B2(n238), .ZN(n171) );
  OAI22_X1 U28 ( .A1(n185), .A2(n239), .B1(n213), .B2(n238), .ZN(n170) );
  OAI22_X1 U29 ( .A1(n186), .A2(n239), .B1(n214), .B2(n238), .ZN(n169) );
  OAI22_X1 U30 ( .A1(n187), .A2(n239), .B1(n215), .B2(n238), .ZN(n168) );
  MUX2_X1 U31 ( .A(n23), .B(N42), .S(n237), .Z(n198) );
  CLKBUF_X1 U32 ( .A(N39), .Z(n15) );
  INV_X1 U33 ( .A(wr_en_y), .ZN(n16) );
  AND2_X1 U34 ( .A1(sel[0]), .A2(sel[1]), .ZN(n20) );
  INV_X1 U35 ( .A(m_ready), .ZN(n19) );
  NAND2_X1 U36 ( .A1(m_valid), .A2(n19), .ZN(n39) );
  OAI211_X1 U37 ( .C1(sel[2]), .C2(n20), .A(sel[3]), .B(n39), .ZN(N27) );
  MUX2_X1 U38 ( .A(n21), .B(N44), .S(n1), .Z(n221) );
  MUX2_X1 U39 ( .A(n21), .B(N44), .S(n237), .Z(n200) );
  MUX2_X1 U40 ( .A(n22), .B(N43), .S(n1), .Z(n222) );
  MUX2_X1 U41 ( .A(n22), .B(N43), .S(n237), .Z(n199) );
  MUX2_X1 U42 ( .A(n23), .B(N42), .S(n1), .Z(n223) );
  MUX2_X1 U43 ( .A(n24), .B(N41), .S(n1), .Z(n224) );
  MUX2_X1 U44 ( .A(n25), .B(N40), .S(n1), .Z(n225) );
  MUX2_X1 U45 ( .A(n26), .B(n15), .S(n1), .Z(n226) );
  MUX2_X1 U46 ( .A(n27), .B(N38), .S(n1), .Z(n227) );
  MUX2_X1 U47 ( .A(n27), .B(N38), .S(n237), .Z(n209) );
  MUX2_X1 U48 ( .A(n28), .B(N37), .S(n1), .Z(n228) );
  MUX2_X1 U49 ( .A(n29), .B(N36), .S(n1), .Z(n229) );
  MUX2_X1 U50 ( .A(n29), .B(N36), .S(n237), .Z(n207) );
  MUX2_X1 U51 ( .A(n32), .B(N35), .S(n1), .Z(n230) );
  MUX2_X1 U52 ( .A(n32), .B(N35), .S(n237), .Z(n206) );
  MUX2_X1 U53 ( .A(n33), .B(N34), .S(n1), .Z(n231) );
  MUX2_X1 U54 ( .A(n33), .B(N34), .S(n237), .Z(n205) );
  MUX2_X1 U55 ( .A(n34), .B(N33), .S(n1), .Z(n232) );
  MUX2_X1 U56 ( .A(n34), .B(N33), .S(n237), .Z(n204) );
  MUX2_X1 U57 ( .A(n35), .B(N32), .S(n1), .Z(n233) );
  MUX2_X1 U58 ( .A(n35), .B(N32), .S(n237), .Z(n203) );
  MUX2_X1 U59 ( .A(n36), .B(N31), .S(n1), .Z(n234) );
  MUX2_X1 U60 ( .A(n36), .B(N31), .S(n237), .Z(n202) );
  MUX2_X1 U61 ( .A(n37), .B(N30), .S(n1), .Z(n235) );
  MUX2_X1 U62 ( .A(n37), .B(N30), .S(n237), .Z(n201) );
  MUX2_X1 U63 ( .A(n38), .B(N29), .S(n1), .Z(n236) );
  MUX2_X1 U64 ( .A(n38), .B(N29), .S(n237), .Z(n194) );
  INV_X1 U65 ( .A(n39), .ZN(n40) );
  OAI21_X1 U66 ( .B1(n40), .B2(n10), .A(n18), .ZN(n41) );
  AOI222_X1 U67 ( .A1(data_out_b[13]), .A2(n17), .B1(adder[13]), .B2(n14), 
        .C1(n63), .C2(n43), .ZN(n44) );
  INV_X1 U68 ( .A(n44), .ZN(n75) );
  AOI222_X1 U69 ( .A1(data_out_b[12]), .A2(n17), .B1(adder[12]), .B2(n14), 
        .C1(n63), .C2(n45), .ZN(n46) );
  INV_X1 U70 ( .A(n46), .ZN(n76) );
  AOI222_X1 U71 ( .A1(data_out_b[11]), .A2(n17), .B1(adder[11]), .B2(n14), 
        .C1(n63), .C2(n47), .ZN(n48) );
  INV_X1 U72 ( .A(n48), .ZN(n77) );
  AOI222_X1 U73 ( .A1(data_out_b[10]), .A2(n17), .B1(adder[10]), .B2(n14), 
        .C1(n63), .C2(n49), .ZN(n50) );
  INV_X1 U74 ( .A(n50), .ZN(n78) );
  AOI222_X1 U75 ( .A1(data_out_b[8]), .A2(n17), .B1(adder[8]), .B2(n14), .C1(
        n63), .C2(f[8]), .ZN(n51) );
  INV_X1 U76 ( .A(n51), .ZN(n80) );
  AOI222_X1 U77 ( .A1(data_out_b[7]), .A2(n17), .B1(adder[7]), .B2(n14), .C1(
        n63), .C2(f[7]), .ZN(n52) );
  INV_X1 U78 ( .A(n52), .ZN(n81) );
  AOI222_X1 U79 ( .A1(data_out_b[6]), .A2(n17), .B1(adder[6]), .B2(n14), .C1(
        n63), .C2(f[6]), .ZN(n53) );
  INV_X1 U80 ( .A(n53), .ZN(n82) );
  AOI222_X1 U81 ( .A1(data_out_b[5]), .A2(n17), .B1(adder[5]), .B2(n14), .C1(
        n63), .C2(f[5]), .ZN(n54) );
  INV_X1 U82 ( .A(n54), .ZN(n83) );
  AOI222_X1 U83 ( .A1(data_out_b[4]), .A2(n17), .B1(adder[4]), .B2(n14), .C1(
        n63), .C2(f[4]), .ZN(n55) );
  INV_X1 U84 ( .A(n55), .ZN(n84) );
  AOI222_X1 U85 ( .A1(data_out_b[3]), .A2(n17), .B1(adder[3]), .B2(n14), .C1(
        n63), .C2(f[3]), .ZN(n56) );
  INV_X1 U86 ( .A(n56), .ZN(n85) );
  AOI222_X1 U87 ( .A1(data_out_b[2]), .A2(n17), .B1(adder[2]), .B2(n14), .C1(
        n63), .C2(n57), .ZN(n58) );
  INV_X1 U88 ( .A(n58), .ZN(n87) );
  AOI222_X1 U89 ( .A1(data_out_b[1]), .A2(n17), .B1(adder[1]), .B2(n14), .C1(
        n63), .C2(n59), .ZN(n60) );
  INV_X1 U90 ( .A(n60), .ZN(n104) );
  AOI222_X1 U91 ( .A1(data_out_b[0]), .A2(n17), .B1(adder[0]), .B2(n14), .C1(
        n63), .C2(n61), .ZN(n62) );
  INV_X1 U92 ( .A(n62), .ZN(n113) );
  AOI222_X1 U93 ( .A1(data_out_b[9]), .A2(n17), .B1(adder[9]), .B2(n14), .C1(
        n63), .C2(f[9]), .ZN(n64) );
  INV_X1 U94 ( .A(n64), .ZN(n79) );
  NOR4_X1 U95 ( .A1(n47), .A2(n45), .A3(n43), .A4(n42), .ZN(n72) );
  NOR4_X1 U96 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n49), .ZN(n71) );
  NAND4_X1 U97 ( .A1(n68), .A2(n67), .A3(n66), .A4(n65), .ZN(n69) );
  NOR4_X1 U98 ( .A1(n69), .A2(n61), .A3(n59), .A4(n57), .ZN(n70) );
  NAND3_X1 U99 ( .A1(n72), .A2(n71), .A3(n70), .ZN(n74) );
  NAND3_X1 U100 ( .A1(wr_en_y), .A2(n74), .A3(n73), .ZN(n238) );
  OAI22_X1 U101 ( .A1(n178), .A2(n239), .B1(n210), .B2(n238), .ZN(n177) );
  OAI22_X1 U102 ( .A1(n179), .A2(n239), .B1(n211), .B2(n238), .ZN(n176) );
  OAI22_X1 U103 ( .A1(n180), .A2(n239), .B1(n212), .B2(n238), .ZN(n175) );
  OAI22_X1 U104 ( .A1(n188), .A2(n239), .B1(n216), .B2(n238), .ZN(n167) );
  OAI22_X1 U105 ( .A1(n189), .A2(n239), .B1(n217), .B2(n238), .ZN(n166) );
  OAI22_X1 U106 ( .A1(n190), .A2(n239), .B1(n218), .B2(n238), .ZN(n165) );
  OAI22_X1 U107 ( .A1(n191), .A2(n239), .B1(n219), .B2(n238), .ZN(n116) );
  OAI22_X1 U108 ( .A1(n192), .A2(n239), .B1(n220), .B2(n238), .ZN(n115) );
  OAI22_X1 U109 ( .A1(n193), .A2(n239), .B1(n73), .B2(n238), .ZN(n114) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_7_DW_mult_tc_1 ( a, b, 
        product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n9, n12, n13, n16, n18, n19, n21, n23, n25, n29, n31, n32,
         n34, n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n50, n53,
         n54, n55, n56, n57, n58, n59, n62, n63, n64, n65, n67, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n93, n95, n96, n97, n98, n99, n103,
         n104, n105, n106, n107, n109, n111, n112, n113, n114, n115, n117,
         n119, n120, n122, n126, n127, n128, n131, n135, n139, n141, n142,
         n143, n144, n145, n146, n147, n148, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n249, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n418,
         n419, n420, n421, n422, n423, n424, n426, n427, n428, n429, n430,
         n433, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U148 ( .A(n265), .B(n144), .Z(n145) );
  XOR2_X1 U150 ( .A(n271), .B(n146), .Z(n147) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U161 ( .A(n177), .B(n168), .CI(n166), .CO(n163), .S(n164) );
  FA_X1 U162 ( .A(n170), .B(n172), .CI(n179), .CO(n165), .S(n166) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n291), .CI(n263), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n317), .B(n252), .CO(n173), .S(n174) );
  FA_X1 U167 ( .A(n180), .B(n187), .CI(n178), .CO(n175), .S(n176) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U169 ( .A(n193), .B(n282), .CI(n191), .CO(n179), .S(n180) );
  FA_X1 U170 ( .A(n268), .B(n292), .CI(n274), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U172 ( .A(n197), .B(n190), .CI(n188), .CO(n185), .S(n186) );
  FA_X1 U173 ( .A(n199), .B(n201), .CI(n192), .CO(n187), .S(n188) );
  FA_X1 U174 ( .A(n275), .B(n293), .CI(n194), .CO(n189), .S(n190) );
  FA_X1 U175 ( .A(n283), .B(n305), .CI(n253), .CO(n191), .S(n192) );
  HA_X1 U176 ( .A(n269), .B(n319), .CO(n193), .S(n194) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U179 ( .A(n276), .B(n284), .CI(n294), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n320), .B(n270), .CI(n306), .CO(n201), .S(n202) );
  FA_X1 U181 ( .A(n208), .B(n213), .CI(n206), .CO(n203), .S(n204) );
  FA_X1 U182 ( .A(n210), .B(n307), .CI(n215), .CO(n205), .S(n206) );
  FA_X1 U183 ( .A(n254), .B(n285), .CI(n295), .CO(n207), .S(n208) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U185 ( .A(n216), .B(n219), .CI(n214), .CO(n211), .S(n212) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n322), .B(n278), .CI(n308), .CO(n215), .S(n216) );
  FA_X1 U188 ( .A(n225), .B(n222), .CI(n220), .CO(n217), .S(n218) );
  FA_X1 U189 ( .A(n255), .B(n309), .CI(n297), .CO(n219), .S(n220) );
  HA_X1 U190 ( .A(n287), .B(n323), .CO(n221), .S(n222) );
  FA_X1 U191 ( .A(n229), .B(n298), .CI(n226), .CO(n223), .S(n224) );
  FA_X1 U192 ( .A(n324), .B(n288), .CI(n310), .CO(n225), .S(n226) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  HA_X1 U194 ( .A(n325), .B(n311), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n312), .B(n300), .CI(n326), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  OR2_X2 U414 ( .A1(n524), .A2(n525), .ZN(n12) );
  INV_X1 U415 ( .A(n503), .ZN(n37) );
  OR2_X1 U416 ( .A1(n164), .A2(n175), .ZN(n490) );
  BUF_X1 U417 ( .A(n9), .Z(n519) );
  OR2_X1 U418 ( .A1(n329), .A2(n258), .ZN(n491) );
  INV_X1 U419 ( .A(n25), .ZN(n492) );
  OR2_X1 U420 ( .A1(n228), .A2(n231), .ZN(n493) );
  OR2_X1 U421 ( .A1(n524), .A2(n525), .ZN(n517) );
  OR2_X1 U422 ( .A1(n524), .A2(n525), .ZN(n516) );
  XNOR2_X1 U423 ( .A(n513), .B(n494), .ZN(product[9]) );
  AND2_X1 U424 ( .A1(n511), .A2(n90), .ZN(n494) );
  INV_X1 U425 ( .A(n547), .ZN(n495) );
  INV_X1 U426 ( .A(n547), .ZN(n21) );
  BUF_X1 U427 ( .A(n562), .Z(n521) );
  OR2_X2 U428 ( .A1(n224), .A2(n227), .ZN(n550) );
  XOR2_X1 U429 ( .A(n205), .B(n200), .Z(n496) );
  XOR2_X1 U430 ( .A(n198), .B(n496), .Z(n196) );
  NAND2_X1 U431 ( .A1(n198), .A2(n205), .ZN(n497) );
  NAND2_X1 U432 ( .A1(n198), .A2(n200), .ZN(n498) );
  NAND2_X1 U433 ( .A1(n205), .A2(n200), .ZN(n499) );
  NAND3_X1 U434 ( .A1(n497), .A2(n498), .A3(n499), .ZN(n195) );
  BUF_X1 U435 ( .A(n539), .Z(n500) );
  INV_X1 U436 ( .A(n492), .ZN(n501) );
  INV_X1 U437 ( .A(n492), .ZN(n502) );
  INV_X1 U438 ( .A(n573), .ZN(n572) );
  INV_X1 U439 ( .A(n526), .ZN(n534) );
  XNOR2_X1 U440 ( .A(n575), .B(a[12]), .ZN(n503) );
  NAND2_X1 U441 ( .A1(n430), .A2(n528), .ZN(n504) );
  NAND2_X1 U442 ( .A1(n430), .A2(n528), .ZN(n505) );
  NAND2_X1 U443 ( .A1(n430), .A2(n528), .ZN(n23) );
  CLKBUF_X2 U444 ( .A(n19), .Z(n515) );
  XNOR2_X1 U445 ( .A(n506), .B(n147), .ZN(n144) );
  XNOR2_X1 U446 ( .A(n301), .B(n148), .ZN(n506) );
  OR2_X1 U447 ( .A1(n531), .A2(n540), .ZN(n512) );
  OR2_X1 U448 ( .A1(n531), .A2(n540), .ZN(n18) );
  INV_X1 U449 ( .A(n570), .ZN(n568) );
  INV_X1 U450 ( .A(n538), .ZN(n507) );
  INV_X1 U451 ( .A(n538), .ZN(n32) );
  INV_X2 U452 ( .A(n577), .ZN(n576) );
  XNOR2_X1 U453 ( .A(n522), .B(b[10]), .ZN(n508) );
  BUF_X2 U454 ( .A(n562), .Z(n522) );
  XOR2_X1 U455 ( .A(n572), .B(a[8]), .Z(n509) );
  BUF_X1 U456 ( .A(n96), .Z(n541) );
  XOR2_X1 U457 ( .A(n570), .B(a[4]), .Z(n531) );
  CLKBUF_X1 U458 ( .A(n567), .Z(n510) );
  INV_X1 U459 ( .A(n1), .ZN(n564) );
  OR2_X1 U460 ( .A1(n204), .A2(n211), .ZN(n511) );
  AOI21_X1 U461 ( .B1(n541), .B2(n549), .A(n93), .ZN(n513) );
  AOI21_X1 U462 ( .B1(n96), .B2(n549), .A(n93), .ZN(n91) );
  CLKBUF_X1 U463 ( .A(n224), .Z(n514) );
  XNOR2_X1 U464 ( .A(n575), .B(a[10]), .ZN(n428) );
  INV_X1 U465 ( .A(n563), .ZN(n518) );
  CLKBUF_X1 U466 ( .A(n9), .Z(n557) );
  NAND2_X1 U467 ( .A1(n428), .A2(n32), .ZN(n520) );
  BUF_X2 U468 ( .A(n562), .Z(n523) );
  INV_X1 U469 ( .A(n564), .ZN(n562) );
  XOR2_X1 U470 ( .A(n567), .B(a[2]), .Z(n524) );
  XNOR2_X1 U471 ( .A(n564), .B(a[2]), .ZN(n525) );
  XNOR2_X2 U472 ( .A(n19), .B(a[8]), .ZN(n526) );
  OAI21_X1 U473 ( .B1(n91), .B2(n89), .A(n90), .ZN(n527) );
  XOR2_X1 U474 ( .A(n570), .B(a[6]), .Z(n528) );
  AOI21_X1 U475 ( .B1(n550), .B2(n104), .A(n545), .ZN(n529) );
  BUF_X2 U476 ( .A(n561), .Z(n530) );
  INV_X1 U477 ( .A(n249), .ZN(n561) );
  INV_X1 U478 ( .A(n540), .ZN(n16) );
  INV_X2 U479 ( .A(n575), .ZN(n574) );
  INV_X1 U480 ( .A(n568), .ZN(n532) );
  NOR2_X1 U481 ( .A1(n164), .A2(n175), .ZN(n533) );
  NOR2_X1 U482 ( .A1(n164), .A2(n175), .ZN(n75) );
  OAI21_X1 U483 ( .B1(n91), .B2(n89), .A(n90), .ZN(n88) );
  XNOR2_X1 U484 ( .A(n571), .B(a[6]), .ZN(n430) );
  XNOR2_X1 U485 ( .A(n527), .B(n535), .ZN(product[10]) );
  NAND2_X1 U486 ( .A1(n128), .A2(n86), .ZN(n535) );
  CLKBUF_X1 U487 ( .A(n107), .Z(n536) );
  NOR2_X1 U488 ( .A1(n186), .A2(n195), .ZN(n537) );
  NOR2_X1 U489 ( .A1(n186), .A2(n195), .ZN(n82) );
  INV_X1 U490 ( .A(n567), .ZN(n565) );
  XNOR2_X1 U491 ( .A(n573), .B(a[10]), .ZN(n538) );
  NAND2_X1 U492 ( .A1(n429), .A2(n526), .ZN(n539) );
  NAND2_X1 U493 ( .A1(n509), .A2(n526), .ZN(n29) );
  XNOR2_X1 U494 ( .A(n564), .B(n249), .ZN(n433) );
  XOR2_X1 U495 ( .A(n564), .B(a[2]), .Z(n9) );
  XNOR2_X1 U496 ( .A(n567), .B(a[4]), .ZN(n540) );
  NOR2_X2 U497 ( .A1(n176), .A2(n185), .ZN(n78) );
  CLKBUF_X1 U498 ( .A(n104), .Z(n542) );
  NAND2_X1 U499 ( .A1(n433), .A2(n561), .ZN(n543) );
  NAND2_X1 U500 ( .A1(n433), .A2(n561), .ZN(n544) );
  NAND2_X1 U501 ( .A1(n433), .A2(n561), .ZN(n6) );
  AND2_X1 U502 ( .A1(n224), .A2(n227), .ZN(n545) );
  AOI21_X1 U503 ( .B1(n88), .B2(n80), .A(n81), .ZN(n546) );
  XNOR2_X1 U504 ( .A(n570), .B(a[6]), .ZN(n547) );
  BUF_X1 U505 ( .A(n43), .Z(n559) );
  XNOR2_X1 U506 ( .A(n70), .B(n47), .ZN(product[14]) );
  NAND2_X1 U507 ( .A1(n548), .A2(n69), .ZN(n47) );
  INV_X1 U508 ( .A(n73), .ZN(n71) );
  AOI21_X1 U509 ( .B1(n548), .B2(n74), .A(n67), .ZN(n65) );
  INV_X1 U510 ( .A(n69), .ZN(n67) );
  INV_X1 U511 ( .A(n74), .ZN(n72) );
  INV_X1 U512 ( .A(n95), .ZN(n93) );
  AOI21_X1 U513 ( .B1(n80), .B2(n527), .A(n81), .ZN(n45) );
  NOR2_X1 U514 ( .A1(n537), .A2(n85), .ZN(n80) );
  OAI21_X1 U515 ( .B1(n82), .B2(n86), .A(n83), .ZN(n81) );
  INV_X1 U516 ( .A(n85), .ZN(n128) );
  INV_X1 U517 ( .A(n78), .ZN(n126) );
  OR2_X1 U518 ( .A1(n152), .A2(n163), .ZN(n548) );
  NAND2_X1 U519 ( .A1(n549), .A2(n95), .ZN(n53) );
  NAND2_X1 U520 ( .A1(n490), .A2(n76), .ZN(n48) );
  OAI21_X1 U521 ( .B1(n533), .B2(n79), .A(n76), .ZN(n74) );
  NOR2_X1 U522 ( .A1(n75), .A2(n78), .ZN(n73) );
  XNOR2_X1 U523 ( .A(n84), .B(n50), .ZN(product[11]) );
  NAND2_X1 U524 ( .A1(n127), .A2(n83), .ZN(n50) );
  INV_X1 U525 ( .A(n537), .ZN(n127) );
  NAND2_X1 U526 ( .A1(n152), .A2(n163), .ZN(n69) );
  OAI21_X1 U527 ( .B1(n113), .B2(n115), .A(n114), .ZN(n112) );
  AOI21_X1 U528 ( .B1(n552), .B2(n112), .A(n109), .ZN(n107) );
  NAND2_X1 U529 ( .A1(n493), .A2(n106), .ZN(n56) );
  NAND2_X1 U530 ( .A1(n131), .A2(n98), .ZN(n54) );
  INV_X1 U531 ( .A(n97), .ZN(n131) );
  NOR2_X1 U532 ( .A1(n196), .A2(n203), .ZN(n85) );
  NAND2_X1 U533 ( .A1(n550), .A2(n103), .ZN(n55) );
  OAI21_X1 U534 ( .B1(n105), .B2(n107), .A(n106), .ZN(n104) );
  AOI21_X1 U535 ( .B1(n551), .B2(n120), .A(n117), .ZN(n115) );
  INV_X1 U536 ( .A(n119), .ZN(n117) );
  INV_X1 U537 ( .A(n122), .ZN(n120) );
  XNOR2_X1 U538 ( .A(n63), .B(n46), .ZN(product[15]) );
  NAND2_X1 U539 ( .A1(n553), .A2(n62), .ZN(n46) );
  NAND2_X1 U540 ( .A1(n73), .A2(n548), .ZN(n64) );
  XNOR2_X1 U541 ( .A(n57), .B(n112), .ZN(product[4]) );
  NAND2_X1 U542 ( .A1(n552), .A2(n111), .ZN(n57) );
  XNOR2_X1 U543 ( .A(n59), .B(n120), .ZN(product[2]) );
  NAND2_X1 U544 ( .A1(n551), .A2(n119), .ZN(n59) );
  NAND2_X1 U545 ( .A1(n186), .A2(n195), .ZN(n83) );
  NAND2_X1 U546 ( .A1(n164), .A2(n175), .ZN(n76) );
  NAND2_X1 U547 ( .A1(n176), .A2(n185), .ZN(n79) );
  NAND2_X1 U548 ( .A1(n196), .A2(n203), .ZN(n86) );
  NAND2_X1 U549 ( .A1(n212), .A2(n217), .ZN(n95) );
  INV_X1 U550 ( .A(n113), .ZN(n135) );
  OR2_X1 U551 ( .A1(n212), .A2(n217), .ZN(n549) );
  NAND2_X1 U552 ( .A1(n204), .A2(n211), .ZN(n90) );
  NOR2_X1 U553 ( .A1(n228), .A2(n231), .ZN(n105) );
  OR2_X1 U554 ( .A1(n328), .A2(n314), .ZN(n551) );
  NOR2_X1 U555 ( .A1(n234), .A2(n257), .ZN(n113) );
  NAND2_X1 U556 ( .A1(n328), .A2(n314), .ZN(n119) );
  NOR2_X1 U557 ( .A1(n218), .A2(n223), .ZN(n97) );
  NAND2_X1 U558 ( .A1(n228), .A2(n231), .ZN(n106) );
  OR2_X1 U559 ( .A1(n232), .A2(n233), .ZN(n552) );
  NAND2_X1 U560 ( .A1(n218), .A2(n223), .ZN(n98) );
  NAND2_X1 U561 ( .A1(n514), .A2(n227), .ZN(n103) );
  NAND2_X1 U562 ( .A1(n232), .A2(n233), .ZN(n111) );
  INV_X1 U563 ( .A(n41), .ZN(n235) );
  OR2_X1 U564 ( .A1(n151), .A2(n139), .ZN(n553) );
  AND2_X1 U565 ( .A1(n491), .A2(n122), .ZN(product[1]) );
  OR2_X1 U566 ( .A1(n559), .A2(n510), .ZN(n392) );
  OAI22_X1 U567 ( .A1(n543), .A2(n407), .B1(n406), .B2(n530), .ZN(n328) );
  XNOR2_X1 U568 ( .A(n576), .B(a[14]), .ZN(n41) );
  XNOR2_X1 U569 ( .A(n569), .B(n559), .ZN(n376) );
  OAI22_X1 U570 ( .A1(n543), .A2(n408), .B1(n407), .B2(n530), .ZN(n329) );
  OAI22_X1 U571 ( .A1(n544), .A2(n406), .B1(n405), .B2(n530), .ZN(n327) );
  OAI22_X1 U572 ( .A1(n543), .A2(n400), .B1(n399), .B2(n530), .ZN(n321) );
  XNOR2_X1 U573 ( .A(n501), .B(n559), .ZN(n352) );
  OAI22_X1 U574 ( .A1(n42), .A2(n579), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U575 ( .A1(n559), .A2(n579), .ZN(n332) );
  OAI22_X1 U576 ( .A1(n6), .A2(n404), .B1(n403), .B2(n561), .ZN(n325) );
  OAI22_X1 U577 ( .A1(n543), .A2(n508), .B1(n397), .B2(n530), .ZN(n319) );
  XNOR2_X1 U578 ( .A(n574), .B(n559), .ZN(n343) );
  XOR2_X1 U579 ( .A(n572), .B(a[8]), .Z(n429) );
  XNOR2_X1 U580 ( .A(n155), .B(n555), .ZN(n139) );
  XNOR2_X1 U581 ( .A(n153), .B(n141), .ZN(n555) );
  XNOR2_X1 U582 ( .A(n157), .B(n556), .ZN(n141) );
  XNOR2_X1 U583 ( .A(n145), .B(n143), .ZN(n556) );
  XOR2_X1 U584 ( .A(n315), .B(n261), .Z(n150) );
  OAI22_X1 U585 ( .A1(n544), .A2(n394), .B1(n393), .B2(n530), .ZN(n315) );
  AND2_X1 U586 ( .A1(n560), .A2(n540), .ZN(n300) );
  OAI22_X1 U587 ( .A1(n6), .A2(n405), .B1(n404), .B2(n561), .ZN(n326) );
  XNOR2_X1 U588 ( .A(n576), .B(n559), .ZN(n336) );
  AND2_X1 U589 ( .A1(n560), .A2(n525), .ZN(n314) );
  NAND2_X1 U590 ( .A1(n427), .A2(n37), .ZN(n39) );
  XOR2_X1 U591 ( .A(n576), .B(a[12]), .Z(n427) );
  AND2_X1 U592 ( .A1(n560), .A2(n534), .ZN(n278) );
  OAI22_X1 U593 ( .A1(n544), .A2(n401), .B1(n400), .B2(n530), .ZN(n322) );
  OAI22_X1 U594 ( .A1(n39), .A2(n336), .B1(n37), .B2(n335), .ZN(n263) );
  AND2_X1 U595 ( .A1(n560), .A2(n503), .ZN(n264) );
  OAI22_X1 U596 ( .A1(n544), .A2(n397), .B1(n396), .B2(n530), .ZN(n318) );
  AND2_X1 U597 ( .A1(n560), .A2(n547), .ZN(n288) );
  OAI22_X1 U598 ( .A1(n403), .A2(n6), .B1(n402), .B2(n561), .ZN(n324) );
  AND2_X1 U599 ( .A1(n560), .A2(n538), .ZN(n270) );
  OAI22_X1 U600 ( .A1(n544), .A2(n399), .B1(n398), .B2(n530), .ZN(n320) );
  AND2_X1 U601 ( .A1(n560), .A2(n235), .ZN(n260) );
  OAI22_X1 U602 ( .A1(n543), .A2(n395), .B1(n394), .B2(n530), .ZN(n316) );
  OAI22_X1 U603 ( .A1(n39), .A2(n335), .B1(n37), .B2(n334), .ZN(n262) );
  INV_X1 U604 ( .A(n25), .ZN(n573) );
  NAND2_X1 U605 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U606 ( .A(n578), .B(a[14]), .Z(n426) );
  INV_X1 U607 ( .A(n13), .ZN(n570) );
  INV_X1 U608 ( .A(n7), .ZN(n567) );
  OAI22_X1 U609 ( .A1(n544), .A2(n402), .B1(n401), .B2(n530), .ZN(n323) );
  XNOR2_X1 U610 ( .A(n515), .B(n559), .ZN(n363) );
  OAI22_X1 U611 ( .A1(n543), .A2(n396), .B1(n395), .B2(n530), .ZN(n317) );
  OAI22_X1 U612 ( .A1(n39), .A2(n577), .B1(n337), .B2(n37), .ZN(n252) );
  OR2_X1 U613 ( .A1(n559), .A2(n577), .ZN(n337) );
  AND2_X1 U614 ( .A1(n560), .A2(n249), .ZN(product[0]) );
  OR2_X1 U615 ( .A1(n559), .A2(n575), .ZN(n344) );
  OR2_X1 U616 ( .A1(n559), .A2(n571), .ZN(n364) );
  OR2_X1 U617 ( .A1(n559), .A2(n492), .ZN(n353) );
  OR2_X1 U618 ( .A1(n559), .A2(n532), .ZN(n377) );
  XNOR2_X1 U619 ( .A(n515), .B(b[9]), .ZN(n354) );
  OAI22_X1 U620 ( .A1(n39), .A2(n334), .B1(n37), .B2(n333), .ZN(n261) );
  XNOR2_X1 U621 ( .A(n576), .B(n422), .ZN(n333) );
  XNOR2_X1 U622 ( .A(n569), .B(b[11]), .ZN(n365) );
  XNOR2_X1 U623 ( .A(n576), .B(n424), .ZN(n335) );
  XNOR2_X1 U624 ( .A(n576), .B(n423), .ZN(n334) );
  OAI22_X1 U625 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U626 ( .A(n578), .B(n424), .ZN(n330) );
  XNOR2_X1 U627 ( .A(n578), .B(n559), .ZN(n331) );
  XNOR2_X1 U628 ( .A(n563), .B(b[11]), .ZN(n397) );
  XNOR2_X1 U629 ( .A(n563), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U630 ( .A(n563), .B(b[13]), .ZN(n395) );
  XNOR2_X1 U631 ( .A(n563), .B(b[14]), .ZN(n394) );
  XNOR2_X1 U632 ( .A(n501), .B(n418), .ZN(n345) );
  XNOR2_X1 U633 ( .A(n574), .B(n420), .ZN(n338) );
  XNOR2_X1 U634 ( .A(n565), .B(b[13]), .ZN(n378) );
  XNOR2_X1 U635 ( .A(n515), .B(n424), .ZN(n362) );
  XNOR2_X1 U636 ( .A(n574), .B(n424), .ZN(n342) );
  XNOR2_X1 U637 ( .A(n502), .B(n424), .ZN(n351) );
  XNOR2_X1 U638 ( .A(n574), .B(n423), .ZN(n341) );
  XNOR2_X1 U639 ( .A(n574), .B(n422), .ZN(n340) );
  XNOR2_X1 U640 ( .A(n574), .B(n421), .ZN(n339) );
  XNOR2_X1 U641 ( .A(n566), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U642 ( .A(n566), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U643 ( .A(n565), .B(n418), .ZN(n384) );
  XNOR2_X1 U644 ( .A(n565), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U645 ( .A(n565), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U646 ( .A(n565), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U647 ( .A(n565), .B(n419), .ZN(n385) );
  XNOR2_X1 U648 ( .A(n569), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U649 ( .A(n569), .B(n418), .ZN(n369) );
  XNOR2_X1 U650 ( .A(n569), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U651 ( .A(n569), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U652 ( .A(n501), .B(n423), .ZN(n350) );
  XNOR2_X1 U653 ( .A(n515), .B(n422), .ZN(n360) );
  XNOR2_X1 U654 ( .A(n501), .B(n422), .ZN(n349) );
  XNOR2_X1 U655 ( .A(n515), .B(n423), .ZN(n361) );
  XNOR2_X1 U656 ( .A(n515), .B(n421), .ZN(n359) );
  XNOR2_X1 U657 ( .A(n515), .B(n420), .ZN(n358) );
  XNOR2_X1 U658 ( .A(n502), .B(n421), .ZN(n348) );
  XNOR2_X1 U659 ( .A(n502), .B(n420), .ZN(n347) );
  XNOR2_X1 U660 ( .A(n515), .B(n418), .ZN(n356) );
  XNOR2_X1 U661 ( .A(n502), .B(n419), .ZN(n346) );
  XNOR2_X1 U662 ( .A(n515), .B(n419), .ZN(n357) );
  XNOR2_X1 U663 ( .A(n515), .B(b[8]), .ZN(n355) );
  XNOR2_X1 U664 ( .A(n563), .B(b[15]), .ZN(n393) );
  BUF_X1 U665 ( .A(n43), .Z(n560) );
  OAI22_X1 U666 ( .A1(n520), .A2(n339), .B1(n338), .B2(n507), .ZN(n265) );
  OAI22_X1 U667 ( .A1(n520), .A2(n340), .B1(n339), .B2(n507), .ZN(n266) );
  OAI22_X1 U668 ( .A1(n520), .A2(n341), .B1(n340), .B2(n507), .ZN(n267) );
  OAI22_X1 U669 ( .A1(n520), .A2(n342), .B1(n341), .B2(n507), .ZN(n268) );
  OAI22_X1 U670 ( .A1(n34), .A2(n343), .B1(n507), .B2(n342), .ZN(n269) );
  OAI22_X1 U671 ( .A1(n34), .A2(n575), .B1(n344), .B2(n507), .ZN(n253) );
  NAND2_X1 U672 ( .A1(n428), .A2(n32), .ZN(n34) );
  XNOR2_X1 U673 ( .A(n558), .B(n45), .ZN(product[12]) );
  AND2_X1 U674 ( .A1(n126), .A2(n79), .ZN(n558) );
  INV_X1 U675 ( .A(n19), .ZN(n571) );
  NOR2_X1 U676 ( .A1(n204), .A2(n211), .ZN(n89) );
  OAI22_X1 U677 ( .A1(n500), .A2(n350), .B1(n349), .B2(n526), .ZN(n275) );
  OAI22_X1 U678 ( .A1(n29), .A2(n346), .B1(n345), .B2(n526), .ZN(n271) );
  OAI22_X1 U679 ( .A1(n500), .A2(n347), .B1(n346), .B2(n526), .ZN(n272) );
  OAI22_X1 U680 ( .A1(n539), .A2(n348), .B1(n347), .B2(n526), .ZN(n273) );
  OAI22_X1 U681 ( .A1(n29), .A2(n349), .B1(n348), .B2(n526), .ZN(n274) );
  OAI22_X1 U682 ( .A1(n539), .A2(n492), .B1(n353), .B2(n526), .ZN(n254) );
  OAI22_X1 U683 ( .A1(n539), .A2(n351), .B1(n350), .B2(n526), .ZN(n276) );
  OAI22_X1 U684 ( .A1(n29), .A2(n352), .B1(n351), .B2(n526), .ZN(n277) );
  OAI21_X1 U685 ( .B1(n87), .B2(n85), .A(n86), .ZN(n84) );
  NAND2_X1 U686 ( .A1(n151), .A2(n139), .ZN(n62) );
  XOR2_X1 U687 ( .A(n58), .B(n115), .Z(product[3]) );
  NAND2_X1 U688 ( .A1(n135), .A2(n114), .ZN(n58) );
  INV_X1 U689 ( .A(n88), .ZN(n87) );
  INV_X1 U690 ( .A(n564), .ZN(n563) );
  OR2_X1 U691 ( .A1(n559), .A2(n518), .ZN(n409) );
  XNOR2_X1 U692 ( .A(n77), .B(n48), .ZN(product[13]) );
  OAI22_X1 U693 ( .A1(n505), .A2(n358), .B1(n357), .B2(n495), .ZN(n282) );
  OAI22_X1 U694 ( .A1(n504), .A2(n356), .B1(n355), .B2(n495), .ZN(n280) );
  OAI22_X1 U695 ( .A1(n504), .A2(n362), .B1(n361), .B2(n495), .ZN(n286) );
  OAI22_X1 U696 ( .A1(n504), .A2(n357), .B1(n356), .B2(n21), .ZN(n281) );
  OAI22_X1 U697 ( .A1(n504), .A2(n360), .B1(n359), .B2(n21), .ZN(n284) );
  OAI22_X1 U698 ( .A1(n505), .A2(n571), .B1(n364), .B2(n495), .ZN(n255) );
  OAI22_X1 U699 ( .A1(n505), .A2(n361), .B1(n360), .B2(n495), .ZN(n285) );
  OAI22_X1 U700 ( .A1(n23), .A2(n363), .B1(n362), .B2(n21), .ZN(n287) );
  XNOR2_X1 U701 ( .A(n568), .B(n424), .ZN(n375) );
  OAI22_X1 U702 ( .A1(n505), .A2(n355), .B1(n354), .B2(n21), .ZN(n279) );
  OAI22_X1 U703 ( .A1(n23), .A2(n359), .B1(n358), .B2(n21), .ZN(n283) );
  XNOR2_X1 U704 ( .A(n568), .B(n421), .ZN(n372) );
  XNOR2_X1 U705 ( .A(n568), .B(n423), .ZN(n374) );
  XNOR2_X1 U706 ( .A(n568), .B(n422), .ZN(n373) );
  XNOR2_X1 U707 ( .A(n568), .B(n419), .ZN(n370) );
  XNOR2_X1 U708 ( .A(n568), .B(n420), .ZN(n371) );
  XNOR2_X1 U709 ( .A(n55), .B(n542), .ZN(product[6]) );
  XOR2_X1 U710 ( .A(n529), .B(n54), .Z(product[7]) );
  OAI21_X1 U711 ( .B1(n99), .B2(n97), .A(n98), .ZN(n96) );
  AOI21_X1 U712 ( .B1(n550), .B2(n104), .A(n545), .ZN(n99) );
  XNOR2_X1 U713 ( .A(n541), .B(n53), .ZN(product[8]) );
  OAI22_X1 U714 ( .A1(n512), .A2(n367), .B1(n366), .B2(n16), .ZN(n290) );
  OAI22_X1 U715 ( .A1(n512), .A2(n370), .B1(n369), .B2(n16), .ZN(n293) );
  OAI22_X1 U716 ( .A1(n18), .A2(n368), .B1(n367), .B2(n16), .ZN(n291) );
  OAI22_X1 U717 ( .A1(n512), .A2(n371), .B1(n370), .B2(n16), .ZN(n294) );
  OAI22_X1 U718 ( .A1(n18), .A2(n373), .B1(n372), .B2(n16), .ZN(n296) );
  OAI22_X1 U719 ( .A1(n18), .A2(n369), .B1(n368), .B2(n16), .ZN(n292) );
  OAI22_X1 U720 ( .A1(n18), .A2(n375), .B1(n374), .B2(n16), .ZN(n298) );
  OAI22_X1 U721 ( .A1(n18), .A2(n372), .B1(n371), .B2(n16), .ZN(n295) );
  OAI22_X1 U722 ( .A1(n512), .A2(n374), .B1(n373), .B2(n16), .ZN(n297) );
  OAI22_X1 U723 ( .A1(n18), .A2(n376), .B1(n375), .B2(n16), .ZN(n299) );
  OAI22_X1 U724 ( .A1(n512), .A2(n532), .B1(n377), .B2(n16), .ZN(n256) );
  OAI22_X1 U725 ( .A1(n512), .A2(n366), .B1(n365), .B2(n16), .ZN(n289) );
  XNOR2_X1 U726 ( .A(n565), .B(n420), .ZN(n386) );
  XNOR2_X1 U727 ( .A(n565), .B(n559), .ZN(n391) );
  XNOR2_X1 U728 ( .A(n566), .B(n422), .ZN(n388) );
  XNOR2_X1 U729 ( .A(n566), .B(n424), .ZN(n390) );
  XNOR2_X1 U730 ( .A(n566), .B(n423), .ZN(n389) );
  XNOR2_X1 U731 ( .A(n566), .B(n421), .ZN(n387) );
  XNOR2_X1 U732 ( .A(n523), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U733 ( .A(n522), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U734 ( .A(n522), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U735 ( .A(n523), .B(n418), .ZN(n401) );
  XNOR2_X1 U736 ( .A(n521), .B(n420), .ZN(n403) );
  XNOR2_X1 U737 ( .A(n523), .B(n421), .ZN(n404) );
  XNOR2_X1 U738 ( .A(n522), .B(n422), .ZN(n405) );
  XNOR2_X1 U739 ( .A(n521), .B(n419), .ZN(n402) );
  XNOR2_X1 U740 ( .A(n523), .B(n559), .ZN(n408) );
  XNOR2_X1 U741 ( .A(n523), .B(n424), .ZN(n407) );
  XNOR2_X1 U742 ( .A(n522), .B(n423), .ZN(n406) );
  OAI21_X1 U743 ( .B1(n64), .B2(n546), .A(n65), .ZN(n63) );
  OAI21_X1 U744 ( .B1(n546), .B2(n71), .A(n72), .ZN(n70) );
  OAI21_X1 U745 ( .B1(n78), .B2(n546), .A(n79), .ZN(n77) );
  XOR2_X1 U746 ( .A(n56), .B(n536), .Z(product[5]) );
  NAND2_X1 U747 ( .A1(n329), .A2(n258), .ZN(n122) );
  INV_X1 U748 ( .A(n111), .ZN(n109) );
  OAI22_X1 U749 ( .A1(n543), .A2(n518), .B1(n409), .B2(n530), .ZN(n258) );
  OAI22_X1 U750 ( .A1(n516), .A2(n379), .B1(n378), .B2(n519), .ZN(n301) );
  OAI22_X1 U751 ( .A1(n517), .A2(n380), .B1(n379), .B2(n519), .ZN(n302) );
  OAI22_X1 U752 ( .A1(n517), .A2(n385), .B1(n384), .B2(n519), .ZN(n307) );
  OAI22_X1 U753 ( .A1(n516), .A2(n382), .B1(n381), .B2(n519), .ZN(n304) );
  OAI22_X1 U754 ( .A1(n517), .A2(n381), .B1(n380), .B2(n519), .ZN(n303) );
  NAND2_X1 U755 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U756 ( .A1(n12), .A2(n383), .B1(n382), .B2(n557), .ZN(n305) );
  OAI22_X1 U757 ( .A1(n517), .A2(n384), .B1(n383), .B2(n519), .ZN(n306) );
  OAI22_X1 U758 ( .A1(n516), .A2(n386), .B1(n385), .B2(n519), .ZN(n308) );
  OAI22_X1 U759 ( .A1(n516), .A2(n387), .B1(n386), .B2(n519), .ZN(n309) );
  OAI22_X1 U760 ( .A1(n516), .A2(n510), .B1(n392), .B2(n519), .ZN(n257) );
  OAI22_X1 U761 ( .A1(n12), .A2(n389), .B1(n388), .B2(n557), .ZN(n311) );
  OAI22_X1 U762 ( .A1(n12), .A2(n388), .B1(n557), .B2(n387), .ZN(n310) );
  OAI22_X1 U763 ( .A1(n12), .A2(n390), .B1(n389), .B2(n557), .ZN(n312) );
  OAI22_X1 U764 ( .A1(n517), .A2(n391), .B1(n390), .B2(n519), .ZN(n313) );
  INV_X1 U765 ( .A(n567), .ZN(n566) );
  INV_X1 U766 ( .A(n570), .ZN(n569) );
  INV_X1 U767 ( .A(n31), .ZN(n575) );
  INV_X1 U768 ( .A(n36), .ZN(n577) );
  INV_X1 U769 ( .A(n579), .ZN(n578) );
  INV_X1 U770 ( .A(n40), .ZN(n579) );
  XOR2_X1 U771 ( .A(n259), .B(n251), .Z(n148) );
  XOR2_X1 U772 ( .A(n289), .B(n279), .Z(n146) );
  XOR2_X1 U773 ( .A(n159), .B(n150), .Z(n142) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_7_DW01_add_2 ( A, B, CI, SUM, 
        CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n7, n8, n9, n10, n11, n12, n13, n14, n15, n18, n19,
         n20, n21, n25, n26, n27, n28, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n48, n49, n51, n53, n54, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n69, n71, n72, n73, n74, n75, n77,
         n79, n80, n81, n82, n83, n85, n87, n88, n90, n98, n99, n100, n102,
         n104, n161, n162, n163, n164, n165, n166, n167, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187;

  OAI21_X1 U126 ( .B1(n40), .B2(n36), .A(n37), .ZN(n161) );
  AOI21_X1 U127 ( .B1(n56), .B2(n64), .A(n57), .ZN(n162) );
  AOI21_X1 U128 ( .B1(n56), .B2(n64), .A(n57), .ZN(n163) );
  OR2_X1 U129 ( .A1(A[11]), .A2(B[11]), .ZN(n164) );
  XNOR2_X1 U130 ( .A(n41), .B(n165), .ZN(SUM[11]) );
  AND2_X1 U131 ( .A1(n164), .A2(n40), .ZN(n165) );
  INV_X1 U132 ( .A(n164), .ZN(n166) );
  OR2_X1 U133 ( .A1(A[12]), .A2(B[12]), .ZN(n167) );
  AND2_X1 U134 ( .A1(n179), .A2(n90), .ZN(SUM[0]) );
  XNOR2_X1 U135 ( .A(n49), .B(n169), .ZN(SUM[10]) );
  AND2_X1 U136 ( .A1(n185), .A2(n48), .ZN(n169) );
  OR2_X1 U137 ( .A1(A[15]), .A2(B[15]), .ZN(n170) );
  NOR2_X1 U138 ( .A1(A[11]), .A2(B[11]), .ZN(n39) );
  AOI21_X1 U139 ( .B1(n185), .B2(n51), .A(n186), .ZN(n171) );
  OAI21_X1 U140 ( .B1(n43), .B2(n162), .A(n44), .ZN(n172) );
  NOR2_X1 U141 ( .A1(A[8]), .A2(B[8]), .ZN(n173) );
  NOR2_X1 U142 ( .A1(A[12]), .A2(B[12]), .ZN(n174) );
  NOR2_X1 U143 ( .A1(A[12]), .A2(B[12]), .ZN(n36) );
  OR2_X1 U144 ( .A1(A[14]), .A2(B[14]), .ZN(n175) );
  OR2_X1 U145 ( .A1(A[13]), .A2(B[13]), .ZN(n176) );
  AND2_X1 U146 ( .A1(A[13]), .A2(B[13]), .ZN(n177) );
  OR2_X2 U147 ( .A1(A[10]), .A2(B[10]), .ZN(n185) );
  AOI21_X1 U148 ( .B1(n42), .B2(n34), .A(n35), .ZN(n178) );
  OR2_X1 U149 ( .A1(A[0]), .A2(B[0]), .ZN(n179) );
  INV_X1 U150 ( .A(n64), .ZN(n63) );
  INV_X1 U151 ( .A(n163), .ZN(n54) );
  INV_X1 U152 ( .A(n79), .ZN(n77) );
  OAI21_X1 U153 ( .B1(n67), .B2(n65), .A(n66), .ZN(n64) );
  AOI21_X1 U154 ( .B1(n172), .B2(n34), .A(n161), .ZN(n33) );
  AOI21_X1 U155 ( .B1(n180), .B2(n88), .A(n85), .ZN(n83) );
  INV_X1 U156 ( .A(n87), .ZN(n85) );
  AOI21_X1 U157 ( .B1(n54), .B2(n183), .A(n51), .ZN(n49) );
  OAI21_X1 U158 ( .B1(n83), .B2(n81), .A(n82), .ZN(n80) );
  INV_X1 U159 ( .A(n90), .ZN(n88) );
  OAI21_X1 U160 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  NAND2_X1 U161 ( .A1(n104), .A2(n82), .ZN(n14) );
  INV_X1 U162 ( .A(n81), .ZN(n104) );
  NAND2_X1 U163 ( .A1(n100), .A2(n66), .ZN(n10) );
  INV_X1 U164 ( .A(n65), .ZN(n100) );
  NAND2_X1 U165 ( .A1(n99), .A2(n62), .ZN(n9) );
  INV_X1 U166 ( .A(n61), .ZN(n99) );
  NAND2_X1 U167 ( .A1(n98), .A2(n59), .ZN(n8) );
  NAND2_X1 U168 ( .A1(n182), .A2(n71), .ZN(n11) );
  NAND2_X1 U169 ( .A1(n180), .A2(n87), .ZN(n15) );
  NAND2_X1 U170 ( .A1(n184), .A2(n79), .ZN(n13) );
  AOI21_X1 U171 ( .B1(n182), .B2(n72), .A(n69), .ZN(n67) );
  INV_X1 U172 ( .A(n71), .ZN(n69) );
  NAND2_X1 U173 ( .A1(n102), .A2(n74), .ZN(n12) );
  INV_X1 U174 ( .A(n73), .ZN(n102) );
  INV_X1 U175 ( .A(n187), .ZN(n25) );
  XOR2_X1 U176 ( .A(n14), .B(n83), .Z(SUM[2]) );
  NAND2_X1 U177 ( .A1(n176), .A2(n28), .ZN(n3) );
  NOR2_X1 U178 ( .A1(A[7]), .A2(B[7]), .ZN(n61) );
  NOR2_X1 U179 ( .A1(A[2]), .A2(B[2]), .ZN(n81) );
  NAND2_X1 U180 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  OR2_X1 U181 ( .A1(A[1]), .A2(B[1]), .ZN(n180) );
  NOR2_X1 U182 ( .A1(A[6]), .A2(B[6]), .ZN(n65) );
  OR2_X1 U183 ( .A1(A[14]), .A2(B[14]), .ZN(n181) );
  XNOR2_X1 U184 ( .A(n60), .B(n8), .ZN(SUM[8]) );
  NOR2_X1 U185 ( .A1(A[4]), .A2(B[4]), .ZN(n73) );
  NAND2_X1 U186 ( .A1(A[7]), .A2(B[7]), .ZN(n62) );
  OR2_X1 U187 ( .A1(A[5]), .A2(B[5]), .ZN(n182) );
  NAND2_X1 U188 ( .A1(A[2]), .A2(B[2]), .ZN(n82) );
  OR2_X1 U189 ( .A1(A[9]), .A2(B[9]), .ZN(n183) );
  NAND2_X1 U190 ( .A1(A[5]), .A2(B[5]), .ZN(n71) );
  NAND2_X1 U191 ( .A1(A[1]), .A2(B[1]), .ZN(n87) );
  NAND2_X1 U192 ( .A1(A[0]), .A2(B[0]), .ZN(n90) );
  NAND2_X1 U193 ( .A1(A[6]), .A2(B[6]), .ZN(n66) );
  OR2_X1 U194 ( .A1(A[3]), .A2(B[3]), .ZN(n184) );
  NAND2_X1 U195 ( .A1(A[4]), .A2(B[4]), .ZN(n74) );
  NAND2_X1 U196 ( .A1(A[3]), .A2(B[3]), .ZN(n79) );
  NAND2_X1 U197 ( .A1(A[8]), .A2(B[8]), .ZN(n59) );
  NAND2_X1 U198 ( .A1(A[9]), .A2(B[9]), .ZN(n53) );
  XNOR2_X1 U199 ( .A(n54), .B(n7), .ZN(SUM[9]) );
  XOR2_X1 U200 ( .A(n63), .B(n9), .Z(SUM[7]) );
  XNOR2_X1 U201 ( .A(n11), .B(n72), .ZN(SUM[5]) );
  XNOR2_X1 U202 ( .A(n13), .B(n80), .ZN(SUM[3]) );
  XNOR2_X1 U203 ( .A(n15), .B(n88), .ZN(SUM[1]) );
  NAND2_X1 U204 ( .A1(n170), .A2(n18), .ZN(n1) );
  INV_X1 U205 ( .A(n173), .ZN(n98) );
  NOR2_X1 U206 ( .A1(n173), .A2(n61), .ZN(n56) );
  OAI21_X1 U207 ( .B1(n58), .B2(n62), .A(n59), .ZN(n57) );
  NOR2_X1 U208 ( .A1(A[8]), .A2(B[8]), .ZN(n58) );
  INV_X1 U209 ( .A(n186), .ZN(n48) );
  XOR2_X1 U210 ( .A(n10), .B(n67), .Z(SUM[6]) );
  NAND2_X1 U211 ( .A1(A[12]), .A2(B[12]), .ZN(n37) );
  NAND2_X1 U212 ( .A1(n167), .A2(n37), .ZN(n4) );
  AND2_X1 U213 ( .A1(A[10]), .A2(B[10]), .ZN(n186) );
  NAND2_X1 U214 ( .A1(n183), .A2(n53), .ZN(n7) );
  INV_X1 U215 ( .A(n53), .ZN(n51) );
  NAND2_X1 U216 ( .A1(A[11]), .A2(B[11]), .ZN(n40) );
  NAND2_X1 U217 ( .A1(n175), .A2(n25), .ZN(n2) );
  NAND2_X1 U218 ( .A1(n175), .A2(n176), .ZN(n20) );
  AOI21_X1 U219 ( .B1(n181), .B2(n177), .A(n187), .ZN(n21) );
  AND2_X1 U220 ( .A1(A[14]), .A2(B[14]), .ZN(n187) );
  AOI21_X1 U221 ( .B1(n184), .B2(n80), .A(n77), .ZN(n75) );
  XOR2_X1 U222 ( .A(n12), .B(n75), .Z(SUM[4]) );
  OAI21_X1 U223 ( .B1(n75), .B2(n73), .A(n74), .ZN(n72) );
  OAI21_X1 U224 ( .B1(n40), .B2(n36), .A(n37), .ZN(n35) );
  NOR2_X1 U225 ( .A1(A[13]), .A2(B[13]), .ZN(n27) );
  OAI21_X1 U226 ( .B1(n41), .B2(n166), .A(n40), .ZN(n38) );
  NOR2_X1 U227 ( .A1(n174), .A2(n39), .ZN(n34) );
  XNOR2_X1 U228 ( .A(n26), .B(n2), .ZN(SUM[14]) );
  NAND2_X1 U229 ( .A1(A[15]), .A2(B[15]), .ZN(n18) );
  INV_X1 U230 ( .A(n172), .ZN(n41) );
  NAND2_X1 U231 ( .A1(n185), .A2(n183), .ZN(n43) );
  AOI21_X1 U232 ( .B1(n185), .B2(n51), .A(n186), .ZN(n44) );
  XNOR2_X1 U233 ( .A(n38), .B(n4), .ZN(SUM[12]) );
  XNOR2_X1 U234 ( .A(n19), .B(n1), .ZN(SUM[15]) );
  XOR2_X1 U235 ( .A(n33), .B(n3), .Z(SUM[13]) );
  OAI21_X1 U236 ( .B1(n178), .B2(n27), .A(n28), .ZN(n26) );
  OAI21_X1 U237 ( .B1(n178), .B2(n20), .A(n21), .ZN(n19) );
  OAI21_X1 U238 ( .B1(n43), .B2(n162), .A(n171), .ZN(n42) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_7 ( clk, clear_acc, 
        data_out_x, data_out, data_out_w, data_out_b, wr_en_y, m_valid, 
        m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [3:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N27, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, n1, n2, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n87, n104, n113, n114, n115, n116, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n17), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n223), .CK(clk), .Q(n22) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n224), .CK(clk), .Q(n23) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n225), .CK(clk), .Q(n24) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n226), .CK(clk), .Q(n25) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n227), .CK(clk), .Q(n26) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n228), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n229), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n230), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n231), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n232), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n233), .CK(clk), .Q(n34) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n234), .CK(clk), .Q(n35) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n235), .CK(clk), .Q(n36) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n236), .CK(clk), .Q(n37) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n237), .CK(clk), .Q(n38) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n238), .CK(clk), .Q(n40) );
  DFF_X1 \f_reg[8]  ( .D(n81), .CK(clk), .Q(f[8]), .QN(n216) );
  DFF_X1 \f_reg[9]  ( .D(n80), .CK(clk), .Q(f[9]), .QN(n217) );
  DFF_X1 \f_reg[10]  ( .D(n79), .CK(clk), .Q(n51), .QN(n218) );
  DFF_X1 \f_reg[11]  ( .D(n78), .CK(clk), .Q(n49), .QN(n219) );
  DFF_X1 \f_reg[12]  ( .D(n1), .CK(clk), .Q(n48), .QN(n220) );
  DFF_X1 \f_reg[13]  ( .D(n77), .CK(clk), .Q(n46), .QN(n221) );
  DFF_X1 \f_reg[14]  ( .D(n4), .CK(clk), .Q(n45), .QN(n222) );
  DFF_X1 \f_reg[15]  ( .D(n2), .CK(clk), .Q(n44), .QN(n75) );
  DFF_X1 \data_out_reg[15]  ( .D(n115), .CK(clk), .Q(data_out[15]), .QN(n195)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n116), .CK(clk), .Q(data_out[14]), .QN(n194)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n166), .CK(clk), .Q(data_out[13]), .QN(n193)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n167), .CK(clk), .Q(data_out[12]), .QN(n192)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n168), .CK(clk), .Q(data_out[11]), .QN(n191)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n169), .CK(clk), .Q(data_out[10]), .QN(n190)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n170), .CK(clk), .Q(data_out[9]), .QN(n189) );
  DFF_X1 \data_out_reg[8]  ( .D(n171), .CK(clk), .Q(data_out[8]), .QN(n188) );
  DFF_X1 \data_out_reg[7]  ( .D(n172), .CK(clk), .Q(data_out[7]), .QN(n187) );
  DFF_X1 \data_out_reg[6]  ( .D(n173), .CK(clk), .Q(data_out[6]), .QN(n186) );
  DFF_X1 \data_out_reg[5]  ( .D(n174), .CK(clk), .Q(data_out[5]), .QN(n185) );
  DFF_X1 \data_out_reg[4]  ( .D(n175), .CK(clk), .Q(data_out[4]), .QN(n184) );
  DFF_X1 \data_out_reg[3]  ( .D(n176), .CK(clk), .Q(data_out[3]), .QN(n183) );
  DFF_X1 \data_out_reg[2]  ( .D(n177), .CK(clk), .Q(data_out[2]), .QN(n182) );
  DFF_X1 \data_out_reg[1]  ( .D(n178), .CK(clk), .Q(data_out[1]), .QN(n181) );
  DFF_X1 \data_out_reg[0]  ( .D(n179), .CK(clk), .Q(data_out[0]), .QN(n180) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_7_DW_mult_tc_1 mult_960 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_7_DW01_add_2 add_961 ( .A({n202, 
        n201, n200, n199, n198, n197, n211, n210, n209, n208, n207, n206, n205, 
        n204, n203, n196}), .B({n44, n45, n46, n48, n49, n51, f[9:3], n59, n61, 
        n63}), .CI(1'b0), .SUM(adder) );
  DFF_X2 delay_reg ( .D(N27), .CK(clk), .Q(n14), .QN(n239) );
  DFF_X1 \f_reg[3]  ( .D(n87), .CK(clk), .Q(f[3]), .QN(n67) );
  DFF_X1 \f_reg[1]  ( .D(n113), .CK(clk), .Q(n61), .QN(n213) );
  DFF_X1 \f_reg[4]  ( .D(n85), .CK(clk), .Q(f[4]), .QN(n68) );
  DFF_X1 \f_reg[2]  ( .D(n104), .CK(clk), .Q(n59), .QN(n214) );
  DFF_X1 \f_reg[0]  ( .D(n114), .CK(clk), .Q(n63), .QN(n212) );
  DFF_X1 \f_reg[5]  ( .D(n84), .CK(clk), .Q(f[5]), .QN(n69) );
  DFF_X1 \f_reg[6]  ( .D(n83), .CK(clk), .Q(f[6]), .QN(n70) );
  DFF_X1 \f_reg[7]  ( .D(n82), .CK(clk), .Q(f[7]), .QN(n215) );
  AND2_X2 U3 ( .A1(n43), .A2(n18), .ZN(n15) );
  MUX2_X1 U4 ( .A(N40), .B(n26), .S(n14), .Z(n198) );
  MUX2_X2 U5 ( .A(n23), .B(N43), .S(n239), .Z(n201) );
  NAND3_X1 U6 ( .A1(n6), .A2(n5), .A3(n7), .ZN(n1) );
  NAND3_X1 U8 ( .A1(n12), .A2(n11), .A3(n13), .ZN(n2) );
  NAND3_X1 U9 ( .A1(n9), .A2(n8), .A3(n10), .ZN(n4) );
  MUX2_X1 U10 ( .A(N39), .B(n27), .S(n14), .Z(n197) );
  NAND2_X1 U11 ( .A1(data_out_b[12]), .A2(n17), .ZN(n5) );
  NAND2_X1 U12 ( .A1(adder[12]), .A2(n15), .ZN(n6) );
  NAND2_X1 U13 ( .A1(n65), .A2(n48), .ZN(n7) );
  NAND2_X1 U14 ( .A1(data_out_b[14]), .A2(n17), .ZN(n8) );
  NAND2_X1 U15 ( .A1(adder[14]), .A2(n15), .ZN(n9) );
  NAND2_X1 U16 ( .A1(n65), .A2(n45), .ZN(n10) );
  NAND2_X1 U17 ( .A1(data_out_b[15]), .A2(n17), .ZN(n11) );
  NAND2_X1 U18 ( .A1(adder[15]), .A2(n15), .ZN(n12) );
  NAND2_X1 U19 ( .A1(n65), .A2(n44), .ZN(n13) );
  INV_X2 U20 ( .A(n43), .ZN(n65) );
  MUX2_X2 U21 ( .A(n29), .B(N37), .S(n239), .Z(n210) );
  MUX2_X2 U22 ( .A(n25), .B(N41), .S(n239), .Z(n199) );
  MUX2_X2 U23 ( .A(n24), .B(N42), .S(n239), .Z(n200) );
  INV_X1 U24 ( .A(n18), .ZN(n17) );
  INV_X1 U25 ( .A(clear_acc), .ZN(n18) );
  NAND2_X1 U26 ( .A1(n16), .A2(N27), .ZN(n241) );
  INV_X1 U27 ( .A(n21), .ZN(n39) );
  OAI22_X1 U28 ( .A1(n183), .A2(n241), .B1(n67), .B2(n240), .ZN(n176) );
  OAI22_X1 U29 ( .A1(n184), .A2(n241), .B1(n68), .B2(n240), .ZN(n175) );
  OAI22_X1 U30 ( .A1(n185), .A2(n241), .B1(n69), .B2(n240), .ZN(n174) );
  OAI22_X1 U31 ( .A1(n186), .A2(n241), .B1(n70), .B2(n240), .ZN(n173) );
  OAI22_X1 U32 ( .A1(n187), .A2(n241), .B1(n215), .B2(n240), .ZN(n172) );
  OAI22_X1 U33 ( .A1(n188), .A2(n241), .B1(n216), .B2(n240), .ZN(n171) );
  OAI22_X1 U34 ( .A1(n189), .A2(n241), .B1(n217), .B2(n240), .ZN(n170) );
  MUX2_X1 U35 ( .A(n36), .B(N32), .S(n239), .Z(n205) );
  INV_X1 U36 ( .A(wr_en_y), .ZN(n16) );
  AND2_X1 U37 ( .A1(sel[0]), .A2(sel[1]), .ZN(n20) );
  INV_X1 U38 ( .A(m_ready), .ZN(n19) );
  NAND2_X1 U39 ( .A1(m_valid), .A2(n19), .ZN(n41) );
  OAI211_X1 U40 ( .C1(sel[2]), .C2(n20), .A(sel[3]), .B(n41), .ZN(N27) );
  NAND2_X1 U41 ( .A1(clear_acc_delay), .A2(n239), .ZN(n21) );
  MUX2_X1 U42 ( .A(n22), .B(N44), .S(n39), .Z(n223) );
  MUX2_X1 U43 ( .A(n22), .B(N44), .S(n239), .Z(n202) );
  MUX2_X1 U44 ( .A(n23), .B(N43), .S(n39), .Z(n224) );
  MUX2_X1 U45 ( .A(n24), .B(N42), .S(n39), .Z(n225) );
  MUX2_X1 U46 ( .A(n25), .B(N41), .S(n39), .Z(n226) );
  MUX2_X1 U47 ( .A(n26), .B(N40), .S(n39), .Z(n227) );
  MUX2_X1 U48 ( .A(n27), .B(N39), .S(n39), .Z(n228) );
  MUX2_X1 U49 ( .A(n28), .B(N38), .S(n39), .Z(n229) );
  MUX2_X1 U50 ( .A(n28), .B(N38), .S(n239), .Z(n211) );
  MUX2_X1 U51 ( .A(n29), .B(N37), .S(n39), .Z(n230) );
  MUX2_X1 U52 ( .A(n32), .B(N36), .S(n39), .Z(n231) );
  MUX2_X1 U53 ( .A(n32), .B(N36), .S(n239), .Z(n209) );
  MUX2_X1 U54 ( .A(n33), .B(N35), .S(n39), .Z(n232) );
  MUX2_X1 U55 ( .A(n33), .B(N35), .S(n239), .Z(n208) );
  MUX2_X1 U56 ( .A(n34), .B(N34), .S(n39), .Z(n233) );
  MUX2_X1 U57 ( .A(n34), .B(N34), .S(n239), .Z(n207) );
  MUX2_X1 U58 ( .A(n35), .B(N33), .S(n39), .Z(n234) );
  MUX2_X1 U59 ( .A(n35), .B(N33), .S(n239), .Z(n206) );
  MUX2_X1 U60 ( .A(n36), .B(N32), .S(n39), .Z(n235) );
  MUX2_X1 U61 ( .A(n37), .B(N31), .S(n39), .Z(n236) );
  MUX2_X1 U62 ( .A(n37), .B(N31), .S(n239), .Z(n204) );
  MUX2_X1 U63 ( .A(n38), .B(N30), .S(n39), .Z(n237) );
  MUX2_X1 U64 ( .A(n38), .B(N30), .S(n239), .Z(n203) );
  MUX2_X1 U65 ( .A(n40), .B(N29), .S(n39), .Z(n238) );
  MUX2_X1 U66 ( .A(n40), .B(N29), .S(n239), .Z(n196) );
  INV_X1 U67 ( .A(n41), .ZN(n42) );
  OAI21_X1 U68 ( .B1(n42), .B2(n14), .A(n18), .ZN(n43) );
  AOI222_X1 U69 ( .A1(data_out_b[13]), .A2(n17), .B1(adder[13]), .B2(n15), 
        .C1(n65), .C2(n46), .ZN(n47) );
  INV_X1 U70 ( .A(n47), .ZN(n77) );
  AOI222_X1 U71 ( .A1(data_out_b[11]), .A2(n17), .B1(adder[11]), .B2(n15), 
        .C1(n65), .C2(n49), .ZN(n50) );
  INV_X1 U72 ( .A(n50), .ZN(n78) );
  AOI222_X1 U73 ( .A1(data_out_b[10]), .A2(n17), .B1(adder[10]), .B2(n15), 
        .C1(n65), .C2(n51), .ZN(n52) );
  INV_X1 U74 ( .A(n52), .ZN(n79) );
  AOI222_X1 U75 ( .A1(data_out_b[8]), .A2(n17), .B1(adder[8]), .B2(n15), .C1(
        n65), .C2(f[8]), .ZN(n53) );
  INV_X1 U76 ( .A(n53), .ZN(n81) );
  AOI222_X1 U77 ( .A1(data_out_b[7]), .A2(n17), .B1(adder[7]), .B2(n15), .C1(
        n65), .C2(f[7]), .ZN(n54) );
  INV_X1 U78 ( .A(n54), .ZN(n82) );
  AOI222_X1 U79 ( .A1(data_out_b[6]), .A2(n17), .B1(adder[6]), .B2(n15), .C1(
        n65), .C2(f[6]), .ZN(n55) );
  INV_X1 U80 ( .A(n55), .ZN(n83) );
  AOI222_X1 U81 ( .A1(data_out_b[5]), .A2(n17), .B1(adder[5]), .B2(n15), .C1(
        n65), .C2(f[5]), .ZN(n56) );
  INV_X1 U82 ( .A(n56), .ZN(n84) );
  AOI222_X1 U83 ( .A1(data_out_b[4]), .A2(n17), .B1(adder[4]), .B2(n15), .C1(
        n65), .C2(f[4]), .ZN(n57) );
  INV_X1 U84 ( .A(n57), .ZN(n85) );
  AOI222_X1 U85 ( .A1(data_out_b[3]), .A2(n17), .B1(adder[3]), .B2(n15), .C1(
        n65), .C2(f[3]), .ZN(n58) );
  INV_X1 U86 ( .A(n58), .ZN(n87) );
  AOI222_X1 U87 ( .A1(data_out_b[2]), .A2(n17), .B1(adder[2]), .B2(n15), .C1(
        n65), .C2(n59), .ZN(n60) );
  INV_X1 U88 ( .A(n60), .ZN(n104) );
  AOI222_X1 U89 ( .A1(data_out_b[1]), .A2(n17), .B1(adder[1]), .B2(n15), .C1(
        n65), .C2(n61), .ZN(n62) );
  INV_X1 U90 ( .A(n62), .ZN(n113) );
  AOI222_X1 U91 ( .A1(data_out_b[0]), .A2(n17), .B1(adder[0]), .B2(n15), .C1(
        n65), .C2(n63), .ZN(n64) );
  INV_X1 U92 ( .A(n64), .ZN(n114) );
  AOI222_X1 U93 ( .A1(data_out_b[9]), .A2(n17), .B1(adder[9]), .B2(n15), .C1(
        n65), .C2(f[9]), .ZN(n66) );
  INV_X1 U94 ( .A(n66), .ZN(n80) );
  NOR4_X1 U95 ( .A1(n49), .A2(n48), .A3(n46), .A4(n45), .ZN(n74) );
  NOR4_X1 U96 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n51), .ZN(n73) );
  NAND4_X1 U97 ( .A1(n70), .A2(n69), .A3(n68), .A4(n67), .ZN(n71) );
  NOR4_X1 U98 ( .A1(n71), .A2(n63), .A3(n61), .A4(n59), .ZN(n72) );
  NAND3_X1 U99 ( .A1(n74), .A2(n73), .A3(n72), .ZN(n76) );
  NAND3_X1 U100 ( .A1(wr_en_y), .A2(n76), .A3(n75), .ZN(n240) );
  OAI22_X1 U101 ( .A1(n180), .A2(n241), .B1(n212), .B2(n240), .ZN(n179) );
  OAI22_X1 U102 ( .A1(n181), .A2(n241), .B1(n213), .B2(n240), .ZN(n178) );
  OAI22_X1 U103 ( .A1(n182), .A2(n241), .B1(n214), .B2(n240), .ZN(n177) );
  OAI22_X1 U104 ( .A1(n190), .A2(n241), .B1(n218), .B2(n240), .ZN(n169) );
  OAI22_X1 U105 ( .A1(n191), .A2(n241), .B1(n219), .B2(n240), .ZN(n168) );
  OAI22_X1 U106 ( .A1(n192), .A2(n241), .B1(n220), .B2(n240), .ZN(n167) );
  OAI22_X1 U107 ( .A1(n193), .A2(n241), .B1(n221), .B2(n240), .ZN(n166) );
  OAI22_X1 U108 ( .A1(n194), .A2(n241), .B1(n222), .B2(n240), .ZN(n116) );
  OAI22_X1 U109 ( .A1(n195), .A2(n241), .B1(n75), .B2(n240), .ZN(n115) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_6_DW_mult_tc_1 ( a, b, 
        product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n9, n12, n13, n16, n18, n19, n21, n23, n25, n27, n29, n31,
         n32, n34, n36, n37, n39, n40, n41, n42, n43, n46, n47, n48, n50, n53,
         n54, n55, n56, n57, n58, n59, n62, n63, n64, n65, n67, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n93, n95, n96, n97, n98, n99, n103,
         n104, n105, n106, n107, n111, n112, n113, n114, n115, n117, n119,
         n120, n122, n127, n131, n135, n139, n141, n142, n143, n144, n145,
         n146, n147, n148, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n237, n239, n245, n247, n249, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n418, n419, n420, n421, n422, n423, n424, n426, n427, n428, n432,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U148 ( .A(n265), .B(n144), .Z(n145) );
  XOR2_X1 U150 ( .A(n271), .B(n146), .Z(n147) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U161 ( .A(n177), .B(n168), .CI(n166), .CO(n163), .S(n164) );
  FA_X1 U162 ( .A(n170), .B(n172), .CI(n179), .CO(n165), .S(n166) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n291), .CI(n263), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n317), .B(n252), .CO(n173), .S(n174) );
  FA_X1 U167 ( .A(n180), .B(n187), .CI(n178), .CO(n175), .S(n176) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U170 ( .A(n268), .B(n292), .CI(n274), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U172 ( .A(n197), .B(n190), .CI(n188), .CO(n185), .S(n186) );
  FA_X1 U173 ( .A(n199), .B(n201), .CI(n192), .CO(n187), .S(n188) );
  FA_X1 U174 ( .A(n275), .B(n293), .CI(n194), .CO(n189), .S(n190) );
  FA_X1 U175 ( .A(n305), .B(n253), .CI(n283), .CO(n191), .S(n192) );
  HA_X1 U176 ( .A(n319), .B(n269), .CO(n193), .S(n194) );
  FA_X1 U177 ( .A(n205), .B(n200), .CI(n198), .CO(n195), .S(n196) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U179 ( .A(n294), .B(n284), .CI(n276), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n320), .B(n270), .CI(n306), .CO(n201), .S(n202) );
  FA_X1 U181 ( .A(n208), .B(n213), .CI(n206), .CO(n203), .S(n204) );
  FA_X1 U182 ( .A(n215), .B(n307), .CI(n210), .CO(n205), .S(n206) );
  FA_X1 U183 ( .A(n295), .B(n285), .CI(n254), .CO(n207), .S(n208) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U185 ( .A(n216), .B(n219), .CI(n214), .CO(n211), .S(n212) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n322), .B(n278), .CI(n308), .CO(n215), .S(n216) );
  FA_X1 U188 ( .A(n225), .B(n222), .CI(n220), .CO(n217), .S(n218) );
  FA_X1 U189 ( .A(n297), .B(n309), .CI(n255), .CO(n219), .S(n220) );
  HA_X1 U190 ( .A(n287), .B(n323), .CO(n221), .S(n222) );
  FA_X1 U191 ( .A(n229), .B(n298), .CI(n226), .CO(n223), .S(n224) );
  FA_X1 U192 ( .A(n310), .B(n288), .CI(n324), .CO(n225), .S(n226) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  HA_X1 U194 ( .A(n325), .B(n311), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n312), .B(n326), .CI(n300), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  OR2_X1 U414 ( .A1(n228), .A2(n231), .ZN(n490) );
  XNOR2_X1 U415 ( .A(n554), .B(n491), .ZN(product[9]) );
  AND2_X1 U416 ( .A1(n550), .A2(n90), .ZN(n491) );
  AOI21_X1 U417 ( .B1(n104), .B2(n565), .A(n556), .ZN(n492) );
  AND2_X1 U418 ( .A1(n232), .A2(n233), .ZN(n544) );
  INV_X1 U419 ( .A(n544), .ZN(n111) );
  BUF_X1 U420 ( .A(n497), .Z(n516) );
  INV_X1 U421 ( .A(n549), .ZN(n27) );
  OR2_X1 U422 ( .A1(n164), .A2(n175), .ZN(n493) );
  OR2_X1 U423 ( .A1(n329), .A2(n258), .ZN(n494) );
  CLKBUF_X1 U424 ( .A(n576), .Z(n557) );
  INV_X1 U425 ( .A(n13), .ZN(n495) );
  BUF_X1 U426 ( .A(n18), .Z(n500) );
  BUF_X1 U427 ( .A(n18), .Z(n501) );
  CLKBUF_X1 U428 ( .A(n86), .Z(n496) );
  BUF_X1 U429 ( .A(n535), .Z(n497) );
  CLKBUF_X1 U430 ( .A(n104), .Z(n498) );
  CLKBUF_X1 U431 ( .A(n18), .Z(n499) );
  OR2_X1 U432 ( .A1(n196), .A2(n203), .ZN(n502) );
  XNOR2_X1 U433 ( .A(n503), .B(n147), .ZN(n144) );
  XNOR2_X1 U434 ( .A(n301), .B(n148), .ZN(n503) );
  BUF_X2 U435 ( .A(n32), .Z(n521) );
  NAND2_X1 U436 ( .A1(n432), .A2(n535), .ZN(n504) );
  INV_X1 U437 ( .A(n245), .ZN(n505) );
  BUF_X1 U438 ( .A(n540), .Z(n506) );
  XOR2_X1 U439 ( .A(n193), .B(n282), .Z(n507) );
  XOR2_X1 U440 ( .A(n191), .B(n507), .Z(n180) );
  NAND2_X1 U441 ( .A1(n191), .A2(n193), .ZN(n508) );
  NAND2_X1 U442 ( .A1(n191), .A2(n282), .ZN(n509) );
  NAND2_X1 U443 ( .A1(n193), .A2(n282), .ZN(n510) );
  NAND3_X1 U444 ( .A1(n509), .A2(n508), .A3(n510), .ZN(n179) );
  CLKBUF_X1 U445 ( .A(n501), .Z(n511) );
  BUF_X1 U446 ( .A(n91), .Z(n554) );
  INV_X1 U447 ( .A(n548), .ZN(n21) );
  AOI21_X1 U448 ( .B1(n88), .B2(n80), .A(n81), .ZN(n512) );
  INV_X2 U449 ( .A(n591), .ZN(n590) );
  NOR2_X1 U450 ( .A1(n164), .A2(n175), .ZN(n513) );
  NOR2_X1 U451 ( .A1(n164), .A2(n175), .ZN(n75) );
  CLKBUF_X1 U452 ( .A(n12), .Z(n514) );
  AOI21_X1 U453 ( .B1(n96), .B2(n561), .A(n93), .ZN(n515) );
  AOI21_X1 U454 ( .B1(n96), .B2(n561), .A(n93), .ZN(n91) );
  XNOR2_X1 U455 ( .A(n576), .B(n249), .ZN(n517) );
  INV_X1 U456 ( .A(n526), .ZN(n518) );
  CLKBUF_X1 U457 ( .A(n575), .Z(n519) );
  XNOR2_X1 U458 ( .A(n589), .B(a[10]), .ZN(n428) );
  OR2_X2 U459 ( .A1(n537), .A2(n522), .ZN(n520) );
  INV_X1 U460 ( .A(n577), .ZN(n570) );
  XOR2_X1 U461 ( .A(n587), .B(a[10]), .Z(n32) );
  XNOR2_X1 U462 ( .A(n583), .B(a[6]), .ZN(n522) );
  BUF_X2 U463 ( .A(n584), .Z(n525) );
  INV_X1 U464 ( .A(n502), .ZN(n523) );
  OR2_X2 U465 ( .A1(n524), .A2(n549), .ZN(n29) );
  XNOR2_X1 U466 ( .A(n586), .B(a[8]), .ZN(n524) );
  BUF_X2 U467 ( .A(n584), .Z(n526) );
  INV_X1 U468 ( .A(n585), .ZN(n584) );
  NAND2_X1 U469 ( .A1(n559), .A2(n16), .ZN(n18) );
  INV_X1 U470 ( .A(n519), .ZN(n527) );
  INV_X1 U471 ( .A(n19), .ZN(n585) );
  INV_X1 U472 ( .A(n579), .ZN(n528) );
  INV_X2 U473 ( .A(n580), .ZN(n579) );
  INV_X1 U474 ( .A(n589), .ZN(n529) );
  INV_X1 U475 ( .A(n589), .ZN(n588) );
  XNOR2_X1 U476 ( .A(n495), .B(a[4]), .ZN(n559) );
  INV_X1 U477 ( .A(n583), .ZN(n581) );
  CLKBUF_X1 U478 ( .A(n107), .Z(n530) );
  BUF_X2 U479 ( .A(n9), .Z(n558) );
  OR2_X1 U480 ( .A1(n176), .A2(n185), .ZN(n531) );
  BUF_X1 U481 ( .A(n37), .Z(n532) );
  XNOR2_X1 U482 ( .A(n588), .B(a[12]), .ZN(n37) );
  OAI21_X1 U483 ( .B1(n515), .B2(n89), .A(n90), .ZN(n533) );
  CLKBUF_X1 U484 ( .A(n500), .Z(n534) );
  XNOR2_X1 U485 ( .A(n575), .B(a[2]), .ZN(n535) );
  XNOR2_X1 U486 ( .A(n575), .B(a[2]), .ZN(n9) );
  NOR2_X1 U487 ( .A1(n186), .A2(n195), .ZN(n536) );
  NOR2_X1 U488 ( .A1(n186), .A2(n195), .ZN(n82) );
  OR2_X2 U489 ( .A1(n537), .A2(n522), .ZN(n23) );
  XOR2_X1 U490 ( .A(n585), .B(a[6]), .Z(n537) );
  CLKBUF_X1 U491 ( .A(n96), .Z(n538) );
  NAND2_X1 U492 ( .A1(n428), .A2(n32), .ZN(n539) );
  AOI21_X1 U493 ( .B1(n533), .B2(n80), .A(n81), .ZN(n540) );
  CLKBUF_X1 U494 ( .A(n97), .Z(n541) );
  XNOR2_X1 U495 ( .A(n533), .B(n542), .ZN(product[10]) );
  NAND2_X1 U496 ( .A1(n502), .A2(n86), .ZN(n542) );
  CLKBUF_X1 U497 ( .A(n565), .Z(n543) );
  CLKBUF_X1 U498 ( .A(n224), .Z(n545) );
  INV_X1 U499 ( .A(n13), .ZN(n583) );
  OR2_X2 U500 ( .A1(n553), .A2(n249), .ZN(n546) );
  OR2_X2 U501 ( .A1(n517), .A2(n249), .ZN(n547) );
  OR2_X1 U502 ( .A1(n517), .A2(n249), .ZN(n6) );
  XNOR2_X1 U503 ( .A(n580), .B(a[2]), .ZN(n432) );
  INV_X1 U504 ( .A(n580), .ZN(n578) );
  XNOR2_X1 U505 ( .A(n583), .B(a[6]), .ZN(n548) );
  XNOR2_X1 U506 ( .A(n585), .B(a[8]), .ZN(n549) );
  XOR2_X1 U507 ( .A(n580), .B(a[4]), .Z(n16) );
  OR2_X1 U508 ( .A1(n204), .A2(n211), .ZN(n550) );
  NAND2_X1 U509 ( .A1(n9), .A2(n432), .ZN(n551) );
  NAND2_X1 U510 ( .A1(n432), .A2(n535), .ZN(n552) );
  NAND2_X1 U511 ( .A1(n9), .A2(n432), .ZN(n12) );
  XNOR2_X1 U512 ( .A(n576), .B(n249), .ZN(n553) );
  CLKBUF_X1 U513 ( .A(n492), .Z(n555) );
  AND2_X1 U514 ( .A1(n224), .A2(n227), .ZN(n556) );
  INV_X1 U515 ( .A(n577), .ZN(n576) );
  INV_X2 U516 ( .A(n587), .ZN(n586) );
  CLKBUF_X3 U517 ( .A(n16), .Z(n569) );
  BUF_X1 U518 ( .A(n43), .Z(n572) );
  NAND2_X1 U519 ( .A1(n560), .A2(n69), .ZN(n47) );
  INV_X1 U520 ( .A(n73), .ZN(n71) );
  AOI21_X1 U521 ( .B1(n560), .B2(n74), .A(n67), .ZN(n65) );
  INV_X1 U522 ( .A(n69), .ZN(n67) );
  NAND2_X1 U523 ( .A1(n73), .A2(n560), .ZN(n64) );
  INV_X1 U524 ( .A(n74), .ZN(n72) );
  OR2_X1 U525 ( .A1(n152), .A2(n163), .ZN(n560) );
  INV_X1 U526 ( .A(n95), .ZN(n93) );
  NAND2_X1 U527 ( .A1(n493), .A2(n76), .ZN(n48) );
  OAI21_X1 U528 ( .B1(n513), .B2(n79), .A(n76), .ZN(n74) );
  NOR2_X1 U529 ( .A1(n75), .A2(n78), .ZN(n73) );
  XNOR2_X1 U530 ( .A(n84), .B(n50), .ZN(product[11]) );
  NAND2_X1 U531 ( .A1(n127), .A2(n83), .ZN(n50) );
  NAND2_X1 U532 ( .A1(n152), .A2(n163), .ZN(n69) );
  NAND2_X1 U533 ( .A1(n561), .A2(n95), .ZN(n53) );
  OAI21_X1 U534 ( .B1(n113), .B2(n115), .A(n114), .ZN(n112) );
  NAND2_X1 U535 ( .A1(n131), .A2(n98), .ZN(n54) );
  INV_X1 U536 ( .A(n541), .ZN(n131) );
  AOI21_X1 U537 ( .B1(n564), .B2(n112), .A(n544), .ZN(n107) );
  NOR2_X1 U538 ( .A1(n176), .A2(n185), .ZN(n78) );
  AOI21_X1 U539 ( .B1(n562), .B2(n120), .A(n117), .ZN(n115) );
  INV_X1 U540 ( .A(n119), .ZN(n117) );
  NOR2_X1 U541 ( .A1(n196), .A2(n203), .ZN(n85) );
  INV_X1 U542 ( .A(n122), .ZN(n120) );
  XNOR2_X1 U543 ( .A(n57), .B(n112), .ZN(product[4]) );
  NAND2_X1 U544 ( .A1(n564), .A2(n111), .ZN(n57) );
  NAND2_X1 U545 ( .A1(n164), .A2(n175), .ZN(n76) );
  OR2_X1 U546 ( .A1(n212), .A2(n217), .ZN(n561) );
  NAND2_X1 U547 ( .A1(n176), .A2(n185), .ZN(n79) );
  NAND2_X1 U548 ( .A1(n212), .A2(n217), .ZN(n95) );
  INV_X1 U549 ( .A(n113), .ZN(n135) );
  NAND2_X1 U550 ( .A1(n204), .A2(n211), .ZN(n90) );
  NAND2_X1 U551 ( .A1(n186), .A2(n195), .ZN(n83) );
  NAND2_X1 U552 ( .A1(n196), .A2(n203), .ZN(n86) );
  XNOR2_X1 U553 ( .A(n59), .B(n120), .ZN(product[2]) );
  NAND2_X1 U554 ( .A1(n562), .A2(n119), .ZN(n59) );
  XNOR2_X1 U555 ( .A(n498), .B(n55), .ZN(product[6]) );
  NAND2_X1 U556 ( .A1(n543), .A2(n103), .ZN(n55) );
  NAND2_X1 U557 ( .A1(n490), .A2(n106), .ZN(n56) );
  NOR2_X1 U558 ( .A1(n234), .A2(n257), .ZN(n113) );
  XNOR2_X1 U559 ( .A(n63), .B(n46), .ZN(product[15]) );
  NAND2_X1 U560 ( .A1(n563), .A2(n62), .ZN(n46) );
  OR2_X1 U561 ( .A1(n328), .A2(n314), .ZN(n562) );
  OR2_X1 U562 ( .A1(n151), .A2(n139), .ZN(n563) );
  NAND2_X1 U563 ( .A1(n328), .A2(n314), .ZN(n119) );
  NOR2_X1 U564 ( .A1(n218), .A2(n223), .ZN(n97) );
  OR2_X1 U565 ( .A1(n232), .A2(n233), .ZN(n564) );
  NAND2_X1 U566 ( .A1(n218), .A2(n223), .ZN(n98) );
  INV_X1 U567 ( .A(n37), .ZN(n237) );
  NAND2_X1 U568 ( .A1(n545), .A2(n227), .ZN(n103) );
  OR2_X1 U569 ( .A1(n224), .A2(n227), .ZN(n565) );
  NAND2_X1 U570 ( .A1(n228), .A2(n231), .ZN(n106) );
  INV_X1 U571 ( .A(n41), .ZN(n235) );
  AND2_X1 U572 ( .A1(n494), .A2(n122), .ZN(product[1]) );
  OAI22_X1 U573 ( .A1(n546), .A2(n407), .B1(n406), .B2(n574), .ZN(n328) );
  XNOR2_X1 U574 ( .A(n590), .B(a[14]), .ZN(n41) );
  OR2_X1 U575 ( .A1(n572), .A2(n528), .ZN(n392) );
  OAI22_X1 U576 ( .A1(n547), .A2(n406), .B1(n405), .B2(n574), .ZN(n327) );
  OAI22_X1 U577 ( .A1(n547), .A2(n405), .B1(n404), .B2(n574), .ZN(n326) );
  AND2_X1 U578 ( .A1(n573), .A2(n245), .ZN(n300) );
  AND2_X1 U579 ( .A1(n573), .A2(n549), .ZN(n278) );
  OAI22_X1 U580 ( .A1(n547), .A2(n401), .B1(n400), .B2(n574), .ZN(n322) );
  OAI22_X1 U581 ( .A1(n6), .A2(n403), .B1(n402), .B2(n574), .ZN(n324) );
  AND2_X1 U582 ( .A1(n573), .A2(n522), .ZN(n288) );
  OAI22_X1 U583 ( .A1(n546), .A2(n397), .B1(n396), .B2(n574), .ZN(n318) );
  AND2_X1 U584 ( .A1(n573), .A2(n237), .ZN(n264) );
  OAI22_X1 U585 ( .A1(n547), .A2(n400), .B1(n399), .B2(n574), .ZN(n321) );
  XNOR2_X1 U586 ( .A(n586), .B(n572), .ZN(n352) );
  OAI22_X1 U587 ( .A1(n546), .A2(n408), .B1(n407), .B2(n574), .ZN(n329) );
  OAI22_X1 U588 ( .A1(n546), .A2(n396), .B1(n395), .B2(n574), .ZN(n317) );
  OAI22_X1 U589 ( .A1(n39), .A2(n591), .B1(n337), .B2(n532), .ZN(n252) );
  OR2_X1 U590 ( .A1(n572), .A2(n591), .ZN(n337) );
  OAI22_X1 U591 ( .A1(n42), .A2(n593), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U592 ( .A1(n572), .A2(n593), .ZN(n332) );
  OAI22_X1 U593 ( .A1(n6), .A2(n404), .B1(n403), .B2(n574), .ZN(n325) );
  OAI22_X1 U594 ( .A1(n547), .A2(n398), .B1(n397), .B2(n574), .ZN(n319) );
  XNOR2_X1 U595 ( .A(n529), .B(n572), .ZN(n343) );
  XNOR2_X1 U596 ( .A(n155), .B(n567), .ZN(n139) );
  XNOR2_X1 U597 ( .A(n153), .B(n141), .ZN(n567) );
  XNOR2_X1 U598 ( .A(n157), .B(n568), .ZN(n141) );
  XNOR2_X1 U599 ( .A(n145), .B(n143), .ZN(n568) );
  XOR2_X1 U600 ( .A(n315), .B(n261), .Z(n150) );
  OAI22_X1 U601 ( .A1(n546), .A2(n394), .B1(n393), .B2(n574), .ZN(n315) );
  XNOR2_X1 U602 ( .A(n582), .B(n572), .ZN(n376) );
  XNOR2_X1 U603 ( .A(n590), .B(n572), .ZN(n336) );
  AND2_X1 U604 ( .A1(n573), .A2(n247), .ZN(n314) );
  NAND2_X1 U605 ( .A1(n427), .A2(n37), .ZN(n39) );
  XOR2_X1 U606 ( .A(n590), .B(a[12]), .Z(n427) );
  OAI22_X1 U607 ( .A1(n39), .A2(n336), .B1(n532), .B2(n335), .ZN(n263) );
  AND2_X1 U608 ( .A1(n573), .A2(n235), .ZN(n260) );
  OAI22_X1 U609 ( .A1(n547), .A2(n395), .B1(n394), .B2(n574), .ZN(n316) );
  OAI22_X1 U610 ( .A1(n39), .A2(n335), .B1(n532), .B2(n334), .ZN(n262) );
  AND2_X1 U611 ( .A1(n573), .A2(n239), .ZN(n270) );
  OAI22_X1 U612 ( .A1(n546), .A2(n399), .B1(n398), .B2(n574), .ZN(n320) );
  INV_X1 U613 ( .A(n25), .ZN(n587) );
  NAND2_X1 U614 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U615 ( .A(n592), .B(a[14]), .Z(n426) );
  INV_X1 U616 ( .A(n7), .ZN(n580) );
  OAI22_X1 U617 ( .A1(n547), .A2(n402), .B1(n401), .B2(n574), .ZN(n323) );
  AND2_X1 U618 ( .A1(n573), .A2(n249), .ZN(product[0]) );
  OR2_X1 U619 ( .A1(n572), .A2(n589), .ZN(n344) );
  OR2_X1 U620 ( .A1(n572), .A2(n518), .ZN(n364) );
  OR2_X1 U621 ( .A1(n572), .A2(n587), .ZN(n353) );
  OR2_X1 U622 ( .A1(n572), .A2(n495), .ZN(n377) );
  OAI22_X1 U623 ( .A1(n39), .A2(n334), .B1(n532), .B2(n333), .ZN(n261) );
  XNOR2_X1 U624 ( .A(n590), .B(n422), .ZN(n333) );
  XNOR2_X1 U625 ( .A(n582), .B(b[11]), .ZN(n365) );
  XNOR2_X1 U626 ( .A(n590), .B(n424), .ZN(n335) );
  XNOR2_X1 U627 ( .A(n590), .B(n423), .ZN(n334) );
  OAI22_X1 U628 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U629 ( .A(n592), .B(n424), .ZN(n330) );
  XNOR2_X1 U630 ( .A(n592), .B(n572), .ZN(n331) );
  XNOR2_X1 U631 ( .A(n570), .B(b[13]), .ZN(n395) );
  XNOR2_X1 U632 ( .A(n570), .B(b[11]), .ZN(n397) );
  XNOR2_X1 U633 ( .A(n570), .B(b[14]), .ZN(n394) );
  XNOR2_X1 U634 ( .A(n557), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U635 ( .A(n586), .B(n418), .ZN(n345) );
  XNOR2_X1 U636 ( .A(n529), .B(n420), .ZN(n338) );
  XNOR2_X1 U637 ( .A(n579), .B(b[13]), .ZN(n378) );
  XNOR2_X1 U638 ( .A(n588), .B(n424), .ZN(n342) );
  XNOR2_X1 U639 ( .A(n529), .B(n423), .ZN(n341) );
  XNOR2_X1 U640 ( .A(n529), .B(n422), .ZN(n340) );
  XNOR2_X1 U641 ( .A(n529), .B(n421), .ZN(n339) );
  XNOR2_X1 U642 ( .A(n579), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U643 ( .A(n578), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U644 ( .A(n579), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U645 ( .A(n579), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U646 ( .A(n579), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U647 ( .A(n579), .B(n419), .ZN(n385) );
  XNOR2_X1 U648 ( .A(n579), .B(n418), .ZN(n384) );
  XNOR2_X1 U649 ( .A(n586), .B(n424), .ZN(n351) );
  XNOR2_X1 U650 ( .A(n582), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U651 ( .A(n582), .B(n418), .ZN(n369) );
  XNOR2_X1 U652 ( .A(n582), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U653 ( .A(n582), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U654 ( .A(n586), .B(n422), .ZN(n349) );
  XNOR2_X1 U655 ( .A(n586), .B(n423), .ZN(n350) );
  XNOR2_X1 U656 ( .A(n586), .B(n421), .ZN(n348) );
  XNOR2_X1 U657 ( .A(n586), .B(n420), .ZN(n347) );
  XNOR2_X1 U658 ( .A(n586), .B(n419), .ZN(n346) );
  XNOR2_X1 U659 ( .A(n557), .B(b[15]), .ZN(n393) );
  BUF_X1 U660 ( .A(n43), .Z(n573) );
  OAI22_X1 U661 ( .A1(n539), .A2(n339), .B1(n338), .B2(n521), .ZN(n265) );
  OAI22_X1 U662 ( .A1(n34), .A2(n340), .B1(n339), .B2(n521), .ZN(n266) );
  INV_X1 U663 ( .A(n32), .ZN(n239) );
  OAI22_X1 U664 ( .A1(n539), .A2(n342), .B1(n341), .B2(n521), .ZN(n268) );
  OAI22_X1 U665 ( .A1(n34), .A2(n341), .B1(n340), .B2(n521), .ZN(n267) );
  OAI22_X1 U666 ( .A1(n539), .A2(n343), .B1(n342), .B2(n521), .ZN(n269) );
  OAI22_X1 U667 ( .A1(n34), .A2(n589), .B1(n344), .B2(n32), .ZN(n253) );
  NAND2_X1 U668 ( .A1(n428), .A2(n32), .ZN(n34) );
  INV_X1 U669 ( .A(n249), .ZN(n574) );
  INV_X1 U670 ( .A(n577), .ZN(n575) );
  OAI22_X1 U671 ( .A1(n546), .A2(n527), .B1(n409), .B2(n574), .ZN(n258) );
  OR2_X1 U672 ( .A1(n572), .A2(n527), .ZN(n409) );
  INV_X1 U673 ( .A(n1), .ZN(n577) );
  NOR2_X1 U674 ( .A1(n204), .A2(n211), .ZN(n89) );
  OAI22_X1 U675 ( .A1(n29), .A2(n350), .B1(n349), .B2(n27), .ZN(n275) );
  OAI22_X1 U676 ( .A1(n29), .A2(n346), .B1(n345), .B2(n27), .ZN(n271) );
  OAI22_X1 U677 ( .A1(n29), .A2(n351), .B1(n350), .B2(n27), .ZN(n276) );
  OAI22_X1 U678 ( .A1(n29), .A2(n347), .B1(n346), .B2(n27), .ZN(n272) );
  OAI22_X1 U679 ( .A1(n29), .A2(n587), .B1(n353), .B2(n27), .ZN(n254) );
  OAI22_X1 U680 ( .A1(n29), .A2(n349), .B1(n348), .B2(n27), .ZN(n274) );
  OAI22_X1 U681 ( .A1(n29), .A2(n348), .B1(n347), .B2(n27), .ZN(n273) );
  XNOR2_X1 U682 ( .A(n525), .B(n422), .ZN(n360) );
  OAI22_X1 U683 ( .A1(n29), .A2(n352), .B1(n351), .B2(n27), .ZN(n277) );
  XNOR2_X1 U684 ( .A(n525), .B(n419), .ZN(n357) );
  XNOR2_X1 U685 ( .A(n525), .B(n423), .ZN(n361) );
  XNOR2_X1 U686 ( .A(n525), .B(n418), .ZN(n356) );
  XNOR2_X1 U687 ( .A(n525), .B(b[9]), .ZN(n354) );
  XNOR2_X1 U688 ( .A(n525), .B(b[8]), .ZN(n355) );
  XNOR2_X1 U689 ( .A(n525), .B(n572), .ZN(n363) );
  XNOR2_X1 U690 ( .A(n526), .B(n420), .ZN(n358) );
  XNOR2_X1 U691 ( .A(n526), .B(n421), .ZN(n359) );
  XNOR2_X1 U692 ( .A(n526), .B(n424), .ZN(n362) );
  XNOR2_X1 U693 ( .A(n540), .B(n571), .ZN(product[12]) );
  AND2_X1 U694 ( .A1(n531), .A2(n79), .ZN(n571) );
  NOR2_X1 U695 ( .A1(n536), .A2(n85), .ZN(n80) );
  INV_X1 U696 ( .A(n536), .ZN(n127) );
  OAI21_X1 U697 ( .B1(n86), .B2(n82), .A(n83), .ZN(n81) );
  XNOR2_X1 U698 ( .A(n70), .B(n47), .ZN(product[14]) );
  XNOR2_X1 U699 ( .A(n77), .B(n48), .ZN(product[13]) );
  OAI21_X1 U700 ( .B1(n107), .B2(n105), .A(n106), .ZN(n104) );
  NOR2_X1 U701 ( .A1(n228), .A2(n231), .ZN(n105) );
  XNOR2_X1 U702 ( .A(n581), .B(n424), .ZN(n375) );
  XNOR2_X1 U703 ( .A(n581), .B(n423), .ZN(n374) );
  XNOR2_X1 U704 ( .A(n581), .B(n422), .ZN(n373) );
  XNOR2_X1 U705 ( .A(n581), .B(n419), .ZN(n370) );
  XNOR2_X1 U706 ( .A(n581), .B(n420), .ZN(n371) );
  XNOR2_X1 U707 ( .A(n581), .B(n421), .ZN(n372) );
  NAND2_X1 U708 ( .A1(n135), .A2(n114), .ZN(n58) );
  OAI21_X1 U709 ( .B1(n87), .B2(n523), .A(n496), .ZN(n84) );
  INV_X1 U710 ( .A(n88), .ZN(n87) );
  OAI21_X1 U711 ( .B1(n91), .B2(n89), .A(n90), .ZN(n88) );
  NAND2_X1 U712 ( .A1(n151), .A2(n139), .ZN(n62) );
  OAI22_X1 U713 ( .A1(n23), .A2(n358), .B1(n357), .B2(n21), .ZN(n282) );
  OAI22_X1 U714 ( .A1(n520), .A2(n356), .B1(n355), .B2(n21), .ZN(n280) );
  OAI22_X1 U715 ( .A1(n520), .A2(n362), .B1(n361), .B2(n21), .ZN(n286) );
  OAI22_X1 U716 ( .A1(n23), .A2(n357), .B1(n356), .B2(n21), .ZN(n281) );
  OAI22_X1 U717 ( .A1(n23), .A2(n360), .B1(n359), .B2(n21), .ZN(n284) );
  OAI22_X1 U718 ( .A1(n520), .A2(n361), .B1(n360), .B2(n21), .ZN(n285) );
  OAI22_X1 U719 ( .A1(n520), .A2(n518), .B1(n364), .B2(n21), .ZN(n255) );
  OAI22_X1 U720 ( .A1(n520), .A2(n363), .B1(n362), .B2(n21), .ZN(n287) );
  OAI22_X1 U721 ( .A1(n359), .A2(n23), .B1(n358), .B2(n21), .ZN(n283) );
  OAI22_X1 U722 ( .A1(n23), .A2(n355), .B1(n354), .B2(n21), .ZN(n279) );
  OAI21_X1 U723 ( .B1(n99), .B2(n97), .A(n98), .ZN(n96) );
  XNOR2_X1 U724 ( .A(n538), .B(n53), .ZN(product[8]) );
  OAI22_X1 U725 ( .A1(n534), .A2(n370), .B1(n369), .B2(n505), .ZN(n293) );
  OAI22_X1 U726 ( .A1(n511), .A2(n367), .B1(n366), .B2(n569), .ZN(n290) );
  OAI22_X1 U727 ( .A1(n501), .A2(n368), .B1(n367), .B2(n569), .ZN(n291) );
  OAI22_X1 U728 ( .A1(n500), .A2(n371), .B1(n370), .B2(n569), .ZN(n294) );
  OAI22_X1 U729 ( .A1(n500), .A2(n369), .B1(n368), .B2(n569), .ZN(n292) );
  OAI22_X1 U730 ( .A1(n501), .A2(n372), .B1(n371), .B2(n569), .ZN(n295) );
  OAI22_X1 U731 ( .A1(n534), .A2(n375), .B1(n374), .B2(n505), .ZN(n298) );
  OAI22_X1 U732 ( .A1(n500), .A2(n376), .B1(n375), .B2(n569), .ZN(n299) );
  OAI22_X1 U733 ( .A1(n500), .A2(n495), .B1(n377), .B2(n569), .ZN(n256) );
  OAI22_X1 U734 ( .A1(n501), .A2(n373), .B1(n372), .B2(n569), .ZN(n296) );
  OAI22_X1 U735 ( .A1(n501), .A2(n366), .B1(n365), .B2(n569), .ZN(n289) );
  OAI22_X1 U736 ( .A1(n374), .A2(n499), .B1(n373), .B2(n569), .ZN(n297) );
  INV_X1 U737 ( .A(n569), .ZN(n245) );
  XNOR2_X1 U738 ( .A(n579), .B(n572), .ZN(n391) );
  XNOR2_X1 U739 ( .A(n579), .B(n420), .ZN(n386) );
  XNOR2_X1 U740 ( .A(n579), .B(n424), .ZN(n390) );
  XNOR2_X1 U741 ( .A(n578), .B(n422), .ZN(n388) );
  XNOR2_X1 U742 ( .A(n578), .B(n423), .ZN(n389) );
  XNOR2_X1 U743 ( .A(n578), .B(n421), .ZN(n387) );
  XOR2_X1 U744 ( .A(n555), .B(n54), .Z(product[7]) );
  AOI21_X1 U745 ( .B1(n104), .B2(n565), .A(n556), .ZN(n99) );
  OAI21_X1 U746 ( .B1(n64), .B2(n506), .A(n65), .ZN(n63) );
  OAI21_X1 U747 ( .B1(n512), .B2(n78), .A(n79), .ZN(n77) );
  OAI21_X1 U748 ( .B1(n512), .B2(n71), .A(n72), .ZN(n70) );
  XNOR2_X1 U749 ( .A(n570), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U750 ( .A(n576), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U751 ( .A(n570), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U752 ( .A(n519), .B(n418), .ZN(n401) );
  XNOR2_X1 U753 ( .A(n557), .B(n572), .ZN(n408) );
  XNOR2_X1 U754 ( .A(n570), .B(n421), .ZN(n404) );
  XNOR2_X1 U755 ( .A(n570), .B(n422), .ZN(n405) );
  XNOR2_X1 U756 ( .A(n576), .B(n420), .ZN(n403) );
  XNOR2_X1 U757 ( .A(n570), .B(n419), .ZN(n402) );
  XNOR2_X1 U758 ( .A(n557), .B(n424), .ZN(n407) );
  XNOR2_X1 U759 ( .A(n570), .B(n423), .ZN(n406) );
  XOR2_X1 U760 ( .A(n56), .B(n530), .Z(product[5]) );
  XOR2_X1 U761 ( .A(n58), .B(n115), .Z(product[3]) );
  NAND2_X1 U762 ( .A1(n329), .A2(n258), .ZN(n122) );
  OAI22_X1 U763 ( .A1(n514), .A2(n379), .B1(n378), .B2(n558), .ZN(n301) );
  OAI22_X1 U764 ( .A1(n514), .A2(n380), .B1(n379), .B2(n558), .ZN(n302) );
  OAI22_X1 U765 ( .A1(n504), .A2(n385), .B1(n384), .B2(n516), .ZN(n307) );
  OAI22_X1 U766 ( .A1(n552), .A2(n382), .B1(n381), .B2(n558), .ZN(n304) );
  OAI22_X1 U767 ( .A1(n551), .A2(n381), .B1(n380), .B2(n558), .ZN(n303) );
  NAND2_X1 U768 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U769 ( .A1(n383), .A2(n552), .B1(n382), .B2(n497), .ZN(n305) );
  OAI22_X1 U770 ( .A1(n551), .A2(n384), .B1(n383), .B2(n558), .ZN(n306) );
  OAI22_X1 U771 ( .A1(n551), .A2(n386), .B1(n385), .B2(n558), .ZN(n308) );
  OAI22_X1 U772 ( .A1(n504), .A2(n387), .B1(n386), .B2(n558), .ZN(n309) );
  OAI22_X1 U773 ( .A1(n504), .A2(n528), .B1(n392), .B2(n516), .ZN(n257) );
  OAI22_X1 U774 ( .A1(n551), .A2(n389), .B1(n388), .B2(n535), .ZN(n311) );
  OAI22_X1 U775 ( .A1(n12), .A2(n388), .B1(n387), .B2(n535), .ZN(n310) );
  OAI22_X1 U776 ( .A1(n551), .A2(n390), .B1(n389), .B2(n558), .ZN(n312) );
  INV_X1 U777 ( .A(n558), .ZN(n247) );
  OAI22_X1 U778 ( .A1(n12), .A2(n391), .B1(n390), .B2(n558), .ZN(n313) );
  INV_X1 U779 ( .A(n583), .ZN(n582) );
  INV_X1 U780 ( .A(n31), .ZN(n589) );
  INV_X1 U781 ( .A(n36), .ZN(n591) );
  INV_X1 U782 ( .A(n593), .ZN(n592) );
  INV_X1 U783 ( .A(n40), .ZN(n593) );
  XOR2_X1 U784 ( .A(n259), .B(n251), .Z(n148) );
  XOR2_X1 U785 ( .A(n289), .B(n279), .Z(n146) );
  XOR2_X1 U786 ( .A(n159), .B(n150), .Z(n142) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_6_DW01_add_2 ( A, B, CI, SUM, 
        CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n18, n19,
         n20, n21, n23, n25, n26, n27, n28, n30, n34, n35, n36, n37, n38, n39,
         n40, n42, n43, n44, n48, n49, n51, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n69, n71, n72, n73, n74, n75,
         n77, n79, n80, n81, n82, n83, n85, n87, n88, n90, n93, n94, n98, n99,
         n100, n102, n104, n161, n162, n163, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182;

  INV_X1 U126 ( .A(n93), .ZN(n161) );
  XNOR2_X1 U127 ( .A(n171), .B(n162), .ZN(SUM[13]) );
  AND2_X1 U128 ( .A1(n93), .A2(n28), .ZN(n162) );
  BUF_X1 U129 ( .A(n40), .Z(n163) );
  AND2_X1 U130 ( .A1(n175), .A2(n90), .ZN(SUM[0]) );
  OR2_X1 U131 ( .A1(A[15]), .A2(B[15]), .ZN(n165) );
  AOI21_X1 U132 ( .B1(n56), .B2(n64), .A(n57), .ZN(n166) );
  OR2_X1 U133 ( .A1(A[11]), .A2(B[11]), .ZN(n167) );
  XNOR2_X1 U134 ( .A(n170), .B(n168), .ZN(SUM[11]) );
  AND2_X1 U135 ( .A1(n167), .A2(n40), .ZN(n168) );
  AOI21_X2 U136 ( .B1(n42), .B2(n34), .A(n35), .ZN(n171) );
  CLKBUF_X1 U137 ( .A(n28), .Z(n169) );
  INV_X1 U138 ( .A(n42), .ZN(n170) );
  NOR2_X1 U139 ( .A1(A[8]), .A2(B[8]), .ZN(n172) );
  INV_X1 U140 ( .A(n167), .ZN(n173) );
  NOR2_X1 U141 ( .A1(A[12]), .A2(B[12]), .ZN(n174) );
  NOR2_X1 U142 ( .A1(A[12]), .A2(B[12]), .ZN(n36) );
  OR2_X2 U143 ( .A1(A[10]), .A2(B[10]), .ZN(n181) );
  OR2_X1 U144 ( .A1(A[0]), .A2(B[0]), .ZN(n175) );
  INV_X1 U145 ( .A(n64), .ZN(n63) );
  INV_X1 U146 ( .A(n166), .ZN(n54) );
  AOI21_X1 U147 ( .B1(n56), .B2(n64), .A(n57), .ZN(n55) );
  AOI21_X1 U148 ( .B1(n176), .B2(n80), .A(n77), .ZN(n75) );
  INV_X1 U149 ( .A(n79), .ZN(n77) );
  OAI21_X1 U150 ( .B1(n67), .B2(n65), .A(n66), .ZN(n64) );
  OAI21_X1 U151 ( .B1(n75), .B2(n73), .A(n74), .ZN(n72) );
  OAI21_X1 U152 ( .B1(n83), .B2(n81), .A(n82), .ZN(n80) );
  AOI21_X1 U153 ( .B1(n177), .B2(n72), .A(n69), .ZN(n67) );
  INV_X1 U154 ( .A(n71), .ZN(n69) );
  AOI21_X1 U155 ( .B1(n54), .B2(n178), .A(n51), .ZN(n49) );
  NAND2_X1 U156 ( .A1(n98), .A2(n59), .ZN(n8) );
  INV_X1 U157 ( .A(n90), .ZN(n88) );
  OAI21_X1 U158 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  INV_X1 U159 ( .A(n27), .ZN(n93) );
  AOI21_X1 U160 ( .B1(n179), .B2(n88), .A(n85), .ZN(n83) );
  INV_X1 U161 ( .A(n87), .ZN(n85) );
  NAND2_X1 U162 ( .A1(n102), .A2(n74), .ZN(n12) );
  INV_X1 U163 ( .A(n73), .ZN(n102) );
  NAND2_X1 U164 ( .A1(n100), .A2(n66), .ZN(n10) );
  INV_X1 U165 ( .A(n65), .ZN(n100) );
  NAND2_X1 U166 ( .A1(n177), .A2(n71), .ZN(n11) );
  NAND2_X1 U167 ( .A1(n178), .A2(n53), .ZN(n7) );
  NAND2_X1 U168 ( .A1(n99), .A2(n62), .ZN(n9) );
  INV_X1 U169 ( .A(n61), .ZN(n99) );
  NAND2_X1 U170 ( .A1(n104), .A2(n82), .ZN(n14) );
  INV_X1 U171 ( .A(n81), .ZN(n104) );
  NAND2_X1 U172 ( .A1(n176), .A2(n79), .ZN(n13) );
  NAND2_X1 U173 ( .A1(n179), .A2(n87), .ZN(n15) );
  INV_X1 U174 ( .A(n25), .ZN(n23) );
  XOR2_X1 U175 ( .A(n49), .B(n6), .Z(SUM[10]) );
  XNOR2_X1 U176 ( .A(n54), .B(n7), .ZN(SUM[9]) );
  XOR2_X1 U177 ( .A(n63), .B(n9), .Z(SUM[7]) );
  XNOR2_X1 U178 ( .A(n13), .B(n80), .ZN(SUM[3]) );
  XNOR2_X1 U179 ( .A(n15), .B(n88), .ZN(SUM[1]) );
  OR2_X1 U180 ( .A1(A[3]), .A2(B[3]), .ZN(n176) );
  OR2_X1 U181 ( .A1(A[5]), .A2(B[5]), .ZN(n177) );
  NOR2_X1 U182 ( .A1(A[7]), .A2(B[7]), .ZN(n61) );
  NOR2_X1 U183 ( .A1(A[11]), .A2(B[11]), .ZN(n39) );
  OR2_X1 U184 ( .A1(A[9]), .A2(B[9]), .ZN(n178) );
  NOR2_X1 U185 ( .A1(A[2]), .A2(B[2]), .ZN(n81) );
  NOR2_X1 U186 ( .A1(A[4]), .A2(B[4]), .ZN(n73) );
  NAND2_X1 U187 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  NAND2_X1 U188 ( .A1(A[11]), .A2(B[11]), .ZN(n40) );
  OR2_X1 U189 ( .A1(A[1]), .A2(B[1]), .ZN(n179) );
  OR2_X1 U190 ( .A1(A[14]), .A2(B[14]), .ZN(n180) );
  NOR2_X1 U191 ( .A1(A[6]), .A2(B[6]), .ZN(n65) );
  NOR2_X1 U192 ( .A1(A[8]), .A2(B[8]), .ZN(n58) );
  XNOR2_X1 U193 ( .A(n60), .B(n8), .ZN(SUM[8]) );
  XNOR2_X1 U194 ( .A(n11), .B(n72), .ZN(SUM[5]) );
  NAND2_X1 U195 ( .A1(A[7]), .A2(B[7]), .ZN(n62) );
  NAND2_X1 U196 ( .A1(A[2]), .A2(B[2]), .ZN(n82) );
  NAND2_X1 U197 ( .A1(A[4]), .A2(B[4]), .ZN(n74) );
  NAND2_X1 U198 ( .A1(A[1]), .A2(B[1]), .ZN(n87) );
  NAND2_X1 U199 ( .A1(A[0]), .A2(B[0]), .ZN(n90) );
  NAND2_X1 U200 ( .A1(A[6]), .A2(B[6]), .ZN(n66) );
  NAND2_X1 U201 ( .A1(A[8]), .A2(B[8]), .ZN(n59) );
  NAND2_X1 U202 ( .A1(A[3]), .A2(B[3]), .ZN(n79) );
  XOR2_X1 U203 ( .A(n12), .B(n75), .Z(SUM[4]) );
  XOR2_X1 U204 ( .A(n14), .B(n83), .Z(SUM[2]) );
  NAND2_X1 U205 ( .A1(n165), .A2(n18), .ZN(n1) );
  NAND2_X1 U206 ( .A1(A[9]), .A2(B[9]), .ZN(n53) );
  INV_X1 U207 ( .A(n182), .ZN(n48) );
  NAND2_X1 U208 ( .A1(A[15]), .A2(B[15]), .ZN(n18) );
  NAND2_X1 U209 ( .A1(A[12]), .A2(B[12]), .ZN(n37) );
  NAND2_X1 U210 ( .A1(n94), .A2(n37), .ZN(n4) );
  INV_X1 U211 ( .A(n174), .ZN(n94) );
  AND2_X1 U212 ( .A1(A[10]), .A2(B[10]), .ZN(n182) );
  INV_X1 U213 ( .A(n53), .ZN(n51) );
  XOR2_X1 U214 ( .A(n10), .B(n67), .Z(SUM[6]) );
  NAND2_X1 U215 ( .A1(A[5]), .A2(B[5]), .ZN(n71) );
  NOR2_X1 U216 ( .A1(A[13]), .A2(B[13]), .ZN(n27) );
  XNOR2_X1 U217 ( .A(n38), .B(n4), .ZN(SUM[12]) );
  INV_X1 U218 ( .A(n172), .ZN(n98) );
  NOR2_X1 U219 ( .A1(n172), .A2(n61), .ZN(n56) );
  OAI21_X1 U220 ( .B1(n58), .B2(n62), .A(n59), .ZN(n57) );
  INV_X1 U221 ( .A(n28), .ZN(n30) );
  AOI21_X1 U222 ( .B1(n180), .B2(n30), .A(n23), .ZN(n21) );
  NAND2_X1 U223 ( .A1(n180), .A2(n93), .ZN(n20) );
  NAND2_X1 U224 ( .A1(n180), .A2(n25), .ZN(n2) );
  NAND2_X1 U225 ( .A1(A[14]), .A2(B[14]), .ZN(n25) );
  OAI21_X1 U226 ( .B1(n36), .B2(n40), .A(n37), .ZN(n35) );
  OAI21_X1 U227 ( .B1(n170), .B2(n173), .A(n163), .ZN(n38) );
  NOR2_X1 U228 ( .A1(n174), .A2(n39), .ZN(n34) );
  OAI21_X1 U229 ( .B1(n43), .B2(n55), .A(n44), .ZN(n42) );
  AOI21_X1 U230 ( .B1(n181), .B2(n51), .A(n182), .ZN(n44) );
  XNOR2_X1 U231 ( .A(n19), .B(n1), .ZN(SUM[15]) );
  NAND2_X1 U232 ( .A1(n181), .A2(n48), .ZN(n6) );
  NAND2_X1 U233 ( .A1(n181), .A2(n178), .ZN(n43) );
  XNOR2_X1 U234 ( .A(n26), .B(n2), .ZN(SUM[14]) );
  OAI21_X1 U235 ( .B1(n171), .B2(n161), .A(n169), .ZN(n26) );
  OAI21_X1 U236 ( .B1(n171), .B2(n20), .A(n21), .ZN(n19) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_6 ( clk, clear_acc, 
        data_out_x, data_out, data_out_w, data_out_b, wr_en_y, m_valid, 
        m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [3:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N27, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, n1, n2, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n87, n104, n113, n114, n115, n116, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n21), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n225), .CK(clk), .Q(n26) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n226), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n227), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n228), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n229), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n230), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n231), .CK(clk), .Q(n34) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n232), .CK(clk), .Q(n35) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n233), .CK(clk), .Q(n36) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n234), .CK(clk), .Q(n37) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n235), .CK(clk), .Q(n38) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n236), .CK(clk), .Q(n39) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n237), .CK(clk), .Q(n40) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n238), .CK(clk), .Q(n41) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n239), .CK(clk), .Q(n42) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n240), .CK(clk), .Q(n44) );
  DFF_X1 \f_reg[7]  ( .D(n83), .CK(clk), .Q(f[7]), .QN(n217) );
  DFF_X1 \f_reg[8]  ( .D(n82), .CK(clk), .Q(f[8]), .QN(n218) );
  DFF_X1 \f_reg[9]  ( .D(n81), .CK(clk), .Q(f[9]), .QN(n219) );
  DFF_X1 \f_reg[10]  ( .D(n80), .CK(clk), .Q(n53), .QN(n220) );
  DFF_X1 \f_reg[11]  ( .D(n79), .CK(clk), .Q(n51), .QN(n221) );
  DFF_X1 \f_reg[12]  ( .D(n1), .CK(clk), .Q(n50), .QN(n222) );
  DFF_X1 \f_reg[13]  ( .D(n16), .CK(clk), .Q(n49), .QN(n223) );
  DFF_X1 \f_reg[14]  ( .D(n7), .CK(clk), .Q(n48), .QN(n224) );
  DFF_X1 \f_reg[15]  ( .D(n6), .CK(clk), .Q(f[15]), .QN(n77) );
  DFF_X1 \data_out_reg[15]  ( .D(n116), .CK(clk), .Q(data_out[15]), .QN(n197)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n167), .CK(clk), .Q(data_out[14]), .QN(n196)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n168), .CK(clk), .Q(data_out[13]), .QN(n195)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n169), .CK(clk), .Q(data_out[12]), .QN(n194)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n170), .CK(clk), .Q(data_out[11]), .QN(n193)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n171), .CK(clk), .Q(data_out[10]), .QN(n192)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n172), .CK(clk), .Q(data_out[9]), .QN(n191) );
  DFF_X1 \data_out_reg[8]  ( .D(n173), .CK(clk), .Q(data_out[8]), .QN(n190) );
  DFF_X1 \data_out_reg[7]  ( .D(n174), .CK(clk), .Q(data_out[7]), .QN(n189) );
  DFF_X1 \data_out_reg[6]  ( .D(n175), .CK(clk), .Q(data_out[6]), .QN(n188) );
  DFF_X1 \data_out_reg[5]  ( .D(n176), .CK(clk), .Q(data_out[5]), .QN(n187) );
  DFF_X1 \data_out_reg[4]  ( .D(n177), .CK(clk), .Q(data_out[4]), .QN(n186) );
  DFF_X1 \data_out_reg[3]  ( .D(n178), .CK(clk), .Q(data_out[3]), .QN(n185) );
  DFF_X1 \data_out_reg[2]  ( .D(n179), .CK(clk), .Q(data_out[2]), .QN(n184) );
  DFF_X1 \data_out_reg[1]  ( .D(n180), .CK(clk), .Q(data_out[1]), .QN(n183) );
  DFF_X1 \data_out_reg[0]  ( .D(n181), .CK(clk), .Q(data_out[0]), .QN(n182) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_6_DW_mult_tc_1 mult_960 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_6_DW01_add_2 add_961 ( .A({n204, 
        n203, n202, n201, n200, n199, n213, n212, n211, n210, n209, n208, n207, 
        n206, n205, n198}), .B({f[15], n48, n49, n50, n51, n53, f[9:3], n61, 
        n63, n65}), .CI(1'b0), .SUM(adder) );
  DFF_X2 delay_reg ( .D(N27), .CK(clk), .Q(n14), .QN(n241) );
  DFF_X1 \f_reg[2]  ( .D(n113), .CK(clk), .Q(n61), .QN(n216) );
  DFF_X1 \f_reg[3]  ( .D(n104), .CK(clk), .Q(f[3]), .QN(n69) );
  DFF_X1 \f_reg[1]  ( .D(n114), .CK(clk), .Q(n63), .QN(n215) );
  DFF_X1 \f_reg[0]  ( .D(n115), .CK(clk), .Q(n65), .QN(n214) );
  DFF_X1 \f_reg[4]  ( .D(n87), .CK(clk), .Q(f[4]), .QN(n70) );
  DFF_X1 \f_reg[5]  ( .D(n85), .CK(clk), .Q(f[5]), .QN(n71) );
  DFF_X1 \f_reg[6]  ( .D(n84), .CK(clk), .Q(f[6]), .QN(n72) );
  AND2_X2 U3 ( .A1(n47), .A2(n22), .ZN(n15) );
  MUX2_X2 U4 ( .A(N41), .B(n29), .S(n14), .Z(n201) );
  MUX2_X1 U5 ( .A(N39), .B(n33), .S(n14), .Z(n199) );
  MUX2_X2 U6 ( .A(n32), .B(N40), .S(n241), .Z(n200) );
  MUX2_X2 U8 ( .A(N43), .B(n27), .S(n14), .Z(n203) );
  NAND3_X1 U9 ( .A1(n4), .A2(n2), .A3(n5), .ZN(n1) );
  NAND2_X1 U10 ( .A1(data_out_b[12]), .A2(n21), .ZN(n2) );
  NAND2_X1 U11 ( .A1(adder[12]), .A2(n15), .ZN(n4) );
  NAND2_X1 U12 ( .A1(n67), .A2(n50), .ZN(n5) );
  NAND3_X1 U13 ( .A1(n12), .A2(n11), .A3(n13), .ZN(n6) );
  NAND3_X1 U14 ( .A1(n9), .A2(n8), .A3(n10), .ZN(n7) );
  MUX2_X2 U15 ( .A(n35), .B(N37), .S(n241), .Z(n212) );
  NAND2_X1 U16 ( .A1(data_out_b[14]), .A2(n21), .ZN(n8) );
  NAND2_X1 U17 ( .A1(adder[14]), .A2(n15), .ZN(n9) );
  NAND2_X1 U18 ( .A1(n67), .A2(n48), .ZN(n10) );
  NAND2_X1 U19 ( .A1(data_out_b[15]), .A2(n21), .ZN(n11) );
  NAND2_X1 U20 ( .A1(adder[15]), .A2(n15), .ZN(n12) );
  NAND2_X1 U21 ( .A1(n67), .A2(f[15]), .ZN(n13) );
  INV_X2 U22 ( .A(n47), .ZN(n67) );
  INV_X1 U23 ( .A(clear_acc), .ZN(n22) );
  NAND2_X1 U24 ( .A1(n20), .A2(N27), .ZN(n243) );
  INV_X1 U25 ( .A(n25), .ZN(n43) );
  OAI22_X1 U26 ( .A1(n185), .A2(n243), .B1(n69), .B2(n242), .ZN(n178) );
  OAI22_X1 U27 ( .A1(n186), .A2(n243), .B1(n70), .B2(n242), .ZN(n177) );
  OAI22_X1 U28 ( .A1(n187), .A2(n243), .B1(n71), .B2(n242), .ZN(n176) );
  OAI22_X1 U29 ( .A1(n188), .A2(n243), .B1(n72), .B2(n242), .ZN(n175) );
  OAI22_X1 U30 ( .A1(n189), .A2(n243), .B1(n217), .B2(n242), .ZN(n174) );
  OAI22_X1 U31 ( .A1(n190), .A2(n243), .B1(n218), .B2(n242), .ZN(n173) );
  OAI22_X1 U32 ( .A1(n191), .A2(n243), .B1(n219), .B2(n242), .ZN(n172) );
  MUX2_X1 U33 ( .A(n40), .B(N32), .S(n241), .Z(n207) );
  MUX2_X1 U34 ( .A(n28), .B(N42), .S(n241), .Z(n202) );
  MUX2_X1 U35 ( .A(n26), .B(N44), .S(n241), .Z(n204) );
  NAND3_X1 U36 ( .A1(n18), .A2(n17), .A3(n19), .ZN(n16) );
  NAND2_X1 U37 ( .A1(data_out_b[13]), .A2(n21), .ZN(n17) );
  NAND2_X1 U38 ( .A1(adder[13]), .A2(n15), .ZN(n18) );
  NAND2_X1 U39 ( .A1(n67), .A2(n49), .ZN(n19) );
  INV_X1 U40 ( .A(n22), .ZN(n21) );
  INV_X1 U41 ( .A(wr_en_y), .ZN(n20) );
  AND2_X1 U42 ( .A1(sel[0]), .A2(sel[1]), .ZN(n24) );
  INV_X1 U43 ( .A(m_ready), .ZN(n23) );
  NAND2_X1 U44 ( .A1(m_valid), .A2(n23), .ZN(n45) );
  OAI211_X1 U45 ( .C1(sel[2]), .C2(n24), .A(sel[3]), .B(n45), .ZN(N27) );
  NAND2_X1 U46 ( .A1(clear_acc_delay), .A2(n241), .ZN(n25) );
  MUX2_X1 U47 ( .A(n26), .B(N44), .S(n43), .Z(n225) );
  MUX2_X1 U48 ( .A(n27), .B(N43), .S(n43), .Z(n226) );
  MUX2_X1 U49 ( .A(n28), .B(N42), .S(n43), .Z(n227) );
  MUX2_X1 U50 ( .A(n29), .B(N41), .S(n43), .Z(n228) );
  MUX2_X1 U51 ( .A(n32), .B(N40), .S(n43), .Z(n229) );
  MUX2_X1 U52 ( .A(n33), .B(N39), .S(n43), .Z(n230) );
  MUX2_X1 U53 ( .A(n34), .B(N38), .S(n43), .Z(n231) );
  MUX2_X1 U54 ( .A(n34), .B(N38), .S(n241), .Z(n213) );
  MUX2_X1 U55 ( .A(n35), .B(N37), .S(n43), .Z(n232) );
  MUX2_X1 U56 ( .A(n36), .B(N36), .S(n43), .Z(n233) );
  MUX2_X1 U57 ( .A(n36), .B(N36), .S(n241), .Z(n211) );
  MUX2_X1 U58 ( .A(n37), .B(N35), .S(n43), .Z(n234) );
  MUX2_X1 U59 ( .A(n37), .B(N35), .S(n241), .Z(n210) );
  MUX2_X1 U60 ( .A(n38), .B(N34), .S(n43), .Z(n235) );
  MUX2_X1 U61 ( .A(n38), .B(N34), .S(n241), .Z(n209) );
  MUX2_X1 U62 ( .A(n39), .B(N33), .S(n43), .Z(n236) );
  MUX2_X1 U63 ( .A(n39), .B(N33), .S(n241), .Z(n208) );
  MUX2_X1 U64 ( .A(n40), .B(N32), .S(n43), .Z(n237) );
  MUX2_X1 U65 ( .A(n41), .B(N31), .S(n43), .Z(n238) );
  MUX2_X1 U66 ( .A(n41), .B(N31), .S(n241), .Z(n206) );
  MUX2_X1 U67 ( .A(n42), .B(N30), .S(n43), .Z(n239) );
  MUX2_X1 U68 ( .A(n42), .B(N30), .S(n241), .Z(n205) );
  MUX2_X1 U69 ( .A(n44), .B(N29), .S(n43), .Z(n240) );
  MUX2_X1 U70 ( .A(n44), .B(N29), .S(n241), .Z(n198) );
  INV_X1 U71 ( .A(n45), .ZN(n46) );
  OAI21_X1 U72 ( .B1(n46), .B2(n14), .A(n22), .ZN(n47) );
  AOI222_X1 U73 ( .A1(data_out_b[11]), .A2(n21), .B1(adder[11]), .B2(n15), 
        .C1(n67), .C2(n51), .ZN(n52) );
  INV_X1 U74 ( .A(n52), .ZN(n79) );
  AOI222_X1 U75 ( .A1(data_out_b[10]), .A2(n21), .B1(adder[10]), .B2(n15), 
        .C1(n67), .C2(n53), .ZN(n54) );
  INV_X1 U76 ( .A(n54), .ZN(n80) );
  AOI222_X1 U77 ( .A1(data_out_b[8]), .A2(n21), .B1(adder[8]), .B2(n15), .C1(
        n67), .C2(f[8]), .ZN(n55) );
  INV_X1 U78 ( .A(n55), .ZN(n82) );
  AOI222_X1 U79 ( .A1(data_out_b[7]), .A2(n21), .B1(adder[7]), .B2(n15), .C1(
        n67), .C2(f[7]), .ZN(n56) );
  INV_X1 U80 ( .A(n56), .ZN(n83) );
  AOI222_X1 U81 ( .A1(data_out_b[6]), .A2(n21), .B1(adder[6]), .B2(n15), .C1(
        n67), .C2(f[6]), .ZN(n57) );
  INV_X1 U82 ( .A(n57), .ZN(n84) );
  AOI222_X1 U83 ( .A1(data_out_b[5]), .A2(n21), .B1(adder[5]), .B2(n15), .C1(
        n67), .C2(f[5]), .ZN(n58) );
  INV_X1 U84 ( .A(n58), .ZN(n85) );
  AOI222_X1 U85 ( .A1(data_out_b[4]), .A2(n21), .B1(adder[4]), .B2(n15), .C1(
        n67), .C2(f[4]), .ZN(n59) );
  INV_X1 U86 ( .A(n59), .ZN(n87) );
  AOI222_X1 U87 ( .A1(data_out_b[3]), .A2(n21), .B1(adder[3]), .B2(n15), .C1(
        n67), .C2(f[3]), .ZN(n60) );
  INV_X1 U88 ( .A(n60), .ZN(n104) );
  AOI222_X1 U89 ( .A1(data_out_b[2]), .A2(n21), .B1(adder[2]), .B2(n15), .C1(
        n67), .C2(n61), .ZN(n62) );
  INV_X1 U90 ( .A(n62), .ZN(n113) );
  AOI222_X1 U91 ( .A1(data_out_b[1]), .A2(n21), .B1(adder[1]), .B2(n15), .C1(
        n67), .C2(n63), .ZN(n64) );
  INV_X1 U92 ( .A(n64), .ZN(n114) );
  AOI222_X1 U93 ( .A1(data_out_b[0]), .A2(n21), .B1(adder[0]), .B2(n15), .C1(
        n67), .C2(n65), .ZN(n66) );
  INV_X1 U94 ( .A(n66), .ZN(n115) );
  AOI222_X1 U95 ( .A1(data_out_b[9]), .A2(n21), .B1(adder[9]), .B2(n15), .C1(
        n67), .C2(f[9]), .ZN(n68) );
  INV_X1 U96 ( .A(n68), .ZN(n81) );
  NOR4_X1 U97 ( .A1(n51), .A2(n50), .A3(n49), .A4(n48), .ZN(n76) );
  NOR4_X1 U98 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n53), .ZN(n75) );
  NAND4_X1 U99 ( .A1(n72), .A2(n71), .A3(n70), .A4(n69), .ZN(n73) );
  NOR4_X1 U100 ( .A1(n73), .A2(n65), .A3(n63), .A4(n61), .ZN(n74) );
  NAND3_X1 U101 ( .A1(n76), .A2(n75), .A3(n74), .ZN(n78) );
  NAND3_X1 U102 ( .A1(wr_en_y), .A2(n78), .A3(n77), .ZN(n242) );
  OAI22_X1 U103 ( .A1(n182), .A2(n243), .B1(n214), .B2(n242), .ZN(n181) );
  OAI22_X1 U104 ( .A1(n183), .A2(n243), .B1(n215), .B2(n242), .ZN(n180) );
  OAI22_X1 U105 ( .A1(n184), .A2(n243), .B1(n216), .B2(n242), .ZN(n179) );
  OAI22_X1 U106 ( .A1(n192), .A2(n243), .B1(n220), .B2(n242), .ZN(n171) );
  OAI22_X1 U107 ( .A1(n193), .A2(n243), .B1(n221), .B2(n242), .ZN(n170) );
  OAI22_X1 U108 ( .A1(n194), .A2(n243), .B1(n222), .B2(n242), .ZN(n169) );
  OAI22_X1 U109 ( .A1(n195), .A2(n243), .B1(n223), .B2(n242), .ZN(n168) );
  OAI22_X1 U110 ( .A1(n196), .A2(n243), .B1(n224), .B2(n242), .ZN(n167) );
  OAI22_X1 U111 ( .A1(n197), .A2(n243), .B1(n77), .B2(n242), .ZN(n116) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_5_DW_mult_tc_1 ( a, b, 
        product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n9, n12, n13, n16, n18, n19, n23, n25, n27, n29, n31, n32,
         n34, n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n62, n63, n64, n65, n67,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n93, n95, n96, n97, n98,
         n99, n103, n104, n105, n106, n107, n109, n111, n112, n113, n114, n115,
         n117, n119, n120, n122, n127, n133, n135, n139, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n237, n249, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n418,
         n419, n420, n421, n422, n423, n424, n426, n427, n429, n430, n432,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U148 ( .A(n265), .B(n144), .Z(n145) );
  XOR2_X1 U150 ( .A(n271), .B(n146), .Z(n147) );
  XOR2_X1 U152 ( .A(n301), .B(n148), .Z(n149) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U161 ( .A(n177), .B(n168), .CI(n166), .CO(n163), .S(n164) );
  FA_X1 U162 ( .A(n170), .B(n172), .CI(n179), .CO(n165), .S(n166) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n263), .CI(n291), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n317), .B(n252), .CO(n173), .S(n174) );
  FA_X1 U167 ( .A(n180), .B(n187), .CI(n178), .CO(n175), .S(n176) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U169 ( .A(n193), .B(n282), .CI(n191), .CO(n179), .S(n180) );
  FA_X1 U170 ( .A(n268), .B(n292), .CI(n274), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U174 ( .A(n275), .B(n293), .CI(n194), .CO(n189), .S(n190) );
  FA_X1 U175 ( .A(n305), .B(n283), .CI(n253), .CO(n191), .S(n192) );
  HA_X1 U176 ( .A(n269), .B(n319), .CO(n193), .S(n194) );
  FA_X1 U177 ( .A(n205), .B(n200), .CI(n198), .CO(n195), .S(n196) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U179 ( .A(n276), .B(n294), .CI(n284), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n306), .B(n270), .CI(n320), .CO(n201), .S(n202) );
  FA_X1 U181 ( .A(n208), .B(n213), .CI(n206), .CO(n203), .S(n204) );
  FA_X1 U182 ( .A(n215), .B(n307), .CI(n210), .CO(n205), .S(n206) );
  FA_X1 U183 ( .A(n295), .B(n285), .CI(n254), .CO(n207), .S(n208) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n308), .B(n278), .CI(n322), .CO(n215), .S(n216) );
  FA_X1 U188 ( .A(n225), .B(n222), .CI(n220), .CO(n217), .S(n218) );
  FA_X1 U189 ( .A(n255), .B(n309), .CI(n297), .CO(n219), .S(n220) );
  HA_X1 U190 ( .A(n287), .B(n323), .CO(n221), .S(n222) );
  FA_X1 U191 ( .A(n229), .B(n298), .CI(n226), .CO(n223), .S(n224) );
  FA_X1 U192 ( .A(n324), .B(n288), .CI(n310), .CO(n225), .S(n226) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  HA_X1 U194 ( .A(n325), .B(n311), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n312), .B(n300), .CI(n326), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  CLKBUF_X1 U414 ( .A(n574), .Z(n490) );
  INV_X1 U415 ( .A(n103), .ZN(n491) );
  AND2_X1 U416 ( .A1(n224), .A2(n227), .ZN(n556) );
  OR2_X1 U417 ( .A1(n176), .A2(n185), .ZN(n492) );
  BUF_X2 U418 ( .A(n9), .Z(n493) );
  OAI21_X1 U419 ( .B1(n524), .B2(n89), .A(n90), .ZN(n494) );
  OAI21_X1 U420 ( .B1(n99), .B2(n97), .A(n98), .ZN(n96) );
  BUF_X2 U421 ( .A(n9), .Z(n532) );
  OR2_X1 U422 ( .A1(n164), .A2(n175), .ZN(n495) );
  OR2_X1 U423 ( .A1(n329), .A2(n258), .ZN(n496) );
  INV_X2 U424 ( .A(n578), .ZN(n508) );
  CLKBUF_X3 U425 ( .A(n13), .Z(n521) );
  OR2_X1 U426 ( .A1(n550), .A2(n531), .ZN(n497) );
  INV_X1 U427 ( .A(n512), .ZN(n498) );
  OR2_X1 U428 ( .A1(n550), .A2(n531), .ZN(n552) );
  OR2_X1 U429 ( .A1(n550), .A2(n531), .ZN(n551) );
  XNOR2_X1 U430 ( .A(n574), .B(a[2]), .ZN(n499) );
  XOR2_X1 U431 ( .A(n575), .B(a[4]), .Z(n511) );
  OR2_X1 U432 ( .A1(n218), .A2(n223), .ZN(n500) );
  CLKBUF_X2 U433 ( .A(n19), .Z(n513) );
  OR2_X1 U434 ( .A1(n196), .A2(n203), .ZN(n501) );
  CLKBUF_X1 U435 ( .A(n541), .Z(n502) );
  BUF_X1 U436 ( .A(n27), .Z(n525) );
  INV_X1 U437 ( .A(n574), .ZN(n572) );
  INV_X2 U438 ( .A(n582), .ZN(n581) );
  NOR2_X1 U439 ( .A1(n164), .A2(n175), .ZN(n503) );
  NOR2_X1 U440 ( .A1(n164), .A2(n175), .ZN(n75) );
  NAND2_X1 U441 ( .A1(n430), .A2(n509), .ZN(n504) );
  NAND2_X1 U442 ( .A1(n430), .A2(n509), .ZN(n23) );
  INV_X1 U443 ( .A(n574), .ZN(n505) );
  INV_X1 U444 ( .A(n574), .ZN(n506) );
  CLKBUF_X1 U445 ( .A(n27), .Z(n507) );
  INV_X1 U446 ( .A(n578), .ZN(n577) );
  AOI21_X1 U447 ( .B1(n542), .B2(n80), .A(n81), .ZN(n541) );
  XOR2_X1 U448 ( .A(n575), .B(a[6]), .Z(n509) );
  OR2_X2 U449 ( .A1(n511), .A2(n512), .ZN(n510) );
  OR2_X2 U450 ( .A1(n511), .A2(n512), .ZN(n18) );
  XNOR2_X1 U451 ( .A(n574), .B(a[4]), .ZN(n512) );
  OR2_X1 U452 ( .A1(n204), .A2(n211), .ZN(n514) );
  INV_X2 U453 ( .A(n7), .ZN(n574) );
  XOR2_X1 U454 ( .A(n571), .B(n249), .Z(n550) );
  INV_X1 U455 ( .A(n540), .ZN(n515) );
  INV_X1 U456 ( .A(n540), .ZN(n516) );
  INV_X1 U457 ( .A(n580), .ZN(n517) );
  INV_X1 U458 ( .A(n580), .ZN(n518) );
  INV_X1 U459 ( .A(n580), .ZN(n579) );
  AOI21_X1 U460 ( .B1(n561), .B2(n553), .A(n491), .ZN(n519) );
  XOR2_X1 U461 ( .A(n574), .B(a[4]), .Z(n16) );
  INV_X1 U462 ( .A(n531), .ZN(n520) );
  INV_X1 U463 ( .A(n531), .ZN(n555) );
  XNOR2_X1 U464 ( .A(n522), .B(n188), .ZN(n186) );
  XNOR2_X1 U465 ( .A(n197), .B(n190), .ZN(n522) );
  XNOR2_X1 U466 ( .A(n523), .B(n192), .ZN(n188) );
  XNOR2_X1 U467 ( .A(n199), .B(n201), .ZN(n523) );
  AOI21_X1 U468 ( .B1(n96), .B2(n558), .A(n93), .ZN(n524) );
  CLKBUF_X1 U469 ( .A(n1), .Z(n543) );
  OR2_X2 U470 ( .A1(n526), .A2(n549), .ZN(n34) );
  XNOR2_X1 U471 ( .A(n517), .B(a[10]), .ZN(n526) );
  XOR2_X1 U472 ( .A(n216), .B(n219), .Z(n527) );
  XOR2_X1 U473 ( .A(n214), .B(n527), .Z(n212) );
  NAND2_X1 U474 ( .A1(n214), .A2(n216), .ZN(n528) );
  NAND2_X1 U475 ( .A1(n214), .A2(n219), .ZN(n529) );
  NAND2_X1 U476 ( .A1(n216), .A2(n219), .ZN(n530) );
  NAND3_X1 U477 ( .A1(n528), .A2(n529), .A3(n530), .ZN(n211) );
  CLKBUF_X1 U478 ( .A(n249), .Z(n531) );
  XNOR2_X1 U479 ( .A(n543), .B(a[2]), .ZN(n533) );
  NAND2_X1 U480 ( .A1(n199), .A2(n201), .ZN(n534) );
  NAND2_X1 U481 ( .A1(n199), .A2(n192), .ZN(n535) );
  NAND2_X1 U482 ( .A1(n201), .A2(n192), .ZN(n536) );
  NAND3_X1 U483 ( .A1(n534), .A2(n535), .A3(n536), .ZN(n187) );
  NAND2_X1 U484 ( .A1(n197), .A2(n190), .ZN(n537) );
  NAND2_X1 U485 ( .A1(n197), .A2(n188), .ZN(n538) );
  NAND2_X1 U486 ( .A1(n190), .A2(n188), .ZN(n539) );
  NAND3_X1 U487 ( .A1(n537), .A2(n538), .A3(n539), .ZN(n185) );
  XNOR2_X1 U488 ( .A(n575), .B(a[6]), .ZN(n540) );
  XNOR2_X1 U489 ( .A(n494), .B(n51), .ZN(product[10]) );
  AOI21_X1 U490 ( .B1(n542), .B2(n80), .A(n81), .ZN(n45) );
  XNOR2_X1 U491 ( .A(n574), .B(a[2]), .ZN(n432) );
  OAI21_X1 U492 ( .B1(n91), .B2(n89), .A(n90), .ZN(n542) );
  OAI21_X1 U493 ( .B1(n524), .B2(n89), .A(n90), .ZN(n88) );
  INV_X1 U494 ( .A(n546), .ZN(n27) );
  BUF_X2 U495 ( .A(n16), .Z(n544) );
  INV_X1 U496 ( .A(n493), .ZN(n545) );
  XNOR2_X1 U497 ( .A(n576), .B(a[8]), .ZN(n546) );
  INV_X1 U498 ( .A(n549), .ZN(n32) );
  NAND2_X2 U499 ( .A1(n429), .A2(n27), .ZN(n29) );
  NAND2_X1 U500 ( .A1(n499), .A2(n533), .ZN(n547) );
  NAND2_X1 U501 ( .A1(n432), .A2(n533), .ZN(n548) );
  NAND2_X1 U502 ( .A1(n432), .A2(n533), .ZN(n12) );
  XNOR2_X1 U503 ( .A(n578), .B(a[10]), .ZN(n549) );
  OR2_X1 U504 ( .A1(n550), .A2(n531), .ZN(n6) );
  CLKBUF_X1 U505 ( .A(n104), .Z(n553) );
  CLKBUF_X1 U506 ( .A(n107), .Z(n554) );
  INV_X1 U507 ( .A(n556), .ZN(n103) );
  INV_X1 U508 ( .A(n571), .ZN(n570) );
  NOR2_X2 U509 ( .A1(n186), .A2(n195), .ZN(n82) );
  XNOR2_X1 U510 ( .A(n543), .B(a[2]), .ZN(n9) );
  NAND2_X1 U511 ( .A1(n557), .A2(n69), .ZN(n47) );
  INV_X1 U512 ( .A(n73), .ZN(n71) );
  AOI21_X1 U513 ( .B1(n74), .B2(n557), .A(n67), .ZN(n65) );
  INV_X1 U514 ( .A(n69), .ZN(n67) );
  NAND2_X1 U515 ( .A1(n73), .A2(n557), .ZN(n64) );
  INV_X1 U516 ( .A(n74), .ZN(n72) );
  INV_X1 U517 ( .A(n95), .ZN(n93) );
  XNOR2_X1 U518 ( .A(n84), .B(n50), .ZN(product[11]) );
  NAND2_X1 U519 ( .A1(n127), .A2(n83), .ZN(n50) );
  NAND2_X1 U520 ( .A1(n501), .A2(n86), .ZN(n51) );
  NAND2_X1 U521 ( .A1(n514), .A2(n90), .ZN(n52) );
  NAND2_X1 U522 ( .A1(n492), .A2(n79), .ZN(n49) );
  OR2_X1 U523 ( .A1(n152), .A2(n163), .ZN(n557) );
  NAND2_X1 U524 ( .A1(n495), .A2(n76), .ZN(n48) );
  OAI21_X1 U525 ( .B1(n503), .B2(n79), .A(n76), .ZN(n74) );
  NOR2_X1 U526 ( .A1(n75), .A2(n78), .ZN(n73) );
  NAND2_X1 U527 ( .A1(n152), .A2(n163), .ZN(n69) );
  OAI21_X1 U528 ( .B1(n113), .B2(n115), .A(n114), .ZN(n112) );
  NAND2_X1 U529 ( .A1(n133), .A2(n106), .ZN(n56) );
  INV_X1 U530 ( .A(n105), .ZN(n133) );
  NAND2_X1 U531 ( .A1(n500), .A2(n98), .ZN(n54) );
  NOR2_X1 U532 ( .A1(n176), .A2(n185), .ZN(n78) );
  NAND2_X1 U533 ( .A1(n561), .A2(n103), .ZN(n55) );
  AOI21_X1 U534 ( .B1(n559), .B2(n120), .A(n117), .ZN(n115) );
  INV_X1 U535 ( .A(n119), .ZN(n117) );
  AOI21_X1 U536 ( .B1(n560), .B2(n112), .A(n109), .ZN(n107) );
  INV_X1 U537 ( .A(n111), .ZN(n109) );
  INV_X1 U538 ( .A(n122), .ZN(n120) );
  NOR2_X1 U539 ( .A1(n196), .A2(n203), .ZN(n85) );
  XNOR2_X1 U540 ( .A(n57), .B(n112), .ZN(product[4]) );
  NAND2_X1 U541 ( .A1(n560), .A2(n111), .ZN(n57) );
  XNOR2_X1 U542 ( .A(n59), .B(n120), .ZN(product[2]) );
  NAND2_X1 U543 ( .A1(n559), .A2(n119), .ZN(n59) );
  NAND2_X1 U544 ( .A1(n176), .A2(n185), .ZN(n79) );
  NAND2_X1 U545 ( .A1(n186), .A2(n195), .ZN(n83) );
  NAND2_X1 U546 ( .A1(n164), .A2(n175), .ZN(n76) );
  NAND2_X1 U547 ( .A1(n196), .A2(n203), .ZN(n86) );
  OR2_X1 U548 ( .A1(n212), .A2(n217), .ZN(n558) );
  NAND2_X1 U549 ( .A1(n204), .A2(n211), .ZN(n90) );
  NAND2_X1 U550 ( .A1(n212), .A2(n217), .ZN(n95) );
  NAND2_X1 U551 ( .A1(n135), .A2(n114), .ZN(n58) );
  INV_X1 U552 ( .A(n113), .ZN(n135) );
  XNOR2_X1 U553 ( .A(n63), .B(n46), .ZN(product[15]) );
  NAND2_X1 U554 ( .A1(n562), .A2(n62), .ZN(n46) );
  OR2_X1 U555 ( .A1(n328), .A2(n314), .ZN(n559) );
  OR2_X1 U556 ( .A1(n232), .A2(n233), .ZN(n560) );
  NOR2_X1 U557 ( .A1(n228), .A2(n231), .ZN(n105) );
  NOR2_X1 U558 ( .A1(n218), .A2(n223), .ZN(n97) );
  NAND2_X1 U559 ( .A1(n228), .A2(n231), .ZN(n106) );
  NAND2_X1 U560 ( .A1(n218), .A2(n223), .ZN(n98) );
  INV_X1 U561 ( .A(n37), .ZN(n237) );
  OR2_X1 U562 ( .A1(n224), .A2(n227), .ZN(n561) );
  INV_X1 U563 ( .A(n41), .ZN(n235) );
  OR2_X1 U564 ( .A1(n151), .A2(n139), .ZN(n562) );
  AND2_X1 U565 ( .A1(n496), .A2(n122), .ZN(product[1]) );
  XNOR2_X1 U566 ( .A(n579), .B(a[12]), .ZN(n37) );
  XNOR2_X1 U567 ( .A(n581), .B(a[14]), .ZN(n41) );
  OR2_X1 U568 ( .A1(n43), .A2(n574), .ZN(n392) );
  XNOR2_X1 U569 ( .A(n513), .B(n43), .ZN(n363) );
  XNOR2_X1 U570 ( .A(n508), .B(n43), .ZN(n352) );
  AND2_X1 U571 ( .A1(n569), .A2(n546), .ZN(n278) );
  AND2_X1 U572 ( .A1(n569), .A2(n237), .ZN(n264) );
  OR2_X1 U573 ( .A1(n43), .A2(n575), .ZN(n377) );
  XNOR2_X1 U574 ( .A(n155), .B(n564), .ZN(n139) );
  XNOR2_X1 U575 ( .A(n153), .B(n141), .ZN(n564) );
  XNOR2_X1 U576 ( .A(n157), .B(n565), .ZN(n141) );
  XNOR2_X1 U577 ( .A(n145), .B(n143), .ZN(n565) );
  OAI22_X1 U578 ( .A1(n39), .A2(n336), .B1(n37), .B2(n335), .ZN(n263) );
  OAI22_X1 U579 ( .A1(n34), .A2(n342), .B1(n341), .B2(n32), .ZN(n268) );
  OAI22_X1 U580 ( .A1(n39), .A2(n582), .B1(n337), .B2(n37), .ZN(n252) );
  OR2_X1 U581 ( .A1(n43), .A2(n582), .ZN(n337) );
  OAI22_X1 U582 ( .A1(n34), .A2(n343), .B1(n342), .B2(n32), .ZN(n269) );
  XNOR2_X1 U583 ( .A(n517), .B(n43), .ZN(n343) );
  OAI22_X1 U584 ( .A1(n42), .A2(n584), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U585 ( .A1(n43), .A2(n584), .ZN(n332) );
  AND2_X1 U586 ( .A1(n569), .A2(n512), .ZN(n300) );
  XOR2_X1 U587 ( .A(n577), .B(a[8]), .Z(n429) );
  XNOR2_X1 U588 ( .A(n159), .B(n566), .ZN(n142) );
  XNOR2_X1 U589 ( .A(n315), .B(n261), .ZN(n566) );
  XNOR2_X1 U590 ( .A(n581), .B(n43), .ZN(n336) );
  XOR2_X1 U591 ( .A(n19), .B(a[6]), .Z(n430) );
  NAND2_X1 U592 ( .A1(n427), .A2(n37), .ZN(n39) );
  XOR2_X1 U593 ( .A(n581), .B(a[12]), .Z(n427) );
  XNOR2_X1 U594 ( .A(n521), .B(n43), .ZN(n376) );
  OAI22_X1 U595 ( .A1(n34), .A2(n341), .B1(n340), .B2(n32), .ZN(n267) );
  AND2_X1 U596 ( .A1(n569), .A2(n235), .ZN(n260) );
  OAI22_X1 U597 ( .A1(n39), .A2(n335), .B1(n37), .B2(n334), .ZN(n262) );
  AND2_X1 U598 ( .A1(n569), .A2(n540), .ZN(n288) );
  AND2_X1 U599 ( .A1(n569), .A2(n549), .ZN(n270) );
  INV_X1 U600 ( .A(n25), .ZN(n578) );
  OAI22_X1 U601 ( .A1(n34), .A2(n580), .B1(n344), .B2(n32), .ZN(n253) );
  INV_X1 U602 ( .A(n13), .ZN(n575) );
  OAI22_X1 U603 ( .A1(n34), .A2(n340), .B1(n339), .B2(n32), .ZN(n266) );
  NAND2_X1 U604 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U605 ( .A(n583), .B(a[14]), .Z(n426) );
  AND2_X1 U606 ( .A1(n569), .A2(n545), .ZN(n314) );
  OR2_X1 U607 ( .A1(n43), .A2(n580), .ZN(n344) );
  AND2_X1 U608 ( .A1(n569), .A2(n249), .ZN(product[0]) );
  OR2_X1 U609 ( .A1(n43), .A2(n576), .ZN(n364) );
  OR2_X1 U610 ( .A1(n43), .A2(n578), .ZN(n353) );
  XNOR2_X1 U611 ( .A(n513), .B(b[9]), .ZN(n354) );
  OAI22_X1 U612 ( .A1(n39), .A2(n334), .B1(n37), .B2(n333), .ZN(n261) );
  XNOR2_X1 U613 ( .A(n581), .B(n422), .ZN(n333) );
  XNOR2_X1 U614 ( .A(n521), .B(b[11]), .ZN(n365) );
  XNOR2_X1 U615 ( .A(n518), .B(n424), .ZN(n342) );
  XNOR2_X1 U616 ( .A(n517), .B(n423), .ZN(n341) );
  XNOR2_X1 U617 ( .A(n518), .B(n422), .ZN(n340) );
  XNOR2_X1 U618 ( .A(n518), .B(n421), .ZN(n339) );
  XNOR2_X1 U619 ( .A(n581), .B(n424), .ZN(n335) );
  XNOR2_X1 U620 ( .A(n581), .B(n423), .ZN(n334) );
  OAI22_X1 U621 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U622 ( .A(n583), .B(n424), .ZN(n330) );
  XNOR2_X1 U623 ( .A(n583), .B(n43), .ZN(n331) );
  XNOR2_X1 U624 ( .A(n508), .B(n418), .ZN(n345) );
  OAI22_X1 U625 ( .A1(n34), .A2(n339), .B1(n338), .B2(n32), .ZN(n265) );
  XNOR2_X1 U626 ( .A(n518), .B(n420), .ZN(n338) );
  XNOR2_X1 U627 ( .A(n506), .B(b[13]), .ZN(n378) );
  XNOR2_X1 U628 ( .A(n513), .B(n424), .ZN(n362) );
  XNOR2_X1 U629 ( .A(n508), .B(n424), .ZN(n351) );
  XNOR2_X1 U630 ( .A(n573), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U631 ( .A(n573), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U632 ( .A(n572), .B(n418), .ZN(n384) );
  XNOR2_X1 U633 ( .A(n506), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U634 ( .A(n506), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U635 ( .A(n505), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U636 ( .A(n572), .B(n419), .ZN(n385) );
  XNOR2_X1 U637 ( .A(n521), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U638 ( .A(n521), .B(n418), .ZN(n369) );
  XNOR2_X1 U639 ( .A(n521), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U640 ( .A(n521), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U641 ( .A(n513), .B(n423), .ZN(n361) );
  XNOR2_X1 U642 ( .A(n513), .B(n422), .ZN(n360) );
  XNOR2_X1 U643 ( .A(n508), .B(n422), .ZN(n349) );
  XNOR2_X1 U644 ( .A(n508), .B(n423), .ZN(n350) );
  XNOR2_X1 U645 ( .A(n513), .B(n421), .ZN(n359) );
  XNOR2_X1 U646 ( .A(n513), .B(n420), .ZN(n358) );
  XNOR2_X1 U647 ( .A(n508), .B(n421), .ZN(n348) );
  XNOR2_X1 U648 ( .A(n508), .B(n420), .ZN(n347) );
  XNOR2_X1 U649 ( .A(n513), .B(n418), .ZN(n356) );
  XNOR2_X1 U650 ( .A(n567), .B(b[14]), .ZN(n394) );
  XNOR2_X1 U651 ( .A(n568), .B(b[11]), .ZN(n397) );
  XNOR2_X1 U652 ( .A(n568), .B(b[13]), .ZN(n395) );
  XNOR2_X1 U653 ( .A(n508), .B(n419), .ZN(n346) );
  XNOR2_X1 U654 ( .A(n513), .B(n419), .ZN(n357) );
  XNOR2_X1 U655 ( .A(n513), .B(b[8]), .ZN(n355) );
  XNOR2_X1 U656 ( .A(n567), .B(b[12]), .ZN(n396) );
  BUF_X1 U657 ( .A(n43), .Z(n569) );
  XNOR2_X1 U658 ( .A(n567), .B(b[15]), .ZN(n393) );
  INV_X1 U659 ( .A(n571), .ZN(n567) );
  INV_X1 U660 ( .A(n571), .ZN(n568) );
  INV_X1 U661 ( .A(n19), .ZN(n576) );
  OR2_X1 U662 ( .A1(n43), .A2(n571), .ZN(n409) );
  INV_X1 U663 ( .A(n1), .ZN(n571) );
  NOR2_X1 U664 ( .A1(n204), .A2(n211), .ZN(n89) );
  OAI22_X1 U665 ( .A1(n29), .A2(n346), .B1(n345), .B2(n525), .ZN(n271) );
  OAI22_X1 U666 ( .A1(n29), .A2(n350), .B1(n349), .B2(n525), .ZN(n275) );
  OAI22_X1 U667 ( .A1(n29), .A2(n351), .B1(n350), .B2(n507), .ZN(n276) );
  OAI22_X1 U668 ( .A1(n29), .A2(n347), .B1(n346), .B2(n525), .ZN(n272) );
  OAI22_X1 U669 ( .A1(n29), .A2(n348), .B1(n347), .B2(n525), .ZN(n273) );
  OAI22_X1 U670 ( .A1(n29), .A2(n349), .B1(n348), .B2(n525), .ZN(n274) );
  OAI22_X1 U671 ( .A1(n29), .A2(n578), .B1(n353), .B2(n507), .ZN(n254) );
  OAI22_X1 U672 ( .A1(n29), .A2(n352), .B1(n351), .B2(n507), .ZN(n277) );
  XNOR2_X1 U673 ( .A(n77), .B(n48), .ZN(product[13]) );
  INV_X1 U674 ( .A(n82), .ZN(n127) );
  NOR2_X1 U675 ( .A1(n82), .A2(n85), .ZN(n80) );
  OAI21_X1 U676 ( .B1(n82), .B2(n86), .A(n83), .ZN(n81) );
  OAI22_X1 U677 ( .A1(n504), .A2(n358), .B1(n357), .B2(n516), .ZN(n282) );
  OAI22_X1 U678 ( .A1(n504), .A2(n356), .B1(n355), .B2(n515), .ZN(n280) );
  OAI22_X1 U679 ( .A1(n504), .A2(n362), .B1(n361), .B2(n515), .ZN(n286) );
  OAI22_X1 U680 ( .A1(n23), .A2(n576), .B1(n364), .B2(n515), .ZN(n255) );
  OAI22_X1 U681 ( .A1(n23), .A2(n357), .B1(n356), .B2(n516), .ZN(n281) );
  OAI22_X1 U682 ( .A1(n504), .A2(n355), .B1(n354), .B2(n515), .ZN(n279) );
  OAI22_X1 U683 ( .A1(n504), .A2(n363), .B1(n362), .B2(n515), .ZN(n287) );
  OAI22_X1 U684 ( .A1(n504), .A2(n360), .B1(n359), .B2(n516), .ZN(n284) );
  OAI22_X1 U685 ( .A1(n23), .A2(n361), .B1(n360), .B2(n516), .ZN(n285) );
  OAI22_X1 U686 ( .A1(n23), .A2(n359), .B1(n358), .B2(n516), .ZN(n283) );
  NAND2_X1 U687 ( .A1(n558), .A2(n95), .ZN(n53) );
  XNOR2_X1 U688 ( .A(n70), .B(n47), .ZN(product[14]) );
  XNOR2_X1 U689 ( .A(n521), .B(n423), .ZN(n374) );
  XNOR2_X1 U690 ( .A(n521), .B(n424), .ZN(n375) );
  XNOR2_X1 U691 ( .A(n521), .B(n422), .ZN(n373) );
  XNOR2_X1 U692 ( .A(n521), .B(n421), .ZN(n372) );
  XNOR2_X1 U693 ( .A(n521), .B(n419), .ZN(n370) );
  XNOR2_X1 U694 ( .A(n521), .B(n420), .ZN(n371) );
  OAI21_X1 U695 ( .B1(n87), .B2(n85), .A(n86), .ZN(n84) );
  XNOR2_X1 U696 ( .A(n55), .B(n553), .ZN(product[6]) );
  AOI21_X1 U697 ( .B1(n561), .B2(n104), .A(n556), .ZN(n99) );
  NAND2_X1 U698 ( .A1(n151), .A2(n139), .ZN(n62) );
  OAI22_X1 U699 ( .A1(n18), .A2(n370), .B1(n369), .B2(n498), .ZN(n293) );
  OAI22_X1 U700 ( .A1(n18), .A2(n367), .B1(n366), .B2(n498), .ZN(n290) );
  OAI22_X1 U701 ( .A1(n510), .A2(n368), .B1(n367), .B2(n544), .ZN(n291) );
  OAI22_X1 U702 ( .A1(n510), .A2(n375), .B1(n374), .B2(n498), .ZN(n298) );
  OAI22_X1 U703 ( .A1(n510), .A2(n373), .B1(n372), .B2(n498), .ZN(n296) );
  OAI22_X1 U704 ( .A1(n510), .A2(n369), .B1(n368), .B2(n544), .ZN(n292) );
  OAI22_X1 U705 ( .A1(n18), .A2(n372), .B1(n371), .B2(n544), .ZN(n295) );
  OAI22_X1 U706 ( .A1(n18), .A2(n374), .B1(n373), .B2(n544), .ZN(n297) );
  OAI22_X1 U707 ( .A1(n510), .A2(n371), .B1(n370), .B2(n498), .ZN(n294) );
  OAI22_X1 U708 ( .A1(n18), .A2(n575), .B1(n377), .B2(n544), .ZN(n256) );
  OAI22_X1 U709 ( .A1(n510), .A2(n376), .B1(n375), .B2(n544), .ZN(n299) );
  OAI22_X1 U710 ( .A1(n18), .A2(n366), .B1(n365), .B2(n544), .ZN(n289) );
  XNOR2_X1 U711 ( .A(n505), .B(n420), .ZN(n386) );
  XNOR2_X1 U712 ( .A(n505), .B(n43), .ZN(n391) );
  XNOR2_X1 U713 ( .A(n573), .B(n422), .ZN(n388) );
  XNOR2_X1 U714 ( .A(n572), .B(n421), .ZN(n387) );
  XNOR2_X1 U715 ( .A(n506), .B(n423), .ZN(n389) );
  XNOR2_X1 U716 ( .A(n505), .B(n424), .ZN(n390) );
  XOR2_X1 U717 ( .A(n56), .B(n554), .Z(product[5]) );
  OAI21_X1 U718 ( .B1(n105), .B2(n107), .A(n106), .ZN(n104) );
  XNOR2_X1 U719 ( .A(n567), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U720 ( .A(n567), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U721 ( .A(n570), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U722 ( .A(n568), .B(n418), .ZN(n401) );
  XNOR2_X1 U723 ( .A(n570), .B(n420), .ZN(n403) );
  XNOR2_X1 U724 ( .A(n570), .B(n419), .ZN(n402) );
  XNOR2_X1 U725 ( .A(n567), .B(n422), .ZN(n405) );
  XNOR2_X1 U726 ( .A(n568), .B(n421), .ZN(n404) );
  XNOR2_X1 U727 ( .A(n570), .B(n423), .ZN(n406) );
  XNOR2_X1 U728 ( .A(n568), .B(n43), .ZN(n408) );
  XNOR2_X1 U729 ( .A(n567), .B(n424), .ZN(n407) );
  NAND2_X1 U730 ( .A1(n232), .A2(n233), .ZN(n111) );
  INV_X1 U731 ( .A(n88), .ZN(n87) );
  NAND2_X1 U732 ( .A1(n328), .A2(n314), .ZN(n119) );
  NOR2_X1 U733 ( .A1(n234), .A2(n257), .ZN(n113) );
  OAI21_X1 U734 ( .B1(n64), .B2(n502), .A(n65), .ZN(n63) );
  OAI21_X1 U735 ( .B1(n541), .B2(n71), .A(n72), .ZN(n70) );
  OAI21_X1 U736 ( .B1(n541), .B2(n78), .A(n79), .ZN(n77) );
  XOR2_X1 U737 ( .A(n45), .B(n49), .Z(product[12]) );
  XOR2_X1 U738 ( .A(n91), .B(n52), .Z(product[9]) );
  XNOR2_X1 U739 ( .A(n96), .B(n53), .ZN(product[8]) );
  AOI21_X1 U740 ( .B1(n96), .B2(n558), .A(n93), .ZN(n91) );
  XOR2_X1 U741 ( .A(n58), .B(n115), .Z(product[3]) );
  OAI22_X1 U742 ( .A1(n551), .A2(n395), .B1(n394), .B2(n520), .ZN(n316) );
  OAI22_X1 U743 ( .A1(n552), .A2(n394), .B1(n393), .B2(n520), .ZN(n315) );
  OAI22_X1 U744 ( .A1(n497), .A2(n396), .B1(n395), .B2(n520), .ZN(n317) );
  OAI22_X1 U745 ( .A1(n497), .A2(n397), .B1(n396), .B2(n520), .ZN(n318) );
  OAI22_X1 U746 ( .A1(n551), .A2(n398), .B1(n397), .B2(n555), .ZN(n319) );
  OAI22_X1 U747 ( .A1(n551), .A2(n400), .B1(n399), .B2(n555), .ZN(n321) );
  OAI22_X1 U748 ( .A1(n6), .A2(n399), .B1(n398), .B2(n555), .ZN(n320) );
  OAI22_X1 U749 ( .A1(n551), .A2(n401), .B1(n400), .B2(n555), .ZN(n322) );
  OAI22_X1 U750 ( .A1(n552), .A2(n402), .B1(n401), .B2(n520), .ZN(n323) );
  NAND2_X1 U751 ( .A1(n329), .A2(n258), .ZN(n122) );
  OAI22_X1 U752 ( .A1(n497), .A2(n404), .B1(n403), .B2(n555), .ZN(n325) );
  OAI22_X1 U753 ( .A1(n6), .A2(n403), .B1(n555), .B2(n402), .ZN(n324) );
  OAI22_X1 U754 ( .A1(n552), .A2(n406), .B1(n405), .B2(n555), .ZN(n327) );
  OAI22_X1 U755 ( .A1(n497), .A2(n405), .B1(n404), .B2(n555), .ZN(n326) );
  OAI22_X1 U756 ( .A1(n552), .A2(n407), .B1(n406), .B2(n520), .ZN(n328) );
  OAI22_X1 U757 ( .A1(n551), .A2(n408), .B1(n407), .B2(n555), .ZN(n329) );
  OAI22_X1 U758 ( .A1(n497), .A2(n571), .B1(n409), .B2(n555), .ZN(n258) );
  XOR2_X1 U759 ( .A(n519), .B(n54), .Z(product[7]) );
  OAI22_X1 U760 ( .A1(n547), .A2(n379), .B1(n378), .B2(n493), .ZN(n301) );
  OAI22_X1 U761 ( .A1(n548), .A2(n380), .B1(n379), .B2(n493), .ZN(n302) );
  OAI22_X1 U762 ( .A1(n12), .A2(n385), .B1(n384), .B2(n532), .ZN(n307) );
  OAI22_X1 U763 ( .A1(n548), .A2(n382), .B1(n381), .B2(n532), .ZN(n304) );
  OAI22_X1 U764 ( .A1(n547), .A2(n381), .B1(n380), .B2(n532), .ZN(n303) );
  NAND2_X1 U765 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U766 ( .A1(n547), .A2(n383), .B1(n382), .B2(n493), .ZN(n305) );
  OAI22_X1 U767 ( .A1(n384), .A2(n547), .B1(n383), .B2(n493), .ZN(n306) );
  OAI22_X1 U768 ( .A1(n547), .A2(n386), .B1(n385), .B2(n493), .ZN(n308) );
  OAI22_X1 U769 ( .A1(n548), .A2(n387), .B1(n386), .B2(n493), .ZN(n309) );
  OAI22_X1 U770 ( .A1(n548), .A2(n490), .B1(n392), .B2(n532), .ZN(n257) );
  OAI22_X1 U771 ( .A1(n12), .A2(n389), .B1(n388), .B2(n532), .ZN(n311) );
  OAI22_X1 U772 ( .A1(n12), .A2(n388), .B1(n387), .B2(n532), .ZN(n310) );
  OAI22_X1 U773 ( .A1(n12), .A2(n390), .B1(n389), .B2(n532), .ZN(n312) );
  OAI22_X1 U774 ( .A1(n548), .A2(n391), .B1(n390), .B2(n532), .ZN(n313) );
  INV_X1 U775 ( .A(n574), .ZN(n573) );
  INV_X1 U776 ( .A(n31), .ZN(n580) );
  INV_X1 U777 ( .A(n36), .ZN(n582) );
  INV_X1 U778 ( .A(n584), .ZN(n583) );
  INV_X1 U779 ( .A(n40), .ZN(n584) );
  XOR2_X1 U780 ( .A(n259), .B(n251), .Z(n148) );
  XOR2_X1 U781 ( .A(n289), .B(n279), .Z(n146) );
  XOR2_X1 U782 ( .A(n149), .B(n147), .Z(n144) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_5_DW01_add_2 ( A, B, CI, SUM, 
        CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n18,
         n19, n20, n21, n25, n26, n27, n28, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n48, n49, n51, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n69, n71, n72, n73, n74, n75,
         n77, n79, n80, n81, n82, n83, n85, n87, n88, n90, n94, n95, n99, n100,
         n102, n104, n161, n162, n163, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182;

  OR2_X1 U126 ( .A1(A[10]), .A2(B[10]), .ZN(n161) );
  OR2_X1 U127 ( .A1(A[10]), .A2(B[10]), .ZN(n180) );
  BUF_X1 U128 ( .A(n39), .Z(n162) );
  XNOR2_X1 U129 ( .A(n163), .B(n41), .ZN(SUM[11]) );
  AND2_X1 U130 ( .A1(n95), .A2(n40), .ZN(n163) );
  AND2_X1 U131 ( .A1(n176), .A2(n90), .ZN(SUM[0]) );
  OR2_X1 U132 ( .A1(A[15]), .A2(B[15]), .ZN(n165) );
  OR2_X1 U133 ( .A1(A[8]), .A2(B[8]), .ZN(n166) );
  NOR2_X1 U134 ( .A1(n172), .A2(n39), .ZN(n167) );
  AND2_X1 U135 ( .A1(A[10]), .A2(B[10]), .ZN(n173) );
  INV_X1 U136 ( .A(n169), .ZN(n25) );
  AND2_X1 U137 ( .A1(A[9]), .A2(B[9]), .ZN(n51) );
  INV_X1 U138 ( .A(n173), .ZN(n48) );
  OR2_X1 U139 ( .A1(A[14]), .A2(B[14]), .ZN(n168) );
  AND2_X1 U140 ( .A1(A[14]), .A2(B[14]), .ZN(n169) );
  OR2_X1 U141 ( .A1(A[13]), .A2(B[13]), .ZN(n170) );
  NOR2_X2 U142 ( .A1(A[11]), .A2(B[11]), .ZN(n39) );
  AND2_X1 U143 ( .A1(A[13]), .A2(B[13]), .ZN(n171) );
  NOR2_X1 U144 ( .A1(A[12]), .A2(B[12]), .ZN(n172) );
  NOR2_X1 U145 ( .A1(A[12]), .A2(B[12]), .ZN(n36) );
  AOI21_X1 U146 ( .B1(n34), .B2(n42), .A(n35), .ZN(n174) );
  AOI21_X1 U147 ( .B1(n167), .B2(n42), .A(n35), .ZN(n175) );
  OR2_X1 U148 ( .A1(A[0]), .A2(B[0]), .ZN(n176) );
  INV_X1 U149 ( .A(n64), .ZN(n63) );
  INV_X1 U150 ( .A(n55), .ZN(n54) );
  INV_X1 U151 ( .A(n42), .ZN(n41) );
  AOI21_X1 U152 ( .B1(n178), .B2(n88), .A(n85), .ZN(n83) );
  INV_X1 U153 ( .A(n87), .ZN(n85) );
  AOI21_X1 U154 ( .B1(n56), .B2(n64), .A(n57), .ZN(n55) );
  NOR2_X1 U155 ( .A1(n58), .A2(n61), .ZN(n56) );
  OAI21_X1 U156 ( .B1(n58), .B2(n62), .A(n59), .ZN(n57) );
  OAI21_X1 U157 ( .B1(n83), .B2(n81), .A(n82), .ZN(n80) );
  AOI21_X1 U158 ( .B1(n182), .B2(n72), .A(n69), .ZN(n67) );
  INV_X1 U159 ( .A(n71), .ZN(n69) );
  OAI21_X1 U160 ( .B1(n75), .B2(n73), .A(n74), .ZN(n72) );
  AOI21_X1 U161 ( .B1(n54), .B2(n181), .A(n51), .ZN(n49) );
  INV_X1 U162 ( .A(n90), .ZN(n88) );
  OAI21_X1 U163 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  AOI21_X1 U164 ( .B1(n177), .B2(n80), .A(n77), .ZN(n75) );
  INV_X1 U165 ( .A(n79), .ZN(n77) );
  NAND2_X1 U166 ( .A1(n166), .A2(n59), .ZN(n8) );
  NAND2_X1 U167 ( .A1(n102), .A2(n74), .ZN(n12) );
  INV_X1 U168 ( .A(n73), .ZN(n102) );
  NAND2_X1 U169 ( .A1(n99), .A2(n62), .ZN(n9) );
  INV_X1 U170 ( .A(n61), .ZN(n99) );
  NAND2_X1 U171 ( .A1(n104), .A2(n82), .ZN(n14) );
  INV_X1 U172 ( .A(n81), .ZN(n104) );
  NAND2_X1 U173 ( .A1(n182), .A2(n71), .ZN(n11) );
  NAND2_X1 U174 ( .A1(n177), .A2(n79), .ZN(n13) );
  NAND2_X1 U175 ( .A1(n178), .A2(n87), .ZN(n15) );
  NAND2_X1 U176 ( .A1(n100), .A2(n66), .ZN(n10) );
  INV_X1 U177 ( .A(n65), .ZN(n100) );
  XNOR2_X1 U178 ( .A(n11), .B(n72), .ZN(SUM[5]) );
  XOR2_X1 U179 ( .A(n12), .B(n75), .Z(SUM[4]) );
  XOR2_X1 U180 ( .A(n14), .B(n83), .Z(SUM[2]) );
  NAND2_X1 U181 ( .A1(n94), .A2(n37), .ZN(n4) );
  XOR2_X1 U182 ( .A(n49), .B(n6), .Z(SUM[10]) );
  NOR2_X1 U183 ( .A1(A[7]), .A2(B[7]), .ZN(n61) );
  NOR2_X1 U184 ( .A1(A[8]), .A2(B[8]), .ZN(n58) );
  NOR2_X1 U185 ( .A1(A[4]), .A2(B[4]), .ZN(n73) );
  NOR2_X1 U186 ( .A1(A[2]), .A2(B[2]), .ZN(n81) );
  NAND2_X1 U187 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  NAND2_X1 U188 ( .A1(A[11]), .A2(B[11]), .ZN(n40) );
  OR2_X1 U189 ( .A1(A[3]), .A2(B[3]), .ZN(n177) );
  OR2_X1 U190 ( .A1(A[1]), .A2(B[1]), .ZN(n178) );
  NAND2_X1 U191 ( .A1(A[7]), .A2(B[7]), .ZN(n62) );
  OR2_X1 U192 ( .A1(A[14]), .A2(B[14]), .ZN(n179) );
  OR2_X1 U193 ( .A1(A[9]), .A2(B[9]), .ZN(n181) );
  NAND2_X1 U194 ( .A1(A[12]), .A2(B[12]), .ZN(n37) );
  XNOR2_X1 U195 ( .A(n13), .B(n80), .ZN(SUM[3]) );
  NOR2_X1 U196 ( .A1(A[6]), .A2(B[6]), .ZN(n65) );
  OR2_X1 U197 ( .A1(A[5]), .A2(B[5]), .ZN(n182) );
  NAND2_X1 U198 ( .A1(A[8]), .A2(B[8]), .ZN(n59) );
  NAND2_X1 U199 ( .A1(A[4]), .A2(B[4]), .ZN(n74) );
  NAND2_X1 U200 ( .A1(A[2]), .A2(B[2]), .ZN(n82) );
  NAND2_X1 U201 ( .A1(A[3]), .A2(B[3]), .ZN(n79) );
  NAND2_X1 U202 ( .A1(A[5]), .A2(B[5]), .ZN(n71) );
  NAND2_X1 U203 ( .A1(A[1]), .A2(B[1]), .ZN(n87) );
  NAND2_X1 U204 ( .A1(A[0]), .A2(B[0]), .ZN(n90) );
  NAND2_X1 U205 ( .A1(A[6]), .A2(B[6]), .ZN(n66) );
  NAND2_X1 U206 ( .A1(A[9]), .A2(B[9]), .ZN(n53) );
  XNOR2_X1 U207 ( .A(n54), .B(n7), .ZN(SUM[9]) );
  XNOR2_X1 U208 ( .A(n60), .B(n8), .ZN(SUM[8]) );
  XOR2_X1 U209 ( .A(n63), .B(n9), .Z(SUM[7]) );
  XNOR2_X1 U210 ( .A(n15), .B(n88), .ZN(SUM[1]) );
  NAND2_X1 U211 ( .A1(n165), .A2(n18), .ZN(n1) );
  NAND2_X1 U212 ( .A1(n170), .A2(n28), .ZN(n3) );
  NAND2_X1 U213 ( .A1(n181), .A2(n53), .ZN(n7) );
  XOR2_X1 U214 ( .A(n10), .B(n67), .Z(SUM[6]) );
  OAI21_X1 U215 ( .B1(n67), .B2(n65), .A(n66), .ZN(n64) );
  AOI21_X1 U216 ( .B1(n179), .B2(n171), .A(n169), .ZN(n21) );
  NAND2_X1 U217 ( .A1(n168), .A2(n25), .ZN(n2) );
  NAND2_X1 U218 ( .A1(n168), .A2(n170), .ZN(n20) );
  OAI21_X1 U219 ( .B1(n40), .B2(n36), .A(n37), .ZN(n35) );
  INV_X1 U220 ( .A(n172), .ZN(n94) );
  NOR2_X1 U221 ( .A1(A[13]), .A2(B[13]), .ZN(n27) );
  OAI21_X1 U222 ( .B1(n43), .B2(n55), .A(n44), .ZN(n42) );
  AOI21_X1 U223 ( .B1(n180), .B2(n51), .A(n173), .ZN(n44) );
  NAND2_X1 U224 ( .A1(n161), .A2(n181), .ZN(n43) );
  NAND2_X1 U225 ( .A1(A[15]), .A2(B[15]), .ZN(n18) );
  OAI21_X1 U226 ( .B1(n41), .B2(n162), .A(n40), .ZN(n38) );
  INV_X1 U227 ( .A(n39), .ZN(n95) );
  NOR2_X1 U228 ( .A1(n172), .A2(n39), .ZN(n34) );
  NAND2_X1 U229 ( .A1(n161), .A2(n48), .ZN(n6) );
  XNOR2_X1 U230 ( .A(n38), .B(n4), .ZN(SUM[12]) );
  XNOR2_X1 U231 ( .A(n19), .B(n1), .ZN(SUM[15]) );
  XNOR2_X1 U232 ( .A(n26), .B(n2), .ZN(SUM[14]) );
  XOR2_X1 U233 ( .A(n174), .B(n3), .Z(SUM[13]) );
  OAI21_X1 U234 ( .B1(n175), .B2(n27), .A(n28), .ZN(n26) );
  OAI21_X1 U235 ( .B1(n174), .B2(n20), .A(n21), .ZN(n19) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_5 ( clk, clear_acc, 
        data_out_x, data_out, data_out_w, data_out_b, wr_en_y, m_valid, 
        m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [3:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N27, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, n1, n2, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n87, n104, n113, n114, n115, n116, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n17), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n221), .CK(clk), .Q(n22) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n222), .CK(clk), .Q(n23) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n223), .CK(clk), .Q(n24) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n224), .CK(clk), .Q(n25) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n225), .CK(clk), .Q(n26) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n226), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n227), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n228), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n229), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n230), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n231), .CK(clk), .Q(n34) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n232), .CK(clk), .Q(n35) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n233), .CK(clk), .Q(n36) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n234), .CK(clk), .Q(n37) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n235), .CK(clk), .Q(n38) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n236), .CK(clk), .Q(n40) );
  DFF_X1 \f_reg[8]  ( .D(n80), .CK(clk), .Q(f[8]), .QN(n214) );
  DFF_X1 \f_reg[9]  ( .D(n79), .CK(clk), .Q(f[9]), .QN(n215) );
  DFF_X1 \f_reg[10]  ( .D(n78), .CK(clk), .Q(n50), .QN(n216) );
  DFF_X1 \f_reg[11]  ( .D(n77), .CK(clk), .Q(n48), .QN(n217) );
  DFF_X1 \f_reg[12]  ( .D(n1), .CK(clk), .Q(n47), .QN(n218) );
  DFF_X1 \f_reg[13]  ( .D(n76), .CK(clk), .Q(n45), .QN(n219) );
  DFF_X1 \f_reg[14]  ( .D(n7), .CK(clk), .Q(n44), .QN(n220) );
  DFF_X1 \f_reg[15]  ( .D(n6), .CK(clk), .Q(f[15]), .QN(n74) );
  DFF_X1 \data_out_reg[15]  ( .D(n114), .CK(clk), .Q(data_out[15]), .QN(n193)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n115), .CK(clk), .Q(data_out[14]), .QN(n192)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n116), .CK(clk), .Q(data_out[13]), .QN(n191)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n165), .CK(clk), .Q(data_out[12]), .QN(n190)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n166), .CK(clk), .Q(data_out[11]), .QN(n189)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n167), .CK(clk), .Q(data_out[10]), .QN(n188)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n168), .CK(clk), .Q(data_out[9]), .QN(n187) );
  DFF_X1 \data_out_reg[8]  ( .D(n169), .CK(clk), .Q(data_out[8]), .QN(n186) );
  DFF_X1 \data_out_reg[7]  ( .D(n170), .CK(clk), .Q(data_out[7]), .QN(n185) );
  DFF_X1 \data_out_reg[6]  ( .D(n171), .CK(clk), .Q(data_out[6]), .QN(n184) );
  DFF_X1 \data_out_reg[5]  ( .D(n172), .CK(clk), .Q(data_out[5]), .QN(n183) );
  DFF_X1 \data_out_reg[4]  ( .D(n173), .CK(clk), .Q(data_out[4]), .QN(n182) );
  DFF_X1 \data_out_reg[3]  ( .D(n174), .CK(clk), .Q(data_out[3]), .QN(n181) );
  DFF_X1 \data_out_reg[2]  ( .D(n175), .CK(clk), .Q(data_out[2]), .QN(n180) );
  DFF_X1 \data_out_reg[1]  ( .D(n176), .CK(clk), .Q(data_out[1]), .QN(n179) );
  DFF_X1 \data_out_reg[0]  ( .D(n177), .CK(clk), .Q(data_out[0]), .QN(n178) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_5_DW_mult_tc_1 mult_960 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_5_DW01_add_2 add_961 ( .A({n200, 
        n199, n198, n197, n196, n195, n209, n208, n207, n206, n205, n204, n203, 
        n202, n201, n194}), .B({f[15], n44, n45, n47, n48, n50, f[9:3], n58, 
        n60, n62}), .CI(1'b0), .SUM(adder) );
  DFF_X2 delay_reg ( .D(N27), .CK(clk), .Q(n14), .QN(n237) );
  DFF_X1 \f_reg[3]  ( .D(n85), .CK(clk), .Q(f[3]), .QN(n66) );
  DFF_X1 \f_reg[1]  ( .D(n104), .CK(clk), .Q(n60), .QN(n211) );
  DFF_X1 \f_reg[4]  ( .D(n84), .CK(clk), .Q(f[4]), .QN(n67) );
  DFF_X1 \f_reg[2]  ( .D(n87), .CK(clk), .Q(n58), .QN(n212) );
  DFF_X1 \f_reg[0]  ( .D(n113), .CK(clk), .Q(n62), .QN(n210) );
  DFF_X1 \f_reg[5]  ( .D(n83), .CK(clk), .Q(f[5]), .QN(n68) );
  DFF_X1 \f_reg[6]  ( .D(n82), .CK(clk), .Q(f[6]), .QN(n69) );
  DFF_X1 \f_reg[7]  ( .D(n81), .CK(clk), .Q(f[7]), .QN(n213) );
  AND2_X2 U3 ( .A1(n43), .A2(n18), .ZN(n15) );
  NAND3_X1 U4 ( .A1(n4), .A2(n2), .A3(n5), .ZN(n1) );
  MUX2_X2 U5 ( .A(n29), .B(N37), .S(n237), .Z(n208) );
  MUX2_X1 U6 ( .A(N39), .B(n27), .S(n14), .Z(n195) );
  NAND2_X1 U8 ( .A1(data_out_b[12]), .A2(n17), .ZN(n2) );
  NAND2_X1 U9 ( .A1(adder[12]), .A2(n15), .ZN(n4) );
  NAND2_X1 U10 ( .A1(n64), .A2(n47), .ZN(n5) );
  NAND3_X1 U11 ( .A1(n12), .A2(n11), .A3(n13), .ZN(n6) );
  NAND3_X1 U12 ( .A1(n9), .A2(n8), .A3(n10), .ZN(n7) );
  NAND2_X1 U13 ( .A1(data_out_b[14]), .A2(n17), .ZN(n8) );
  NAND2_X1 U14 ( .A1(adder[14]), .A2(n15), .ZN(n9) );
  NAND2_X1 U15 ( .A1(n64), .A2(n44), .ZN(n10) );
  MUX2_X2 U16 ( .A(N43), .B(n23), .S(n14), .Z(n199) );
  MUX2_X2 U17 ( .A(n26), .B(N40), .S(n237), .Z(n196) );
  MUX2_X2 U18 ( .A(n25), .B(N41), .S(n237), .Z(n197) );
  NAND2_X1 U19 ( .A1(data_out_b[15]), .A2(n17), .ZN(n11) );
  NAND2_X1 U20 ( .A1(adder[15]), .A2(n15), .ZN(n12) );
  NAND2_X1 U21 ( .A1(n64), .A2(f[15]), .ZN(n13) );
  INV_X2 U22 ( .A(n43), .ZN(n64) );
  MUX2_X2 U23 ( .A(N42), .B(n24), .S(n14), .Z(n198) );
  INV_X1 U24 ( .A(n18), .ZN(n17) );
  INV_X1 U25 ( .A(clear_acc), .ZN(n18) );
  NAND2_X1 U26 ( .A1(n16), .A2(N27), .ZN(n239) );
  OAI22_X1 U27 ( .A1(n181), .A2(n239), .B1(n66), .B2(n238), .ZN(n174) );
  OAI22_X1 U28 ( .A1(n182), .A2(n239), .B1(n67), .B2(n238), .ZN(n173) );
  OAI22_X1 U29 ( .A1(n183), .A2(n239), .B1(n68), .B2(n238), .ZN(n172) );
  OAI22_X1 U30 ( .A1(n184), .A2(n239), .B1(n69), .B2(n238), .ZN(n171) );
  OAI22_X1 U31 ( .A1(n185), .A2(n239), .B1(n213), .B2(n238), .ZN(n170) );
  OAI22_X1 U32 ( .A1(n186), .A2(n239), .B1(n214), .B2(n238), .ZN(n169) );
  OAI22_X1 U33 ( .A1(n187), .A2(n239), .B1(n215), .B2(n238), .ZN(n168) );
  INV_X1 U34 ( .A(n21), .ZN(n39) );
  INV_X1 U35 ( .A(wr_en_y), .ZN(n16) );
  AND2_X1 U36 ( .A1(sel[0]), .A2(sel[1]), .ZN(n20) );
  INV_X1 U37 ( .A(m_ready), .ZN(n19) );
  NAND2_X1 U38 ( .A1(m_valid), .A2(n19), .ZN(n41) );
  OAI211_X1 U39 ( .C1(sel[2]), .C2(n20), .A(sel[3]), .B(n41), .ZN(N27) );
  NAND2_X1 U40 ( .A1(clear_acc_delay), .A2(n237), .ZN(n21) );
  MUX2_X1 U41 ( .A(n22), .B(N44), .S(n39), .Z(n221) );
  MUX2_X1 U42 ( .A(n22), .B(N44), .S(n237), .Z(n200) );
  MUX2_X1 U43 ( .A(n23), .B(N43), .S(n39), .Z(n222) );
  MUX2_X1 U44 ( .A(n24), .B(N42), .S(n39), .Z(n223) );
  MUX2_X1 U45 ( .A(n25), .B(N41), .S(n39), .Z(n224) );
  MUX2_X1 U46 ( .A(n26), .B(N40), .S(n39), .Z(n225) );
  MUX2_X1 U47 ( .A(n27), .B(N39), .S(n39), .Z(n226) );
  MUX2_X1 U48 ( .A(n28), .B(N38), .S(n39), .Z(n227) );
  MUX2_X1 U49 ( .A(n28), .B(N38), .S(n237), .Z(n209) );
  MUX2_X1 U50 ( .A(n29), .B(N37), .S(n39), .Z(n228) );
  MUX2_X1 U51 ( .A(n32), .B(N36), .S(n39), .Z(n229) );
  MUX2_X1 U52 ( .A(n32), .B(N36), .S(n237), .Z(n207) );
  MUX2_X1 U53 ( .A(n33), .B(N35), .S(n39), .Z(n230) );
  MUX2_X1 U54 ( .A(n33), .B(N35), .S(n237), .Z(n206) );
  MUX2_X1 U55 ( .A(n34), .B(N34), .S(n39), .Z(n231) );
  MUX2_X1 U56 ( .A(n34), .B(N34), .S(n237), .Z(n205) );
  MUX2_X1 U57 ( .A(n35), .B(N33), .S(n39), .Z(n232) );
  MUX2_X1 U58 ( .A(n35), .B(N33), .S(n237), .Z(n204) );
  MUX2_X1 U59 ( .A(n36), .B(N32), .S(n39), .Z(n233) );
  MUX2_X1 U60 ( .A(n36), .B(N32), .S(n237), .Z(n203) );
  MUX2_X1 U61 ( .A(n37), .B(N31), .S(n39), .Z(n234) );
  MUX2_X1 U62 ( .A(n37), .B(N31), .S(n237), .Z(n202) );
  MUX2_X1 U63 ( .A(n38), .B(N30), .S(n39), .Z(n235) );
  MUX2_X1 U64 ( .A(n38), .B(N30), .S(n237), .Z(n201) );
  MUX2_X1 U65 ( .A(n40), .B(N29), .S(n39), .Z(n236) );
  MUX2_X1 U66 ( .A(n40), .B(N29), .S(n237), .Z(n194) );
  INV_X1 U67 ( .A(n41), .ZN(n42) );
  OAI21_X1 U68 ( .B1(n42), .B2(n14), .A(n18), .ZN(n43) );
  AOI222_X1 U69 ( .A1(data_out_b[13]), .A2(n17), .B1(adder[13]), .B2(n15), 
        .C1(n64), .C2(n45), .ZN(n46) );
  INV_X1 U70 ( .A(n46), .ZN(n76) );
  AOI222_X1 U71 ( .A1(data_out_b[11]), .A2(n17), .B1(adder[11]), .B2(n15), 
        .C1(n64), .C2(n48), .ZN(n49) );
  INV_X1 U72 ( .A(n49), .ZN(n77) );
  AOI222_X1 U73 ( .A1(data_out_b[10]), .A2(n17), .B1(adder[10]), .B2(n15), 
        .C1(n64), .C2(n50), .ZN(n51) );
  INV_X1 U74 ( .A(n51), .ZN(n78) );
  AOI222_X1 U75 ( .A1(data_out_b[8]), .A2(n17), .B1(adder[8]), .B2(n15), .C1(
        n64), .C2(f[8]), .ZN(n52) );
  INV_X1 U76 ( .A(n52), .ZN(n80) );
  AOI222_X1 U77 ( .A1(data_out_b[7]), .A2(n17), .B1(adder[7]), .B2(n15), .C1(
        n64), .C2(f[7]), .ZN(n53) );
  INV_X1 U78 ( .A(n53), .ZN(n81) );
  AOI222_X1 U79 ( .A1(data_out_b[6]), .A2(n17), .B1(adder[6]), .B2(n15), .C1(
        n64), .C2(f[6]), .ZN(n54) );
  INV_X1 U80 ( .A(n54), .ZN(n82) );
  AOI222_X1 U81 ( .A1(data_out_b[5]), .A2(n17), .B1(adder[5]), .B2(n15), .C1(
        n64), .C2(f[5]), .ZN(n55) );
  INV_X1 U82 ( .A(n55), .ZN(n83) );
  AOI222_X1 U83 ( .A1(data_out_b[4]), .A2(n17), .B1(adder[4]), .B2(n15), .C1(
        n64), .C2(f[4]), .ZN(n56) );
  INV_X1 U84 ( .A(n56), .ZN(n84) );
  AOI222_X1 U85 ( .A1(data_out_b[3]), .A2(n17), .B1(adder[3]), .B2(n15), .C1(
        n64), .C2(f[3]), .ZN(n57) );
  INV_X1 U86 ( .A(n57), .ZN(n85) );
  AOI222_X1 U87 ( .A1(data_out_b[2]), .A2(n17), .B1(adder[2]), .B2(n15), .C1(
        n64), .C2(n58), .ZN(n59) );
  INV_X1 U88 ( .A(n59), .ZN(n87) );
  AOI222_X1 U89 ( .A1(data_out_b[1]), .A2(n17), .B1(adder[1]), .B2(n15), .C1(
        n64), .C2(n60), .ZN(n61) );
  INV_X1 U90 ( .A(n61), .ZN(n104) );
  AOI222_X1 U91 ( .A1(data_out_b[0]), .A2(n17), .B1(adder[0]), .B2(n15), .C1(
        n64), .C2(n62), .ZN(n63) );
  INV_X1 U92 ( .A(n63), .ZN(n113) );
  AOI222_X1 U93 ( .A1(data_out_b[9]), .A2(n17), .B1(adder[9]), .B2(n15), .C1(
        n64), .C2(f[9]), .ZN(n65) );
  INV_X1 U94 ( .A(n65), .ZN(n79) );
  NOR4_X1 U95 ( .A1(n48), .A2(n47), .A3(n45), .A4(n44), .ZN(n73) );
  NOR4_X1 U96 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n50), .ZN(n72) );
  NAND4_X1 U97 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(n70) );
  NOR4_X1 U98 ( .A1(n70), .A2(n62), .A3(n60), .A4(n58), .ZN(n71) );
  NAND3_X1 U99 ( .A1(n73), .A2(n72), .A3(n71), .ZN(n75) );
  NAND3_X1 U100 ( .A1(wr_en_y), .A2(n75), .A3(n74), .ZN(n238) );
  OAI22_X1 U101 ( .A1(n178), .A2(n239), .B1(n210), .B2(n238), .ZN(n177) );
  OAI22_X1 U102 ( .A1(n179), .A2(n239), .B1(n211), .B2(n238), .ZN(n176) );
  OAI22_X1 U103 ( .A1(n180), .A2(n239), .B1(n212), .B2(n238), .ZN(n175) );
  OAI22_X1 U104 ( .A1(n188), .A2(n239), .B1(n216), .B2(n238), .ZN(n167) );
  OAI22_X1 U105 ( .A1(n189), .A2(n239), .B1(n217), .B2(n238), .ZN(n166) );
  OAI22_X1 U106 ( .A1(n190), .A2(n239), .B1(n218), .B2(n238), .ZN(n165) );
  OAI22_X1 U107 ( .A1(n191), .A2(n239), .B1(n219), .B2(n238), .ZN(n116) );
  OAI22_X1 U108 ( .A1(n192), .A2(n239), .B1(n220), .B2(n238), .ZN(n115) );
  OAI22_X1 U109 ( .A1(n193), .A2(n239), .B1(n74), .B2(n238), .ZN(n114) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_4_DW_mult_tc_1 ( a, b, 
        product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n9, n12, n13, n16, n18, n19, n23, n25, n27, n29, n31, n32,
         n34, n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n50, n52,
         n53, n54, n55, n56, n57, n58, n59, n62, n63, n64, n65, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n95, n96, n97, n98, n99, n101,
         n103, n104, n105, n107, n109, n111, n112, n113, n114, n115, n117,
         n119, n120, n122, n125, n127, n129, n135, n139, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n237, n245, n247, n249, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n418, n419, n420, n421, n422, n423, n424, n426, n427, n429,
         n431, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U148 ( .A(n265), .B(n144), .Z(n145) );
  XOR2_X1 U150 ( .A(n271), .B(n146), .Z(n147) );
  XOR2_X1 U152 ( .A(n301), .B(n148), .Z(n149) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U162 ( .A(n170), .B(n172), .CI(n179), .CO(n165), .S(n166) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n291), .CI(n263), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n317), .B(n252), .CO(n173), .S(n174) );
  FA_X1 U167 ( .A(n180), .B(n187), .CI(n178), .CO(n175), .S(n176) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U169 ( .A(n193), .B(n282), .CI(n191), .CO(n179), .S(n180) );
  FA_X1 U170 ( .A(n268), .B(n274), .CI(n292), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U172 ( .A(n197), .B(n190), .CI(n188), .CO(n185), .S(n186) );
  FA_X1 U173 ( .A(n199), .B(n201), .CI(n192), .CO(n187), .S(n188) );
  FA_X1 U174 ( .A(n275), .B(n293), .CI(n194), .CO(n189), .S(n190) );
  FA_X1 U175 ( .A(n305), .B(n283), .CI(n253), .CO(n191), .S(n192) );
  HA_X1 U176 ( .A(n319), .B(n269), .CO(n193), .S(n194) );
  FA_X1 U177 ( .A(n205), .B(n200), .CI(n198), .CO(n195), .S(n196) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U179 ( .A(n276), .B(n284), .CI(n294), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n320), .B(n270), .CI(n306), .CO(n201), .S(n202) );
  FA_X1 U181 ( .A(n208), .B(n213), .CI(n206), .CO(n203), .S(n204) );
  FA_X1 U182 ( .A(n210), .B(n307), .CI(n215), .CO(n205), .S(n206) );
  FA_X1 U183 ( .A(n254), .B(n285), .CI(n295), .CO(n207), .S(n208) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U185 ( .A(n216), .B(n219), .CI(n214), .CO(n211), .S(n212) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n322), .B(n278), .CI(n308), .CO(n215), .S(n216) );
  FA_X1 U188 ( .A(n225), .B(n222), .CI(n220), .CO(n217), .S(n218) );
  FA_X1 U189 ( .A(n255), .B(n309), .CI(n297), .CO(n219), .S(n220) );
  HA_X1 U190 ( .A(n287), .B(n323), .CO(n221), .S(n222) );
  FA_X1 U192 ( .A(n324), .B(n288), .CI(n310), .CO(n225), .S(n226) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  HA_X1 U194 ( .A(n311), .B(n325), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n326), .B(n300), .CI(n312), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  INV_X1 U414 ( .A(n13), .ZN(n490) );
  BUF_X1 U415 ( .A(n572), .Z(n491) );
  BUF_X1 U416 ( .A(n563), .Z(n492) );
  OR2_X2 U417 ( .A1(n545), .A2(n549), .ZN(n6) );
  AND2_X1 U418 ( .A1(n212), .A2(n217), .ZN(n547) );
  INV_X1 U419 ( .A(n547), .ZN(n95) );
  NOR2_X1 U420 ( .A1(n164), .A2(n175), .ZN(n75) );
  OR2_X1 U421 ( .A1(n329), .A2(n258), .ZN(n493) );
  XOR2_X1 U422 ( .A(n583), .B(a[14]), .Z(n41) );
  XNOR2_X1 U423 ( .A(n576), .B(a[6]), .ZN(n494) );
  BUF_X1 U424 ( .A(n83), .Z(n495) );
  INV_X1 U425 ( .A(n580), .ZN(n496) );
  XNOR2_X1 U426 ( .A(n576), .B(a[6]), .ZN(n546) );
  INV_X2 U427 ( .A(n583), .ZN(n582) );
  BUF_X2 U428 ( .A(n9), .Z(n563) );
  XOR2_X1 U429 ( .A(n577), .B(a[6]), .Z(n519) );
  BUF_X2 U430 ( .A(n19), .Z(n530) );
  INV_X1 U431 ( .A(n491), .ZN(n497) );
  XNOR2_X1 U432 ( .A(n166), .B(n498), .ZN(n164) );
  XNOR2_X1 U433 ( .A(n177), .B(n168), .ZN(n498) );
  OR2_X1 U434 ( .A1(n218), .A2(n223), .ZN(n499) );
  OR2_X1 U435 ( .A1(n176), .A2(n185), .ZN(n500) );
  NOR2_X1 U436 ( .A1(n186), .A2(n195), .ZN(n501) );
  NOR2_X1 U437 ( .A1(n186), .A2(n195), .ZN(n82) );
  INV_X1 U438 ( .A(n546), .ZN(n502) );
  INV_X1 U439 ( .A(n494), .ZN(n503) );
  NAND2_X1 U440 ( .A1(n228), .A2(n231), .ZN(n504) );
  INV_X1 U441 ( .A(n576), .ZN(n574) );
  INV_X2 U442 ( .A(n490), .ZN(n575) );
  INV_X1 U443 ( .A(n500), .ZN(n505) );
  NOR2_X1 U444 ( .A1(n176), .A2(n185), .ZN(n78) );
  INV_X1 U445 ( .A(n532), .ZN(n506) );
  INV_X1 U446 ( .A(n532), .ZN(n27) );
  NAND2_X1 U447 ( .A1(n166), .A2(n177), .ZN(n507) );
  NAND2_X1 U448 ( .A1(n166), .A2(n168), .ZN(n508) );
  NAND2_X1 U449 ( .A1(n177), .A2(n168), .ZN(n509) );
  NAND3_X1 U450 ( .A1(n507), .A2(n508), .A3(n509), .ZN(n163) );
  INV_X2 U451 ( .A(n581), .ZN(n523) );
  XOR2_X1 U452 ( .A(n25), .B(a[10]), .Z(n536) );
  OR2_X2 U453 ( .A1(n519), .A2(n494), .ZN(n510) );
  OR2_X1 U454 ( .A1(n519), .A2(n546), .ZN(n23) );
  CLKBUF_X1 U455 ( .A(n74), .Z(n511) );
  CLKBUF_X1 U456 ( .A(n12), .Z(n512) );
  AOI21_X1 U457 ( .B1(n557), .B2(n112), .A(n109), .ZN(n513) );
  NAND2_X1 U458 ( .A1(n431), .A2(n561), .ZN(n514) );
  NAND2_X1 U459 ( .A1(n431), .A2(n561), .ZN(n515) );
  NAND2_X1 U460 ( .A1(n431), .A2(n561), .ZN(n18) );
  CLKBUF_X1 U461 ( .A(n572), .Z(n516) );
  CLKBUF_X1 U462 ( .A(n534), .Z(n517) );
  AOI21_X1 U463 ( .B1(n88), .B2(n80), .A(n81), .ZN(n534) );
  CLKBUF_X1 U464 ( .A(n562), .Z(n518) );
  OR2_X2 U465 ( .A1(n545), .A2(n549), .ZN(n520) );
  OR2_X1 U466 ( .A1(n196), .A2(n203), .ZN(n521) );
  BUF_X2 U467 ( .A(n569), .Z(n522) );
  INV_X1 U468 ( .A(n581), .ZN(n580) );
  INV_X1 U469 ( .A(n1), .ZN(n524) );
  XOR2_X1 U470 ( .A(n573), .B(a[4]), .Z(n16) );
  BUF_X1 U471 ( .A(n37), .Z(n525) );
  OAI21_X1 U472 ( .B1(n91), .B2(n89), .A(n90), .ZN(n526) );
  OAI21_X1 U473 ( .B1(n513), .B2(n105), .A(n504), .ZN(n527) );
  OAI21_X1 U474 ( .B1(n91), .B2(n89), .A(n90), .ZN(n88) );
  XNOR2_X1 U475 ( .A(n579), .B(a[8]), .ZN(n429) );
  OR2_X2 U476 ( .A1(n528), .A2(n536), .ZN(n34) );
  XNOR2_X1 U477 ( .A(n580), .B(a[10]), .ZN(n528) );
  INV_X1 U478 ( .A(n249), .ZN(n569) );
  XNOR2_X1 U479 ( .A(n45), .B(n529), .ZN(product[12]) );
  AND2_X1 U480 ( .A1(n500), .A2(n79), .ZN(n529) );
  XNOR2_X1 U481 ( .A(a[2]), .B(n1), .ZN(n9) );
  INV_X1 U482 ( .A(n1), .ZN(n571) );
  XNOR2_X1 U483 ( .A(n226), .B(n531), .ZN(n224) );
  XNOR2_X1 U484 ( .A(n229), .B(n298), .ZN(n531) );
  XNOR2_X1 U485 ( .A(n577), .B(a[8]), .ZN(n532) );
  OR2_X1 U486 ( .A1(n228), .A2(n231), .ZN(n533) );
  CLKBUF_X1 U487 ( .A(n91), .Z(n535) );
  AOI21_X1 U488 ( .B1(n526), .B2(n80), .A(n81), .ZN(n45) );
  INV_X1 U489 ( .A(n536), .ZN(n32) );
  NAND2_X1 U490 ( .A1(n226), .A2(n229), .ZN(n537) );
  NAND2_X1 U491 ( .A1(n226), .A2(n298), .ZN(n538) );
  NAND2_X1 U492 ( .A1(n229), .A2(n298), .ZN(n539) );
  NAND3_X1 U493 ( .A1(n537), .A2(n538), .A3(n539), .ZN(n223) );
  AOI21_X1 U494 ( .B1(n553), .B2(n527), .A(n101), .ZN(n540) );
  OR2_X1 U495 ( .A1(n12), .A2(n388), .ZN(n541) );
  OR2_X1 U496 ( .A1(n387), .A2(n563), .ZN(n542) );
  NAND2_X1 U497 ( .A1(n541), .A2(n542), .ZN(n310) );
  INV_X2 U498 ( .A(n573), .ZN(n572) );
  BUF_X2 U499 ( .A(n16), .Z(n562) );
  NAND2_X1 U500 ( .A1(n429), .A2(n27), .ZN(n543) );
  NAND2_X1 U501 ( .A1(n429), .A2(n27), .ZN(n544) );
  NAND2_X1 U502 ( .A1(n429), .A2(n27), .ZN(n29) );
  XOR2_X1 U503 ( .A(n571), .B(n249), .Z(n545) );
  XNOR2_X1 U504 ( .A(n573), .B(a[2]), .ZN(n551) );
  OR2_X1 U505 ( .A1(n212), .A2(n217), .ZN(n548) );
  INV_X1 U506 ( .A(n571), .ZN(n570) );
  INV_X1 U507 ( .A(n569), .ZN(n549) );
  XNOR2_X1 U508 ( .A(n526), .B(n550), .ZN(product[10]) );
  NAND2_X1 U509 ( .A1(n521), .A2(n86), .ZN(n550) );
  OR2_X1 U510 ( .A1(n152), .A2(n163), .ZN(n552) );
  INV_X2 U511 ( .A(n579), .ZN(n578) );
  OR2_X1 U512 ( .A1(n328), .A2(n314), .ZN(n556) );
  OR2_X1 U513 ( .A1(n224), .A2(n227), .ZN(n553) );
  NAND2_X2 U514 ( .A1(n9), .A2(n551), .ZN(n12) );
  AOI21_X1 U515 ( .B1(n552), .B2(n511), .A(n67), .ZN(n65) );
  INV_X1 U516 ( .A(n69), .ZN(n67) );
  NAND2_X1 U517 ( .A1(n552), .A2(n69), .ZN(n47) );
  INV_X1 U518 ( .A(n73), .ZN(n71) );
  INV_X1 U519 ( .A(n74), .ZN(n72) );
  NAND2_X1 U520 ( .A1(n73), .A2(n552), .ZN(n64) );
  NOR2_X1 U521 ( .A1(n501), .A2(n85), .ZN(n80) );
  XNOR2_X1 U522 ( .A(n77), .B(n48), .ZN(product[13]) );
  NAND2_X1 U523 ( .A1(n125), .A2(n76), .ZN(n48) );
  INV_X1 U524 ( .A(n75), .ZN(n125) );
  NAND2_X1 U525 ( .A1(n129), .A2(n90), .ZN(n52) );
  INV_X1 U526 ( .A(n89), .ZN(n129) );
  NAND2_X1 U527 ( .A1(n548), .A2(n95), .ZN(n53) );
  OAI21_X1 U528 ( .B1(n75), .B2(n79), .A(n76), .ZN(n74) );
  NOR2_X1 U529 ( .A1(n75), .A2(n78), .ZN(n73) );
  XNOR2_X1 U530 ( .A(n84), .B(n50), .ZN(product[11]) );
  NAND2_X1 U531 ( .A1(n127), .A2(n495), .ZN(n50) );
  INV_X1 U532 ( .A(n501), .ZN(n127) );
  NAND2_X1 U533 ( .A1(n152), .A2(n163), .ZN(n69) );
  INV_X1 U534 ( .A(n103), .ZN(n101) );
  AOI21_X1 U535 ( .B1(n557), .B2(n112), .A(n109), .ZN(n107) );
  INV_X1 U536 ( .A(n111), .ZN(n109) );
  OAI21_X1 U537 ( .B1(n113), .B2(n115), .A(n114), .ZN(n112) );
  NAND2_X1 U538 ( .A1(n499), .A2(n98), .ZN(n54) );
  NOR2_X1 U539 ( .A1(n196), .A2(n203), .ZN(n85) );
  NAND2_X1 U540 ( .A1(n553), .A2(n103), .ZN(n55) );
  NAND2_X1 U541 ( .A1(n557), .A2(n111), .ZN(n57) );
  OAI21_X1 U542 ( .B1(n105), .B2(n107), .A(n504), .ZN(n104) );
  AOI21_X1 U543 ( .B1(n556), .B2(n120), .A(n117), .ZN(n115) );
  INV_X1 U544 ( .A(n119), .ZN(n117) );
  INV_X1 U545 ( .A(n122), .ZN(n120) );
  NAND2_X1 U546 ( .A1(n176), .A2(n185), .ZN(n79) );
  NAND2_X1 U547 ( .A1(n164), .A2(n175), .ZN(n76) );
  NAND2_X1 U548 ( .A1(n196), .A2(n203), .ZN(n86) );
  NAND2_X1 U549 ( .A1(n186), .A2(n195), .ZN(n83) );
  NAND2_X1 U550 ( .A1(n204), .A2(n211), .ZN(n90) );
  NAND2_X1 U551 ( .A1(n135), .A2(n114), .ZN(n58) );
  INV_X1 U552 ( .A(n113), .ZN(n135) );
  XNOR2_X1 U553 ( .A(n59), .B(n120), .ZN(product[2]) );
  NAND2_X1 U554 ( .A1(n556), .A2(n119), .ZN(n59) );
  NAND2_X1 U555 ( .A1(n533), .A2(n504), .ZN(n56) );
  AND2_X1 U556 ( .A1(n493), .A2(n122), .ZN(product[1]) );
  NAND2_X1 U557 ( .A1(n328), .A2(n314), .ZN(n119) );
  NOR2_X1 U558 ( .A1(n228), .A2(n231), .ZN(n105) );
  NOR2_X1 U559 ( .A1(n234), .A2(n257), .ZN(n113) );
  OR2_X1 U560 ( .A1(n151), .A2(n139), .ZN(n555) );
  XNOR2_X1 U561 ( .A(n63), .B(n46), .ZN(product[15]) );
  NAND2_X1 U562 ( .A1(n555), .A2(n62), .ZN(n46) );
  NOR2_X1 U563 ( .A1(n218), .A2(n223), .ZN(n97) );
  NAND2_X1 U564 ( .A1(n218), .A2(n223), .ZN(n98) );
  OR2_X1 U565 ( .A1(n232), .A2(n233), .ZN(n557) );
  INV_X1 U566 ( .A(n37), .ZN(n237) );
  NAND2_X1 U567 ( .A1(n224), .A2(n227), .ZN(n103) );
  INV_X1 U568 ( .A(n41), .ZN(n235) );
  XNOR2_X1 U569 ( .A(n523), .B(a[12]), .ZN(n37) );
  OR2_X1 U570 ( .A1(n567), .A2(n497), .ZN(n392) );
  XNOR2_X1 U571 ( .A(n530), .B(n567), .ZN(n363) );
  XNOR2_X1 U572 ( .A(n578), .B(n567), .ZN(n352) );
  AND2_X1 U573 ( .A1(n532), .A2(n568), .ZN(n278) );
  XNOR2_X1 U574 ( .A(n575), .B(n567), .ZN(n376) );
  XNOR2_X1 U575 ( .A(n155), .B(n558), .ZN(n139) );
  XNOR2_X1 U576 ( .A(n153), .B(n141), .ZN(n558) );
  XNOR2_X1 U577 ( .A(n157), .B(n559), .ZN(n141) );
  XNOR2_X1 U578 ( .A(n145), .B(n143), .ZN(n559) );
  OAI22_X1 U579 ( .A1(n39), .A2(n336), .B1(n525), .B2(n335), .ZN(n263) );
  OAI22_X1 U580 ( .A1(n39), .A2(n583), .B1(n337), .B2(n525), .ZN(n252) );
  OR2_X1 U581 ( .A1(n567), .A2(n583), .ZN(n337) );
  OAI22_X1 U582 ( .A1(n42), .A2(n585), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U583 ( .A1(n567), .A2(n585), .ZN(n332) );
  XNOR2_X1 U584 ( .A(n523), .B(n567), .ZN(n343) );
  AND2_X1 U585 ( .A1(n568), .A2(n245), .ZN(n300) );
  XNOR2_X1 U586 ( .A(n159), .B(n560), .ZN(n142) );
  XNOR2_X1 U587 ( .A(n315), .B(n261), .ZN(n560) );
  XNOR2_X1 U588 ( .A(n582), .B(n567), .ZN(n336) );
  NAND2_X1 U589 ( .A1(n427), .A2(n37), .ZN(n39) );
  XOR2_X1 U590 ( .A(n582), .B(a[12]), .Z(n427) );
  AND2_X1 U591 ( .A1(n568), .A2(n237), .ZN(n264) );
  AND2_X1 U592 ( .A1(n568), .A2(n494), .ZN(n288) );
  AND2_X1 U593 ( .A1(n568), .A2(n536), .ZN(n270) );
  AND2_X1 U594 ( .A1(n568), .A2(n235), .ZN(n260) );
  OAI22_X1 U595 ( .A1(n39), .A2(n335), .B1(n525), .B2(n334), .ZN(n262) );
  INV_X1 U596 ( .A(n25), .ZN(n579) );
  INV_X1 U597 ( .A(n13), .ZN(n576) );
  NAND2_X1 U598 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U599 ( .A(n584), .B(a[14]), .Z(n426) );
  INV_X1 U600 ( .A(n7), .ZN(n573) );
  AND2_X1 U601 ( .A1(n568), .A2(n247), .ZN(n314) );
  AND2_X1 U602 ( .A1(n568), .A2(n549), .ZN(product[0]) );
  OR2_X1 U603 ( .A1(n567), .A2(n490), .ZN(n377) );
  OR2_X1 U604 ( .A1(n567), .A2(n577), .ZN(n364) );
  OR2_X1 U605 ( .A1(n567), .A2(n579), .ZN(n353) );
  OR2_X1 U606 ( .A1(n567), .A2(n496), .ZN(n344) );
  XNOR2_X1 U607 ( .A(n530), .B(b[9]), .ZN(n354) );
  OAI22_X1 U608 ( .A1(n39), .A2(n334), .B1(n525), .B2(n333), .ZN(n261) );
  XNOR2_X1 U609 ( .A(n582), .B(n422), .ZN(n333) );
  XNOR2_X1 U610 ( .A(n575), .B(b[11]), .ZN(n365) );
  XNOR2_X1 U611 ( .A(n582), .B(n424), .ZN(n335) );
  XNOR2_X1 U612 ( .A(n582), .B(n423), .ZN(n334) );
  OAI22_X1 U613 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U614 ( .A(n584), .B(n424), .ZN(n330) );
  XNOR2_X1 U615 ( .A(n584), .B(n567), .ZN(n331) );
  XNOR2_X1 U616 ( .A(n523), .B(n420), .ZN(n338) );
  XNOR2_X1 U617 ( .A(n578), .B(n418), .ZN(n345) );
  XNOR2_X1 U618 ( .A(n516), .B(b[13]), .ZN(n378) );
  XNOR2_X1 U619 ( .A(n530), .B(n424), .ZN(n362) );
  XNOR2_X1 U620 ( .A(n523), .B(n424), .ZN(n342) );
  XNOR2_X1 U621 ( .A(n578), .B(n424), .ZN(n351) );
  XNOR2_X1 U622 ( .A(n523), .B(n423), .ZN(n341) );
  XNOR2_X1 U623 ( .A(n523), .B(n422), .ZN(n340) );
  XNOR2_X1 U624 ( .A(n523), .B(n421), .ZN(n339) );
  XNOR2_X1 U625 ( .A(n572), .B(n418), .ZN(n384) );
  XNOR2_X1 U626 ( .A(n572), .B(n419), .ZN(n385) );
  XNOR2_X1 U627 ( .A(n516), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U628 ( .A(n491), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U629 ( .A(n572), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U630 ( .A(n572), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U631 ( .A(n516), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U632 ( .A(n575), .B(n418), .ZN(n369) );
  XNOR2_X1 U633 ( .A(n575), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U634 ( .A(n575), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U635 ( .A(n575), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U636 ( .A(n530), .B(n423), .ZN(n361) );
  XNOR2_X1 U637 ( .A(n530), .B(n422), .ZN(n360) );
  XNOR2_X1 U638 ( .A(n578), .B(n423), .ZN(n350) );
  XNOR2_X1 U639 ( .A(n578), .B(n422), .ZN(n349) );
  XNOR2_X1 U640 ( .A(n530), .B(n420), .ZN(n358) );
  XNOR2_X1 U641 ( .A(n578), .B(n421), .ZN(n348) );
  XNOR2_X1 U642 ( .A(n530), .B(n421), .ZN(n359) );
  XNOR2_X1 U643 ( .A(n578), .B(n420), .ZN(n347) );
  XNOR2_X1 U644 ( .A(n530), .B(n418), .ZN(n356) );
  XNOR2_X1 U645 ( .A(n565), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U646 ( .A(n564), .B(b[11]), .ZN(n397) );
  XNOR2_X1 U647 ( .A(n564), .B(b[14]), .ZN(n394) );
  XNOR2_X1 U648 ( .A(n530), .B(n419), .ZN(n357) );
  XNOR2_X1 U649 ( .A(n578), .B(n419), .ZN(n346) );
  XNOR2_X1 U650 ( .A(n530), .B(b[8]), .ZN(n355) );
  XNOR2_X1 U651 ( .A(n570), .B(b[13]), .ZN(n395) );
  BUF_X1 U652 ( .A(n43), .Z(n568) );
  XNOR2_X1 U653 ( .A(n570), .B(b[15]), .ZN(n393) );
  CLKBUF_X1 U654 ( .A(n16), .Z(n561) );
  XNOR2_X1 U655 ( .A(n70), .B(n47), .ZN(product[14]) );
  OAI22_X1 U656 ( .A1(n34), .A2(n339), .B1(n338), .B2(n32), .ZN(n265) );
  OAI22_X1 U657 ( .A1(n34), .A2(n340), .B1(n339), .B2(n32), .ZN(n266) );
  OAI22_X1 U658 ( .A1(n34), .A2(n342), .B1(n341), .B2(n32), .ZN(n268) );
  OAI22_X1 U659 ( .A1(n34), .A2(n343), .B1(n342), .B2(n32), .ZN(n269) );
  OAI22_X1 U660 ( .A1(n34), .A2(n341), .B1(n340), .B2(n32), .ZN(n267) );
  OAI22_X1 U661 ( .A1(n34), .A2(n496), .B1(n344), .B2(n32), .ZN(n253) );
  INV_X1 U662 ( .A(n19), .ZN(n577) );
  OR2_X1 U663 ( .A1(n571), .A2(n567), .ZN(n409) );
  INV_X1 U664 ( .A(n524), .ZN(n564) );
  INV_X1 U665 ( .A(n524), .ZN(n565) );
  NAND2_X1 U666 ( .A1(n232), .A2(n233), .ZN(n111) );
  OAI22_X1 U667 ( .A1(n510), .A2(n358), .B1(n357), .B2(n502), .ZN(n282) );
  OAI22_X1 U668 ( .A1(n510), .A2(n362), .B1(n361), .B2(n503), .ZN(n286) );
  OAI22_X1 U669 ( .A1(n510), .A2(n360), .B1(n359), .B2(n502), .ZN(n284) );
  OAI22_X1 U670 ( .A1(n510), .A2(n356), .B1(n355), .B2(n503), .ZN(n280) );
  OAI22_X1 U671 ( .A1(n510), .A2(n577), .B1(n364), .B2(n503), .ZN(n255) );
  OAI22_X1 U672 ( .A1(n510), .A2(n357), .B1(n356), .B2(n502), .ZN(n281) );
  OAI22_X1 U673 ( .A1(n23), .A2(n363), .B1(n502), .B2(n362), .ZN(n287) );
  OAI22_X1 U674 ( .A1(n510), .A2(n361), .B1(n360), .B2(n503), .ZN(n285) );
  OAI22_X1 U675 ( .A1(n23), .A2(n359), .B1(n358), .B2(n502), .ZN(n283) );
  OAI22_X1 U676 ( .A1(n510), .A2(n355), .B1(n354), .B2(n502), .ZN(n279) );
  NOR2_X1 U677 ( .A1(n204), .A2(n211), .ZN(n89) );
  OAI22_X1 U678 ( .A1(n29), .A2(n350), .B1(n349), .B2(n506), .ZN(n275) );
  OAI22_X1 U679 ( .A1(n544), .A2(n346), .B1(n345), .B2(n506), .ZN(n271) );
  OAI22_X1 U680 ( .A1(n544), .A2(n351), .B1(n350), .B2(n506), .ZN(n276) );
  OAI22_X1 U681 ( .A1(n29), .A2(n347), .B1(n346), .B2(n506), .ZN(n272) );
  OAI22_X1 U682 ( .A1(n544), .A2(n348), .B1(n347), .B2(n506), .ZN(n273) );
  OAI22_X1 U683 ( .A1(n29), .A2(n349), .B1(n348), .B2(n506), .ZN(n274) );
  OAI22_X1 U684 ( .A1(n543), .A2(n579), .B1(n353), .B2(n506), .ZN(n254) );
  OAI22_X1 U685 ( .A1(n543), .A2(n352), .B1(n351), .B2(n506), .ZN(n277) );
  XNOR2_X1 U686 ( .A(n572), .B(n420), .ZN(n386) );
  XNOR2_X1 U687 ( .A(n491), .B(n567), .ZN(n391) );
  XNOR2_X1 U688 ( .A(n572), .B(n422), .ZN(n388) );
  XNOR2_X1 U689 ( .A(n572), .B(n424), .ZN(n390) );
  XNOR2_X1 U690 ( .A(n572), .B(n421), .ZN(n387) );
  XNOR2_X1 U691 ( .A(n572), .B(n423), .ZN(n389) );
  CLKBUF_X1 U692 ( .A(n96), .Z(n566) );
  XNOR2_X1 U693 ( .A(n575), .B(n424), .ZN(n375) );
  XNOR2_X1 U694 ( .A(n575), .B(n419), .ZN(n370) );
  XNOR2_X1 U695 ( .A(n575), .B(n420), .ZN(n371) );
  XNOR2_X1 U696 ( .A(n575), .B(n423), .ZN(n374) );
  XNOR2_X1 U697 ( .A(n575), .B(n421), .ZN(n372) );
  XNOR2_X1 U698 ( .A(n574), .B(n422), .ZN(n373) );
  XOR2_X1 U699 ( .A(n574), .B(a[4]), .Z(n431) );
  OAI21_X1 U700 ( .B1(n99), .B2(n97), .A(n98), .ZN(n96) );
  XNOR2_X1 U701 ( .A(n55), .B(n527), .ZN(product[6]) );
  AOI21_X1 U702 ( .B1(n104), .B2(n553), .A(n101), .ZN(n99) );
  OAI21_X1 U703 ( .B1(n82), .B2(n86), .A(n83), .ZN(n81) );
  OAI21_X1 U704 ( .B1(n87), .B2(n85), .A(n86), .ZN(n84) );
  XNOR2_X1 U705 ( .A(n565), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U706 ( .A(n570), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U707 ( .A(n564), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U708 ( .A(n565), .B(n418), .ZN(n401) );
  XNOR2_X1 U709 ( .A(n565), .B(n567), .ZN(n408) );
  XNOR2_X1 U710 ( .A(n570), .B(n421), .ZN(n404) );
  XNOR2_X1 U711 ( .A(n564), .B(n422), .ZN(n405) );
  XNOR2_X1 U712 ( .A(n565), .B(n420), .ZN(n403) );
  XNOR2_X1 U713 ( .A(n570), .B(n419), .ZN(n402) );
  XNOR2_X1 U714 ( .A(n564), .B(n424), .ZN(n407) );
  XNOR2_X1 U715 ( .A(n565), .B(n423), .ZN(n406) );
  NAND2_X1 U716 ( .A1(n151), .A2(n139), .ZN(n62) );
  OAI22_X1 U717 ( .A1(n514), .A2(n367), .B1(n366), .B2(n518), .ZN(n290) );
  OAI22_X1 U718 ( .A1(n515), .A2(n370), .B1(n369), .B2(n518), .ZN(n293) );
  OAI22_X1 U719 ( .A1(n18), .A2(n368), .B1(n367), .B2(n562), .ZN(n291) );
  OAI22_X1 U720 ( .A1(n514), .A2(n375), .B1(n374), .B2(n518), .ZN(n298) );
  OAI22_X1 U721 ( .A1(n18), .A2(n369), .B1(n368), .B2(n562), .ZN(n292) );
  OAI22_X1 U722 ( .A1(n514), .A2(n373), .B1(n372), .B2(n562), .ZN(n296) );
  OAI22_X1 U723 ( .A1(n514), .A2(n371), .B1(n370), .B2(n562), .ZN(n294) );
  OAI22_X1 U724 ( .A1(n515), .A2(n372), .B1(n371), .B2(n562), .ZN(n295) );
  OAI22_X1 U725 ( .A1(n18), .A2(n374), .B1(n373), .B2(n562), .ZN(n297) );
  OAI22_X1 U726 ( .A1(n514), .A2(n490), .B1(n377), .B2(n562), .ZN(n256) );
  OAI22_X1 U727 ( .A1(n515), .A2(n376), .B1(n375), .B2(n562), .ZN(n299) );
  OAI22_X1 U728 ( .A1(n515), .A2(n366), .B1(n365), .B2(n562), .ZN(n289) );
  INV_X1 U729 ( .A(n562), .ZN(n245) );
  XOR2_X1 U730 ( .A(n56), .B(n513), .Z(product[5]) );
  XNOR2_X1 U731 ( .A(n57), .B(n112), .ZN(product[4]) );
  INV_X1 U732 ( .A(n88), .ZN(n87) );
  OAI21_X1 U733 ( .B1(n64), .B2(n517), .A(n65), .ZN(n63) );
  OAI21_X1 U734 ( .B1(n534), .B2(n71), .A(n72), .ZN(n70) );
  OAI21_X1 U735 ( .B1(n534), .B2(n505), .A(n79), .ZN(n77) );
  XOR2_X1 U736 ( .A(n535), .B(n52), .Z(product[9]) );
  XNOR2_X1 U737 ( .A(n566), .B(n53), .ZN(product[8]) );
  AOI21_X1 U738 ( .B1(n96), .B2(n548), .A(n547), .ZN(n91) );
  XOR2_X1 U739 ( .A(n58), .B(n115), .Z(product[3]) );
  OAI22_X1 U740 ( .A1(n520), .A2(n395), .B1(n394), .B2(n522), .ZN(n316) );
  OAI22_X1 U741 ( .A1(n520), .A2(n394), .B1(n393), .B2(n522), .ZN(n315) );
  OAI22_X1 U742 ( .A1(n520), .A2(n396), .B1(n395), .B2(n522), .ZN(n317) );
  OAI22_X1 U743 ( .A1(n520), .A2(n397), .B1(n396), .B2(n522), .ZN(n318) );
  OAI22_X1 U744 ( .A1(n520), .A2(n398), .B1(n397), .B2(n522), .ZN(n319) );
  OAI22_X1 U745 ( .A1(n520), .A2(n400), .B1(n399), .B2(n522), .ZN(n321) );
  OAI22_X1 U746 ( .A1(n6), .A2(n399), .B1(n398), .B2(n522), .ZN(n320) );
  OAI22_X1 U747 ( .A1(n6), .A2(n401), .B1(n400), .B2(n522), .ZN(n322) );
  OAI22_X1 U748 ( .A1(n6), .A2(n402), .B1(n401), .B2(n522), .ZN(n323) );
  NAND2_X1 U749 ( .A1(n329), .A2(n258), .ZN(n122) );
  OAI22_X1 U750 ( .A1(n6), .A2(n404), .B1(n403), .B2(n569), .ZN(n325) );
  OAI22_X1 U751 ( .A1(n6), .A2(n403), .B1(n402), .B2(n522), .ZN(n324) );
  OAI22_X1 U752 ( .A1(n520), .A2(n406), .B1(n405), .B2(n522), .ZN(n327) );
  OAI22_X1 U753 ( .A1(n520), .A2(n405), .B1(n404), .B2(n522), .ZN(n326) );
  OAI22_X1 U754 ( .A1(n520), .A2(n407), .B1(n406), .B2(n522), .ZN(n328) );
  OAI22_X1 U755 ( .A1(n520), .A2(n408), .B1(n407), .B2(n522), .ZN(n329) );
  OAI22_X1 U756 ( .A1(n520), .A2(n524), .B1(n409), .B2(n522), .ZN(n258) );
  XOR2_X1 U757 ( .A(n540), .B(n54), .Z(product[7]) );
  OAI22_X1 U758 ( .A1(n512), .A2(n379), .B1(n378), .B2(n492), .ZN(n301) );
  OAI22_X1 U759 ( .A1(n512), .A2(n380), .B1(n379), .B2(n563), .ZN(n302) );
  OAI22_X1 U760 ( .A1(n512), .A2(n385), .B1(n384), .B2(n492), .ZN(n307) );
  OAI22_X1 U761 ( .A1(n12), .A2(n382), .B1(n381), .B2(n563), .ZN(n304) );
  OAI22_X1 U762 ( .A1(n12), .A2(n381), .B1(n380), .B2(n563), .ZN(n303) );
  NAND2_X1 U763 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U764 ( .A1(n12), .A2(n383), .B1(n382), .B2(n563), .ZN(n305) );
  OAI22_X1 U765 ( .A1(n12), .A2(n384), .B1(n383), .B2(n563), .ZN(n306) );
  OAI22_X1 U766 ( .A1(n12), .A2(n386), .B1(n385), .B2(n563), .ZN(n308) );
  OAI22_X1 U767 ( .A1(n12), .A2(n387), .B1(n386), .B2(n563), .ZN(n309) );
  OAI22_X1 U768 ( .A1(n12), .A2(n497), .B1(n392), .B2(n563), .ZN(n257) );
  OAI22_X1 U769 ( .A1(n12), .A2(n389), .B1(n388), .B2(n563), .ZN(n311) );
  OAI22_X1 U770 ( .A1(n12), .A2(n390), .B1(n389), .B2(n563), .ZN(n312) );
  INV_X1 U771 ( .A(n563), .ZN(n247) );
  OAI22_X1 U772 ( .A1(n12), .A2(n391), .B1(n390), .B2(n563), .ZN(n313) );
  BUF_X4 U773 ( .A(n43), .Z(n567) );
  INV_X1 U774 ( .A(n31), .ZN(n581) );
  INV_X1 U775 ( .A(n36), .ZN(n583) );
  INV_X1 U776 ( .A(n585), .ZN(n584) );
  INV_X1 U777 ( .A(n40), .ZN(n585) );
  XOR2_X1 U778 ( .A(n259), .B(n251), .Z(n148) );
  XOR2_X1 U779 ( .A(n289), .B(n279), .Z(n146) );
  XOR2_X1 U780 ( .A(n149), .B(n147), .Z(n144) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_4_DW01_add_2 ( A, B, CI, SUM, 
        CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n18,
         n19, n20, n21, n23, n25, n26, n27, n28, n30, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n46, n48, n49, n51, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n71,
         n72, n73, n74, n75, n77, n79, n80, n81, n82, n83, n85, n87, n88, n90,
         n93, n94, n98, n99, n100, n102, n104, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179;

  AND2_X1 U126 ( .A1(n174), .A2(n90), .ZN(SUM[0]) );
  OR2_X1 U127 ( .A1(A[15]), .A2(B[15]), .ZN(n162) );
  XNOR2_X1 U128 ( .A(n41), .B(n163), .ZN(SUM[11]) );
  AND2_X1 U129 ( .A1(n172), .A2(n166), .ZN(n163) );
  BUF_X1 U130 ( .A(n27), .Z(n164) );
  OR2_X1 U131 ( .A1(A[14]), .A2(B[14]), .ZN(n175) );
  OR2_X1 U132 ( .A1(A[10]), .A2(B[10]), .ZN(n165) );
  NAND2_X1 U133 ( .A1(A[11]), .A2(B[11]), .ZN(n166) );
  NOR2_X1 U134 ( .A1(A[8]), .A2(B[8]), .ZN(n167) );
  NOR2_X1 U135 ( .A1(A[8]), .A2(B[8]), .ZN(n58) );
  AOI21_X1 U136 ( .B1(n165), .B2(n51), .A(n46), .ZN(n168) );
  OAI21_X1 U137 ( .B1(n55), .B2(n43), .A(n168), .ZN(n169) );
  NOR2_X1 U138 ( .A1(A[12]), .A2(B[12]), .ZN(n170) );
  NOR2_X1 U139 ( .A1(A[12]), .A2(B[12]), .ZN(n36) );
  AOI21_X1 U140 ( .B1(n56), .B2(n64), .A(n57), .ZN(n171) );
  OR2_X1 U141 ( .A1(A[11]), .A2(B[11]), .ZN(n172) );
  AOI21_X1 U142 ( .B1(n42), .B2(n34), .A(n35), .ZN(n173) );
  AOI21_X1 U143 ( .B1(n169), .B2(n34), .A(n35), .ZN(n33) );
  NOR2_X1 U144 ( .A1(A[7]), .A2(B[7]), .ZN(n61) );
  OR2_X1 U145 ( .A1(A[9]), .A2(B[9]), .ZN(n177) );
  OR2_X1 U146 ( .A1(A[0]), .A2(B[0]), .ZN(n174) );
  INV_X1 U147 ( .A(n64), .ZN(n63) );
  INV_X1 U148 ( .A(n171), .ZN(n54) );
  INV_X1 U149 ( .A(n42), .ZN(n41) );
  INV_X1 U150 ( .A(n71), .ZN(n69) );
  AOI21_X1 U151 ( .B1(n178), .B2(n88), .A(n85), .ZN(n83) );
  INV_X1 U152 ( .A(n87), .ZN(n85) );
  AOI21_X1 U153 ( .B1(n56), .B2(n64), .A(n57), .ZN(n55) );
  AOI21_X1 U154 ( .B1(n176), .B2(n80), .A(n77), .ZN(n75) );
  INV_X1 U155 ( .A(n79), .ZN(n77) );
  NAND2_X1 U156 ( .A1(n175), .A2(n93), .ZN(n20) );
  INV_X1 U157 ( .A(n28), .ZN(n30) );
  OAI21_X1 U158 ( .B1(n83), .B2(n81), .A(n82), .ZN(n80) );
  AOI21_X1 U159 ( .B1(n54), .B2(n177), .A(n51), .ZN(n49) );
  NAND2_X1 U160 ( .A1(n98), .A2(n59), .ZN(n8) );
  INV_X1 U161 ( .A(n90), .ZN(n88) );
  OAI21_X1 U162 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  INV_X1 U163 ( .A(n53), .ZN(n51) );
  NAND2_X1 U164 ( .A1(n99), .A2(n62), .ZN(n9) );
  INV_X1 U165 ( .A(n61), .ZN(n99) );
  NAND2_X1 U166 ( .A1(n177), .A2(n53), .ZN(n7) );
  NAND2_X1 U167 ( .A1(n104), .A2(n82), .ZN(n14) );
  INV_X1 U168 ( .A(n81), .ZN(n104) );
  NAND2_X1 U169 ( .A1(n176), .A2(n79), .ZN(n13) );
  NAND2_X1 U170 ( .A1(n179), .A2(n71), .ZN(n11) );
  NAND2_X1 U171 ( .A1(n178), .A2(n87), .ZN(n15) );
  INV_X1 U172 ( .A(n25), .ZN(n23) );
  AOI21_X1 U173 ( .B1(n165), .B2(n51), .A(n46), .ZN(n44) );
  INV_X1 U174 ( .A(n48), .ZN(n46) );
  NAND2_X1 U175 ( .A1(n100), .A2(n66), .ZN(n10) );
  INV_X1 U176 ( .A(n65), .ZN(n100) );
  NAND2_X1 U177 ( .A1(n102), .A2(n74), .ZN(n12) );
  INV_X1 U178 ( .A(n73), .ZN(n102) );
  NAND2_X1 U179 ( .A1(n175), .A2(n25), .ZN(n2) );
  XNOR2_X1 U180 ( .A(n38), .B(n4), .ZN(SUM[12]) );
  NAND2_X1 U181 ( .A1(n94), .A2(n37), .ZN(n4) );
  XNOR2_X1 U182 ( .A(n54), .B(n7), .ZN(SUM[9]) );
  XOR2_X1 U183 ( .A(n63), .B(n9), .Z(SUM[7]) );
  XNOR2_X1 U184 ( .A(n11), .B(n72), .ZN(SUM[5]) );
  XNOR2_X1 U185 ( .A(n13), .B(n80), .ZN(SUM[3]) );
  XOR2_X1 U186 ( .A(n14), .B(n83), .Z(SUM[2]) );
  XNOR2_X1 U187 ( .A(n15), .B(n88), .ZN(SUM[1]) );
  NOR2_X1 U188 ( .A1(A[11]), .A2(B[11]), .ZN(n39) );
  OR2_X1 U189 ( .A1(A[3]), .A2(B[3]), .ZN(n176) );
  NAND2_X1 U190 ( .A1(n93), .A2(n28), .ZN(n3) );
  NOR2_X1 U191 ( .A1(A[2]), .A2(B[2]), .ZN(n81) );
  XOR2_X1 U192 ( .A(n49), .B(n6), .Z(SUM[10]) );
  NAND2_X1 U193 ( .A1(A[11]), .A2(B[11]), .ZN(n40) );
  OR2_X1 U194 ( .A1(A[1]), .A2(B[1]), .ZN(n178) );
  NAND2_X1 U195 ( .A1(A[12]), .A2(B[12]), .ZN(n37) );
  XNOR2_X1 U196 ( .A(n60), .B(n8), .ZN(SUM[8]) );
  NOR2_X1 U197 ( .A1(A[6]), .A2(B[6]), .ZN(n65) );
  NOR2_X1 U198 ( .A1(A[4]), .A2(B[4]), .ZN(n73) );
  NAND2_X1 U199 ( .A1(A[7]), .A2(B[7]), .ZN(n62) );
  NAND2_X1 U200 ( .A1(A[2]), .A2(B[2]), .ZN(n82) );
  NAND2_X1 U201 ( .A1(A[9]), .A2(B[9]), .ZN(n53) );
  NAND2_X1 U202 ( .A1(A[5]), .A2(B[5]), .ZN(n71) );
  NAND2_X1 U203 ( .A1(A[1]), .A2(B[1]), .ZN(n87) );
  NAND2_X1 U204 ( .A1(A[0]), .A2(B[0]), .ZN(n90) );
  OR2_X1 U205 ( .A1(A[5]), .A2(B[5]), .ZN(n179) );
  NAND2_X1 U206 ( .A1(A[6]), .A2(B[6]), .ZN(n66) );
  NAND2_X1 U207 ( .A1(A[4]), .A2(B[4]), .ZN(n74) );
  NAND2_X1 U208 ( .A1(A[3]), .A2(B[3]), .ZN(n79) );
  NAND2_X1 U209 ( .A1(n162), .A2(n18), .ZN(n1) );
  INV_X1 U210 ( .A(n27), .ZN(n93) );
  NAND2_X1 U211 ( .A1(A[15]), .A2(B[15]), .ZN(n18) );
  OAI21_X1 U212 ( .B1(n41), .B2(n39), .A(n166), .ZN(n38) );
  INV_X1 U213 ( .A(n170), .ZN(n94) );
  NOR2_X1 U214 ( .A1(n170), .A2(n39), .ZN(n34) );
  OAI21_X1 U215 ( .B1(n36), .B2(n40), .A(n37), .ZN(n35) );
  AOI21_X1 U216 ( .B1(n175), .B2(n30), .A(n23), .ZN(n21) );
  NAND2_X1 U217 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  NOR2_X1 U218 ( .A1(A[13]), .A2(B[13]), .ZN(n27) );
  INV_X1 U219 ( .A(n167), .ZN(n98) );
  NOR2_X1 U220 ( .A1(n167), .A2(n61), .ZN(n56) );
  OAI21_X1 U221 ( .B1(n58), .B2(n62), .A(n59), .ZN(n57) );
  NAND2_X1 U222 ( .A1(A[8]), .A2(B[8]), .ZN(n59) );
  XOR2_X1 U223 ( .A(n10), .B(n67), .Z(SUM[6]) );
  OAI21_X1 U224 ( .B1(n67), .B2(n65), .A(n66), .ZN(n64) );
  AOI21_X1 U225 ( .B1(n179), .B2(n72), .A(n69), .ZN(n67) );
  OAI21_X1 U226 ( .B1(n75), .B2(n73), .A(n74), .ZN(n72) );
  XOR2_X1 U227 ( .A(n12), .B(n75), .Z(SUM[4]) );
  OAI21_X1 U228 ( .B1(n55), .B2(n43), .A(n44), .ZN(n42) );
  NAND2_X1 U229 ( .A1(n165), .A2(n48), .ZN(n6) );
  NAND2_X1 U230 ( .A1(n165), .A2(n177), .ZN(n43) );
  XNOR2_X1 U231 ( .A(n19), .B(n1), .ZN(SUM[15]) );
  NAND2_X1 U232 ( .A1(A[14]), .A2(B[14]), .ZN(n25) );
  XNOR2_X1 U233 ( .A(n26), .B(n2), .ZN(SUM[14]) );
  XOR2_X1 U234 ( .A(n173), .B(n3), .Z(SUM[13]) );
  OAI21_X1 U235 ( .B1(n33), .B2(n164), .A(n28), .ZN(n26) );
  OAI21_X1 U236 ( .B1(n173), .B2(n20), .A(n21), .ZN(n19) );
  NAND2_X1 U237 ( .A1(A[10]), .A2(B[10]), .ZN(n48) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_4 ( clk, clear_acc, 
        data_out_x, data_out, data_out_w, data_out_b, wr_en_y, m_valid, 
        m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [3:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N27, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, n1, n2, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n87, n104, n113, n114, n115, n116, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n18), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n219), .CK(clk), .Q(n22) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n220), .CK(clk), .Q(n23) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n221), .CK(clk), .Q(n24) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n222), .CK(clk), .Q(n25) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n223), .CK(clk), .Q(n26) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n224), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n225), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n226), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n227), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n228), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n229), .CK(clk), .Q(n34) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n230), .CK(clk), .Q(n35) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n231), .CK(clk), .Q(n36) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n232), .CK(clk), .Q(n37) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n233), .CK(clk), .Q(n38) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n234), .CK(clk), .Q(n39) );
  DFF_X1 \f_reg[8]  ( .D(n79), .CK(clk), .Q(f[8]), .QN(n212) );
  DFF_X1 \f_reg[9]  ( .D(n78), .CK(clk), .Q(f[9]), .QN(n213) );
  DFF_X1 \f_reg[10]  ( .D(n77), .CK(clk), .Q(n49), .QN(n214) );
  DFF_X1 \f_reg[11]  ( .D(n76), .CK(clk), .Q(n47), .QN(n215) );
  DFF_X1 \f_reg[12]  ( .D(n4), .CK(clk), .Q(n46), .QN(n216) );
  DFF_X1 \f_reg[13]  ( .D(n75), .CK(clk), .Q(n44), .QN(n217) );
  DFF_X1 \f_reg[14]  ( .D(n5), .CK(clk), .Q(n43), .QN(n218) );
  DFF_X1 \f_reg[15]  ( .D(n9), .CK(clk), .Q(f[15]), .QN(n73) );
  DFF_X1 \data_out_reg[15]  ( .D(n113), .CK(clk), .Q(data_out[15]), .QN(n191)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n114), .CK(clk), .Q(data_out[14]), .QN(n190)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n115), .CK(clk), .Q(data_out[13]), .QN(n189)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n116), .CK(clk), .Q(data_out[12]), .QN(n188)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n164), .CK(clk), .Q(data_out[11]), .QN(n187)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n165), .CK(clk), .Q(data_out[10]), .QN(n186)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n166), .CK(clk), .Q(data_out[9]), .QN(n185) );
  DFF_X1 \data_out_reg[8]  ( .D(n167), .CK(clk), .Q(data_out[8]), .QN(n184) );
  DFF_X1 \data_out_reg[7]  ( .D(n168), .CK(clk), .Q(data_out[7]), .QN(n183) );
  DFF_X1 \data_out_reg[6]  ( .D(n169), .CK(clk), .Q(data_out[6]), .QN(n182) );
  DFF_X1 \data_out_reg[5]  ( .D(n170), .CK(clk), .Q(data_out[5]), .QN(n181) );
  DFF_X1 \data_out_reg[4]  ( .D(n171), .CK(clk), .Q(data_out[4]), .QN(n180) );
  DFF_X1 \data_out_reg[3]  ( .D(n172), .CK(clk), .Q(data_out[3]), .QN(n179) );
  DFF_X1 \data_out_reg[2]  ( .D(n173), .CK(clk), .Q(data_out[2]), .QN(n178) );
  DFF_X1 \data_out_reg[1]  ( .D(n174), .CK(clk), .Q(data_out[1]), .QN(n177) );
  DFF_X1 \data_out_reg[0]  ( .D(n175), .CK(clk), .Q(data_out[0]), .QN(n176) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_4_DW_mult_tc_1 mult_960 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_4_DW01_add_2 add_961 ( .A({n198, 
        n197, n196, n195, n194, n193, n207, n206, n205, n204, n203, n202, n201, 
        n200, n199, n192}), .B({f[15], n43, n44, n46, n47, n49, f[9:3], n57, 
        n59, n61}), .CI(1'b0), .SUM(adder) );
  DFF_X2 delay_reg ( .D(N27), .CK(clk), .Q(n2), .QN(n235) );
  DFF_X1 \f_reg[4]  ( .D(n83), .CK(clk), .Q(f[4]), .QN(n66) );
  DFF_X1 \f_reg[3]  ( .D(n84), .CK(clk), .Q(f[3]), .QN(n65) );
  DFF_X1 \f_reg[2]  ( .D(n85), .CK(clk), .Q(n57), .QN(n210) );
  DFF_X1 \f_reg[1]  ( .D(n87), .CK(clk), .Q(n59), .QN(n209) );
  DFF_X1 \f_reg[0]  ( .D(n104), .CK(clk), .Q(n61), .QN(n208) );
  DFF_X1 \f_reg[5]  ( .D(n82), .CK(clk), .Q(f[5]), .QN(n67) );
  DFF_X1 \f_reg[6]  ( .D(n81), .CK(clk), .Q(f[6]), .QN(n68) );
  DFF_X1 \f_reg[7]  ( .D(n80), .CK(clk), .Q(f[7]), .QN(n211) );
  MUX2_X2 U3 ( .A(N41), .B(n25), .S(n2), .Z(n195) );
  AND2_X1 U4 ( .A1(clear_acc_delay), .A2(n235), .ZN(n1) );
  AND2_X2 U5 ( .A1(n42), .A2(n19), .ZN(n16) );
  NAND3_X1 U6 ( .A1(n7), .A2(n6), .A3(n8), .ZN(n4) );
  NAND3_X1 U8 ( .A1(n14), .A2(n13), .A3(n15), .ZN(n5) );
  NAND2_X1 U9 ( .A1(data_out_b[12]), .A2(n18), .ZN(n6) );
  NAND2_X1 U10 ( .A1(adder[12]), .A2(n16), .ZN(n7) );
  NAND2_X1 U11 ( .A1(n63), .A2(n46), .ZN(n8) );
  NAND3_X1 U12 ( .A1(n11), .A2(n10), .A3(n12), .ZN(n9) );
  MUX2_X2 U13 ( .A(n26), .B(N40), .S(n235), .Z(n194) );
  MUX2_X2 U14 ( .A(n29), .B(N37), .S(n235), .Z(n206) );
  NAND2_X1 U15 ( .A1(data_out_b[15]), .A2(n18), .ZN(n10) );
  NAND2_X1 U16 ( .A1(adder[15]), .A2(n16), .ZN(n11) );
  NAND2_X1 U17 ( .A1(n63), .A2(f[15]), .ZN(n12) );
  NAND2_X1 U18 ( .A1(data_out_b[14]), .A2(n18), .ZN(n13) );
  NAND2_X1 U19 ( .A1(adder[14]), .A2(n16), .ZN(n14) );
  NAND2_X1 U20 ( .A1(n63), .A2(n43), .ZN(n15) );
  INV_X1 U21 ( .A(n19), .ZN(n18) );
  INV_X1 U22 ( .A(clear_acc), .ZN(n19) );
  NAND2_X1 U23 ( .A1(n17), .A2(N27), .ZN(n237) );
  OAI22_X1 U24 ( .A1(n179), .A2(n237), .B1(n65), .B2(n236), .ZN(n172) );
  OAI22_X1 U25 ( .A1(n180), .A2(n237), .B1(n66), .B2(n236), .ZN(n171) );
  OAI22_X1 U26 ( .A1(n181), .A2(n237), .B1(n67), .B2(n236), .ZN(n170) );
  OAI22_X1 U27 ( .A1(n182), .A2(n237), .B1(n68), .B2(n236), .ZN(n169) );
  OAI22_X1 U28 ( .A1(n183), .A2(n237), .B1(n211), .B2(n236), .ZN(n168) );
  OAI22_X1 U29 ( .A1(n184), .A2(n237), .B1(n212), .B2(n236), .ZN(n167) );
  OAI22_X1 U30 ( .A1(n185), .A2(n237), .B1(n213), .B2(n236), .ZN(n166) );
  MUX2_X1 U31 ( .A(n36), .B(N32), .S(n235), .Z(n201) );
  INV_X2 U32 ( .A(n42), .ZN(n63) );
  INV_X1 U33 ( .A(wr_en_y), .ZN(n17) );
  AND2_X1 U34 ( .A1(sel[0]), .A2(sel[1]), .ZN(n21) );
  INV_X1 U35 ( .A(m_ready), .ZN(n20) );
  NAND2_X1 U36 ( .A1(m_valid), .A2(n20), .ZN(n40) );
  OAI211_X1 U37 ( .C1(sel[2]), .C2(n21), .A(sel[3]), .B(n40), .ZN(N27) );
  MUX2_X1 U38 ( .A(n22), .B(N44), .S(n1), .Z(n219) );
  MUX2_X1 U39 ( .A(n22), .B(N44), .S(n235), .Z(n198) );
  MUX2_X1 U40 ( .A(n23), .B(N43), .S(n1), .Z(n220) );
  MUX2_X1 U41 ( .A(n23), .B(N43), .S(n235), .Z(n197) );
  MUX2_X1 U42 ( .A(n24), .B(N42), .S(n1), .Z(n221) );
  MUX2_X1 U43 ( .A(n24), .B(N42), .S(n235), .Z(n196) );
  MUX2_X1 U44 ( .A(n25), .B(N41), .S(n1), .Z(n222) );
  MUX2_X1 U45 ( .A(n26), .B(N40), .S(n1), .Z(n223) );
  MUX2_X1 U46 ( .A(n27), .B(N39), .S(n1), .Z(n224) );
  MUX2_X1 U47 ( .A(n27), .B(N39), .S(n235), .Z(n193) );
  MUX2_X1 U48 ( .A(n28), .B(N38), .S(n1), .Z(n225) );
  MUX2_X1 U49 ( .A(n28), .B(N38), .S(n235), .Z(n207) );
  MUX2_X1 U50 ( .A(n29), .B(N37), .S(n1), .Z(n226) );
  MUX2_X1 U51 ( .A(n32), .B(N36), .S(n1), .Z(n227) );
  MUX2_X1 U52 ( .A(n32), .B(N36), .S(n235), .Z(n205) );
  MUX2_X1 U53 ( .A(n33), .B(N35), .S(n1), .Z(n228) );
  MUX2_X1 U54 ( .A(n33), .B(N35), .S(n235), .Z(n204) );
  MUX2_X1 U55 ( .A(n34), .B(N34), .S(n1), .Z(n229) );
  MUX2_X1 U56 ( .A(n34), .B(N34), .S(n235), .Z(n203) );
  MUX2_X1 U57 ( .A(n35), .B(N33), .S(n1), .Z(n230) );
  MUX2_X1 U58 ( .A(n35), .B(N33), .S(n235), .Z(n202) );
  MUX2_X1 U59 ( .A(n36), .B(N32), .S(n1), .Z(n231) );
  MUX2_X1 U60 ( .A(n37), .B(N31), .S(n1), .Z(n232) );
  MUX2_X1 U61 ( .A(n37), .B(N31), .S(n235), .Z(n200) );
  MUX2_X1 U62 ( .A(n38), .B(N30), .S(n1), .Z(n233) );
  MUX2_X1 U63 ( .A(n38), .B(N30), .S(n235), .Z(n199) );
  MUX2_X1 U64 ( .A(n39), .B(N29), .S(n1), .Z(n234) );
  MUX2_X1 U65 ( .A(n39), .B(N29), .S(n235), .Z(n192) );
  INV_X1 U66 ( .A(n40), .ZN(n41) );
  OAI21_X1 U67 ( .B1(n41), .B2(n2), .A(n19), .ZN(n42) );
  AOI222_X1 U68 ( .A1(data_out_b[13]), .A2(n18), .B1(adder[13]), .B2(n16), 
        .C1(n63), .C2(n44), .ZN(n45) );
  INV_X1 U69 ( .A(n45), .ZN(n75) );
  AOI222_X1 U70 ( .A1(data_out_b[11]), .A2(n18), .B1(adder[11]), .B2(n16), 
        .C1(n63), .C2(n47), .ZN(n48) );
  INV_X1 U71 ( .A(n48), .ZN(n76) );
  AOI222_X1 U72 ( .A1(data_out_b[10]), .A2(n18), .B1(adder[10]), .B2(n16), 
        .C1(n63), .C2(n49), .ZN(n50) );
  INV_X1 U73 ( .A(n50), .ZN(n77) );
  AOI222_X1 U74 ( .A1(data_out_b[8]), .A2(n18), .B1(adder[8]), .B2(n16), .C1(
        n63), .C2(f[8]), .ZN(n51) );
  INV_X1 U75 ( .A(n51), .ZN(n79) );
  AOI222_X1 U76 ( .A1(data_out_b[7]), .A2(n18), .B1(adder[7]), .B2(n16), .C1(
        n63), .C2(f[7]), .ZN(n52) );
  INV_X1 U77 ( .A(n52), .ZN(n80) );
  AOI222_X1 U78 ( .A1(data_out_b[6]), .A2(n18), .B1(adder[6]), .B2(n16), .C1(
        n63), .C2(f[6]), .ZN(n53) );
  INV_X1 U79 ( .A(n53), .ZN(n81) );
  AOI222_X1 U80 ( .A1(data_out_b[5]), .A2(n18), .B1(adder[5]), .B2(n16), .C1(
        n63), .C2(f[5]), .ZN(n54) );
  INV_X1 U81 ( .A(n54), .ZN(n82) );
  AOI222_X1 U82 ( .A1(data_out_b[4]), .A2(n18), .B1(adder[4]), .B2(n16), .C1(
        n63), .C2(f[4]), .ZN(n55) );
  INV_X1 U83 ( .A(n55), .ZN(n83) );
  AOI222_X1 U84 ( .A1(data_out_b[3]), .A2(n18), .B1(adder[3]), .B2(n16), .C1(
        n63), .C2(f[3]), .ZN(n56) );
  INV_X1 U85 ( .A(n56), .ZN(n84) );
  AOI222_X1 U86 ( .A1(data_out_b[2]), .A2(n18), .B1(adder[2]), .B2(n16), .C1(
        n63), .C2(n57), .ZN(n58) );
  INV_X1 U87 ( .A(n58), .ZN(n85) );
  AOI222_X1 U88 ( .A1(data_out_b[1]), .A2(n18), .B1(adder[1]), .B2(n16), .C1(
        n63), .C2(n59), .ZN(n60) );
  INV_X1 U89 ( .A(n60), .ZN(n87) );
  AOI222_X1 U90 ( .A1(data_out_b[0]), .A2(n18), .B1(adder[0]), .B2(n16), .C1(
        n63), .C2(n61), .ZN(n62) );
  INV_X1 U91 ( .A(n62), .ZN(n104) );
  AOI222_X1 U92 ( .A1(data_out_b[9]), .A2(n18), .B1(adder[9]), .B2(n16), .C1(
        n63), .C2(f[9]), .ZN(n64) );
  INV_X1 U93 ( .A(n64), .ZN(n78) );
  NOR4_X1 U94 ( .A1(n47), .A2(n46), .A3(n44), .A4(n43), .ZN(n72) );
  NOR4_X1 U95 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n49), .ZN(n71) );
  NAND4_X1 U96 ( .A1(n68), .A2(n67), .A3(n66), .A4(n65), .ZN(n69) );
  NOR4_X1 U97 ( .A1(n69), .A2(n61), .A3(n59), .A4(n57), .ZN(n70) );
  NAND3_X1 U98 ( .A1(n72), .A2(n71), .A3(n70), .ZN(n74) );
  NAND3_X1 U99 ( .A1(wr_en_y), .A2(n74), .A3(n73), .ZN(n236) );
  OAI22_X1 U100 ( .A1(n176), .A2(n237), .B1(n208), .B2(n236), .ZN(n175) );
  OAI22_X1 U101 ( .A1(n177), .A2(n237), .B1(n209), .B2(n236), .ZN(n174) );
  OAI22_X1 U102 ( .A1(n178), .A2(n237), .B1(n210), .B2(n236), .ZN(n173) );
  OAI22_X1 U103 ( .A1(n186), .A2(n237), .B1(n214), .B2(n236), .ZN(n165) );
  OAI22_X1 U104 ( .A1(n187), .A2(n237), .B1(n215), .B2(n236), .ZN(n164) );
  OAI22_X1 U105 ( .A1(n188), .A2(n237), .B1(n216), .B2(n236), .ZN(n116) );
  OAI22_X1 U106 ( .A1(n189), .A2(n237), .B1(n217), .B2(n236), .ZN(n115) );
  OAI22_X1 U107 ( .A1(n190), .A2(n237), .B1(n218), .B2(n236), .ZN(n114) );
  OAI22_X1 U108 ( .A1(n191), .A2(n237), .B1(n73), .B2(n236), .ZN(n113) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_3_DW_mult_tc_1 ( a, b, 
        product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n9, n12, n13, n16, n18, n19, n21, n23, n25, n27, n29, n31,
         n32, n34, n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n50,
         n52, n53, n55, n56, n57, n58, n59, n62, n63, n64, n65, n67, n69, n70,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n93, n95, n96, n97, n98, n99, n101, n103,
         n104, n105, n106, n107, n109, n111, n112, n113, n114, n115, n117,
         n119, n120, n122, n125, n127, n135, n139, n141, n142, n143, n144,
         n145, n147, n148, n149, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n239, n241, n243, n247, n249, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n418, n419, n420, n421, n422, n423, n424, n426, n427, n428, n429,
         n430, n432, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U148 ( .A(n265), .B(n144), .Z(n145) );
  XOR2_X1 U152 ( .A(n301), .B(n148), .Z(n149) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U161 ( .A(n177), .B(n168), .CI(n166), .CO(n163), .S(n164) );
  FA_X1 U162 ( .A(n170), .B(n172), .CI(n179), .CO(n165), .S(n166) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n291), .CI(n263), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n252), .B(n317), .CO(n173), .S(n174) );
  FA_X1 U167 ( .A(n180), .B(n187), .CI(n178), .CO(n175), .S(n176) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U169 ( .A(n193), .B(n282), .CI(n191), .CO(n179), .S(n180) );
  FA_X1 U170 ( .A(n268), .B(n274), .CI(n292), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U172 ( .A(n197), .B(n190), .CI(n188), .CO(n185), .S(n186) );
  FA_X1 U173 ( .A(n199), .B(n201), .CI(n192), .CO(n187), .S(n188) );
  FA_X1 U174 ( .A(n275), .B(n293), .CI(n194), .CO(n189), .S(n190) );
  FA_X1 U175 ( .A(n283), .B(n253), .CI(n305), .CO(n191), .S(n192) );
  HA_X1 U176 ( .A(n319), .B(n269), .CO(n193), .S(n194) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U179 ( .A(n276), .B(n284), .CI(n294), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n320), .B(n270), .CI(n306), .CO(n201), .S(n202) );
  FA_X1 U181 ( .A(n208), .B(n213), .CI(n206), .CO(n203), .S(n204) );
  FA_X1 U182 ( .A(n215), .B(n307), .CI(n210), .CO(n205), .S(n206) );
  FA_X1 U183 ( .A(n254), .B(n285), .CI(n295), .CO(n207), .S(n208) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U187 ( .A(n322), .B(n278), .CI(n308), .CO(n215), .S(n216) );
  FA_X1 U189 ( .A(n255), .B(n309), .CI(n297), .CO(n219), .S(n220) );
  FA_X1 U192 ( .A(n324), .B(n288), .CI(n310), .CO(n225), .S(n226) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  HA_X1 U194 ( .A(n311), .B(n325), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n326), .B(n300), .CI(n312), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  BUF_X1 U414 ( .A(n45), .Z(n490) );
  BUF_X2 U415 ( .A(n584), .Z(n528) );
  BUF_X1 U416 ( .A(n76), .Z(n491) );
  INV_X1 U417 ( .A(n523), .ZN(n37) );
  OR2_X2 U418 ( .A1(n539), .A2(n564), .ZN(n18) );
  AOI21_X1 U419 ( .B1(n568), .B2(n120), .A(n117), .ZN(n115) );
  OR2_X1 U420 ( .A1(n329), .A2(n258), .ZN(n492) );
  XNOR2_X1 U421 ( .A(n536), .B(n493), .ZN(product[7]) );
  AND2_X1 U422 ( .A1(n521), .A2(n98), .ZN(n493) );
  BUF_X1 U423 ( .A(n104), .Z(n535) );
  BUF_X2 U424 ( .A(n584), .Z(n529) );
  INV_X1 U425 ( .A(n241), .ZN(n494) );
  INV_X1 U426 ( .A(n241), .ZN(n548) );
  XNOR2_X1 U427 ( .A(n45), .B(n495), .ZN(product[12]) );
  AND2_X1 U428 ( .A1(n542), .A2(n79), .ZN(n495) );
  CLKBUF_X1 U429 ( .A(n39), .Z(n496) );
  AOI21_X1 U430 ( .B1(n96), .B2(n567), .A(n93), .ZN(n497) );
  XOR2_X1 U431 ( .A(n594), .B(a[10]), .Z(n498) );
  NAND2_X1 U432 ( .A1(n432), .A2(n578), .ZN(n499) );
  INV_X1 U433 ( .A(n587), .ZN(n500) );
  INV_X1 U434 ( .A(n590), .ZN(n501) );
  OAI21_X1 U435 ( .B1(n99), .B2(n97), .A(n98), .ZN(n502) );
  CLKBUF_X1 U436 ( .A(n591), .Z(n503) );
  CLKBUF_X3 U437 ( .A(n9), .Z(n579) );
  CLKBUF_X1 U438 ( .A(n222), .Z(n504) );
  AOI21_X1 U439 ( .B1(n502), .B2(n567), .A(n93), .ZN(n505) );
  INV_X2 U440 ( .A(n588), .ZN(n587) );
  XOR2_X1 U441 ( .A(n296), .B(n286), .Z(n506) );
  XOR2_X1 U442 ( .A(n506), .B(n221), .Z(n214) );
  XOR2_X1 U443 ( .A(n216), .B(n219), .Z(n507) );
  XOR2_X1 U444 ( .A(n507), .B(n214), .Z(n212) );
  NAND2_X1 U445 ( .A1(n296), .A2(n286), .ZN(n508) );
  NAND2_X1 U446 ( .A1(n296), .A2(n221), .ZN(n509) );
  NAND2_X1 U447 ( .A1(n286), .A2(n221), .ZN(n510) );
  NAND3_X1 U448 ( .A1(n508), .A2(n509), .A3(n510), .ZN(n213) );
  NAND2_X1 U449 ( .A1(n216), .A2(n219), .ZN(n511) );
  NAND2_X1 U450 ( .A1(n216), .A2(n214), .ZN(n512) );
  NAND2_X1 U451 ( .A1(n219), .A2(n214), .ZN(n513) );
  NAND3_X1 U452 ( .A1(n511), .A2(n512), .A3(n513), .ZN(n211) );
  BUF_X1 U453 ( .A(n591), .Z(n534) );
  XNOR2_X1 U454 ( .A(n226), .B(n514), .ZN(n224) );
  XNOR2_X1 U455 ( .A(n229), .B(n298), .ZN(n514) );
  XOR2_X1 U456 ( .A(n225), .B(n222), .Z(n515) );
  XOR2_X1 U457 ( .A(n220), .B(n515), .Z(n218) );
  NAND2_X1 U458 ( .A1(n220), .A2(n225), .ZN(n516) );
  NAND2_X1 U459 ( .A1(n220), .A2(n504), .ZN(n517) );
  NAND2_X1 U460 ( .A1(n225), .A2(n504), .ZN(n518) );
  NAND3_X1 U461 ( .A1(n516), .A2(n517), .A3(n518), .ZN(n217) );
  OR2_X1 U462 ( .A1(n228), .A2(n231), .ZN(n519) );
  XNOR2_X1 U463 ( .A(n88), .B(n520), .ZN(product[10]) );
  NAND2_X1 U464 ( .A1(n538), .A2(n86), .ZN(n520) );
  CLKBUF_X3 U465 ( .A(n21), .Z(n577) );
  OR2_X1 U466 ( .A1(n218), .A2(n223), .ZN(n521) );
  XOR2_X1 U467 ( .A(n287), .B(n323), .Z(n222) );
  BUF_X1 U468 ( .A(n21), .Z(n576) );
  XNOR2_X1 U469 ( .A(n198), .B(n522), .ZN(n196) );
  XNOR2_X1 U470 ( .A(n205), .B(n200), .ZN(n522) );
  AND2_X1 U471 ( .A1(n323), .A2(n287), .ZN(n221) );
  XNOR2_X1 U472 ( .A(n596), .B(a[12]), .ZN(n523) );
  OR2_X2 U473 ( .A1(n556), .A2(n565), .ZN(n524) );
  OR2_X2 U474 ( .A1(n556), .A2(n565), .ZN(n525) );
  OR2_X1 U475 ( .A1(n556), .A2(n565), .ZN(n6) );
  OR2_X1 U476 ( .A1(n551), .A2(n78), .ZN(n526) );
  INV_X1 U477 ( .A(n583), .ZN(n527) );
  INV_X1 U478 ( .A(n239), .ZN(n530) );
  XOR2_X1 U479 ( .A(n594), .B(a[10]), .Z(n32) );
  INV_X1 U480 ( .A(n591), .ZN(n531) );
  NAND2_X1 U481 ( .A1(n432), .A2(n578), .ZN(n532) );
  BUF_X2 U482 ( .A(n9), .Z(n578) );
  INV_X1 U483 ( .A(n501), .ZN(n533) );
  NAND2_X1 U484 ( .A1(n429), .A2(n27), .ZN(n29) );
  XNOR2_X1 U485 ( .A(n594), .B(a[8]), .ZN(n429) );
  AOI21_X1 U486 ( .B1(n569), .B2(n535), .A(n101), .ZN(n536) );
  XNOR2_X1 U487 ( .A(n597), .B(a[14]), .ZN(n537) );
  INV_X2 U488 ( .A(n598), .ZN(n597) );
  XNOR2_X1 U489 ( .A(n596), .B(a[10]), .ZN(n428) );
  OAI21_X1 U490 ( .B1(n113), .B2(n115), .A(n114), .ZN(n112) );
  OR2_X1 U491 ( .A1(n196), .A2(n203), .ZN(n538) );
  XNOR2_X1 U492 ( .A(n501), .B(a[4]), .ZN(n539) );
  AOI21_X1 U493 ( .B1(n555), .B2(n80), .A(n81), .ZN(n540) );
  AOI21_X1 U494 ( .B1(n555), .B2(n80), .A(n81), .ZN(n45) );
  BUF_X2 U495 ( .A(n582), .Z(n541) );
  OR2_X1 U496 ( .A1(n176), .A2(n185), .ZN(n542) );
  NAND2_X1 U497 ( .A1(n428), .A2(n498), .ZN(n543) );
  NAND2_X1 U498 ( .A1(n428), .A2(n32), .ZN(n34) );
  INV_X1 U499 ( .A(n564), .ZN(n16) );
  NAND2_X1 U500 ( .A1(n430), .A2(n576), .ZN(n544) );
  NAND2_X1 U501 ( .A1(n430), .A2(n576), .ZN(n545) );
  NAND2_X1 U502 ( .A1(n430), .A2(n576), .ZN(n23) );
  CLKBUF_X1 U503 ( .A(n584), .Z(n546) );
  CLKBUF_X3 U504 ( .A(n584), .Z(n547) );
  INV_X1 U505 ( .A(n585), .ZN(n584) );
  XOR2_X1 U506 ( .A(n592), .B(a[8]), .Z(n27) );
  XNOR2_X1 U507 ( .A(n271), .B(n549), .ZN(n147) );
  XNOR2_X1 U508 ( .A(n289), .B(n279), .ZN(n549) );
  CLKBUF_X1 U509 ( .A(n107), .Z(n550) );
  NOR2_X1 U510 ( .A1(n164), .A2(n175), .ZN(n551) );
  NOR2_X1 U511 ( .A1(n164), .A2(n175), .ZN(n75) );
  INV_X1 U512 ( .A(n13), .ZN(n590) );
  XOR2_X1 U513 ( .A(a[2]), .B(n585), .Z(n9) );
  NAND2_X1 U514 ( .A1(n198), .A2(n205), .ZN(n552) );
  NAND2_X1 U515 ( .A1(n198), .A2(n200), .ZN(n553) );
  NAND2_X1 U516 ( .A1(n205), .A2(n200), .ZN(n554) );
  NAND3_X1 U517 ( .A1(n552), .A2(n553), .A3(n554), .ZN(n195) );
  NOR2_X1 U518 ( .A1(n196), .A2(n203), .ZN(n85) );
  XNOR2_X1 U519 ( .A(a[6]), .B(n592), .ZN(n430) );
  OAI21_X1 U520 ( .B1(n497), .B2(n89), .A(n90), .ZN(n555) );
  INV_X2 U521 ( .A(n596), .ZN(n595) );
  XNOR2_X1 U522 ( .A(n588), .B(a[2]), .ZN(n432) );
  INV_X1 U523 ( .A(n588), .ZN(n586) );
  XNOR2_X1 U524 ( .A(n583), .B(n249), .ZN(n556) );
  NAND2_X1 U525 ( .A1(n226), .A2(n229), .ZN(n557) );
  NAND2_X1 U526 ( .A1(n226), .A2(n298), .ZN(n558) );
  NAND2_X1 U527 ( .A1(n229), .A2(n298), .ZN(n559) );
  NAND3_X1 U528 ( .A1(n557), .A2(n558), .A3(n559), .ZN(n223) );
  OR2_X1 U529 ( .A1(n204), .A2(n211), .ZN(n560) );
  NAND2_X1 U530 ( .A1(n578), .A2(n432), .ZN(n561) );
  NAND2_X1 U531 ( .A1(n578), .A2(n432), .ZN(n562) );
  NAND2_X1 U532 ( .A1(n432), .A2(n578), .ZN(n12) );
  NOR2_X1 U533 ( .A1(n186), .A2(n195), .ZN(n563) );
  NOR2_X1 U534 ( .A1(n186), .A2(n195), .ZN(n82) );
  XOR2_X1 U535 ( .A(n590), .B(a[6]), .Z(n21) );
  XNOR2_X1 U536 ( .A(n588), .B(a[4]), .ZN(n564) );
  INV_X1 U537 ( .A(n582), .ZN(n565) );
  INV_X2 U538 ( .A(n594), .ZN(n593) );
  INV_X2 U539 ( .A(n592), .ZN(n591) );
  BUF_X1 U540 ( .A(n43), .Z(n580) );
  NAND2_X1 U541 ( .A1(n566), .A2(n69), .ZN(n47) );
  INV_X1 U542 ( .A(n74), .ZN(n72) );
  INV_X1 U543 ( .A(n69), .ZN(n67) );
  NAND2_X1 U544 ( .A1(n73), .A2(n566), .ZN(n64) );
  INV_X1 U545 ( .A(n95), .ZN(n93) );
  OAI21_X1 U546 ( .B1(n505), .B2(n89), .A(n90), .ZN(n88) );
  NAND2_X1 U547 ( .A1(n90), .A2(n560), .ZN(n52) );
  OR2_X1 U548 ( .A1(n152), .A2(n163), .ZN(n566) );
  NOR2_X1 U549 ( .A1(n563), .A2(n85), .ZN(n80) );
  OAI21_X1 U550 ( .B1(n82), .B2(n86), .A(n83), .ZN(n81) );
  NAND2_X1 U551 ( .A1(n567), .A2(n95), .ZN(n53) );
  OAI21_X1 U552 ( .B1(n75), .B2(n79), .A(n76), .ZN(n74) );
  NAND2_X1 U553 ( .A1(n125), .A2(n491), .ZN(n48) );
  INV_X1 U554 ( .A(n551), .ZN(n125) );
  NOR2_X1 U555 ( .A1(n551), .A2(n78), .ZN(n73) );
  NAND2_X1 U556 ( .A1(n152), .A2(n163), .ZN(n69) );
  NAND2_X1 U557 ( .A1(n127), .A2(n83), .ZN(n50) );
  OAI21_X1 U558 ( .B1(n87), .B2(n85), .A(n86), .ZN(n84) );
  INV_X1 U559 ( .A(n563), .ZN(n127) );
  NAND2_X1 U560 ( .A1(n135), .A2(n114), .ZN(n58) );
  INV_X1 U561 ( .A(n113), .ZN(n135) );
  NAND2_X1 U562 ( .A1(n106), .A2(n519), .ZN(n56) );
  AOI21_X1 U563 ( .B1(n104), .B2(n569), .A(n101), .ZN(n99) );
  INV_X1 U564 ( .A(n103), .ZN(n101) );
  AOI21_X1 U565 ( .B1(n570), .B2(n112), .A(n109), .ZN(n107) );
  INV_X1 U566 ( .A(n111), .ZN(n109) );
  NOR2_X1 U567 ( .A1(n176), .A2(n185), .ZN(n78) );
  OR2_X1 U568 ( .A1(n212), .A2(n217), .ZN(n567) );
  INV_X1 U569 ( .A(n119), .ZN(n117) );
  INV_X1 U570 ( .A(n122), .ZN(n120) );
  XNOR2_X1 U571 ( .A(n57), .B(n112), .ZN(product[4]) );
  NAND2_X1 U572 ( .A1(n570), .A2(n111), .ZN(n57) );
  XNOR2_X1 U573 ( .A(n59), .B(n120), .ZN(product[2]) );
  NAND2_X1 U574 ( .A1(n568), .A2(n119), .ZN(n59) );
  NAND2_X1 U575 ( .A1(n176), .A2(n185), .ZN(n79) );
  NAND2_X1 U576 ( .A1(n196), .A2(n203), .ZN(n86) );
  NAND2_X1 U577 ( .A1(n164), .A2(n175), .ZN(n76) );
  NAND2_X1 U578 ( .A1(n186), .A2(n195), .ZN(n83) );
  NAND2_X1 U579 ( .A1(n212), .A2(n217), .ZN(n95) );
  XNOR2_X1 U580 ( .A(n63), .B(n46), .ZN(product[15]) );
  NAND2_X1 U581 ( .A1(n571), .A2(n62), .ZN(n46) );
  AOI21_X1 U582 ( .B1(n566), .B2(n74), .A(n67), .ZN(n65) );
  XNOR2_X1 U583 ( .A(n55), .B(n535), .ZN(product[6]) );
  NAND2_X1 U584 ( .A1(n569), .A2(n103), .ZN(n55) );
  NOR2_X1 U585 ( .A1(n234), .A2(n257), .ZN(n113) );
  OR2_X1 U586 ( .A1(n328), .A2(n314), .ZN(n568) );
  NOR2_X1 U587 ( .A1(n228), .A2(n231), .ZN(n105) );
  NOR2_X1 U588 ( .A1(n218), .A2(n223), .ZN(n97) );
  NAND2_X1 U589 ( .A1(n224), .A2(n227), .ZN(n103) );
  OR2_X1 U590 ( .A1(n224), .A2(n227), .ZN(n569) );
  OR2_X1 U591 ( .A1(n232), .A2(n233), .ZN(n570) );
  NAND2_X1 U592 ( .A1(n218), .A2(n223), .ZN(n98) );
  NAND2_X1 U593 ( .A1(n228), .A2(n231), .ZN(n106) );
  NAND2_X1 U594 ( .A1(n232), .A2(n233), .ZN(n111) );
  INV_X1 U595 ( .A(n537), .ZN(n235) );
  OR2_X1 U596 ( .A1(n151), .A2(n139), .ZN(n571) );
  AND2_X1 U597 ( .A1(n492), .A2(n122), .ZN(product[1]) );
  XNOR2_X1 U598 ( .A(n597), .B(a[14]), .ZN(n41) );
  INV_X1 U599 ( .A(n249), .ZN(n582) );
  OR2_X1 U600 ( .A1(n580), .A2(n500), .ZN(n392) );
  OAI22_X1 U601 ( .A1(n39), .A2(n336), .B1(n37), .B2(n335), .ZN(n263) );
  XNOR2_X1 U602 ( .A(n589), .B(n580), .ZN(n376) );
  AND2_X1 U603 ( .A1(n581), .A2(n564), .ZN(n300) );
  XNOR2_X1 U604 ( .A(n593), .B(n580), .ZN(n352) );
  XNOR2_X1 U605 ( .A(n155), .B(n573), .ZN(n139) );
  XNOR2_X1 U606 ( .A(n153), .B(n141), .ZN(n573) );
  XNOR2_X1 U607 ( .A(n157), .B(n574), .ZN(n141) );
  XNOR2_X1 U608 ( .A(n145), .B(n143), .ZN(n574) );
  OAI22_X1 U609 ( .A1(n39), .A2(n598), .B1(n337), .B2(n37), .ZN(n252) );
  OR2_X1 U610 ( .A1(n580), .A2(n598), .ZN(n337) );
  OAI22_X1 U611 ( .A1(n42), .A2(n599), .B1(n332), .B2(n537), .ZN(n251) );
  OR2_X1 U612 ( .A1(n580), .A2(n599), .ZN(n332) );
  XNOR2_X1 U613 ( .A(n595), .B(n580), .ZN(n343) );
  XNOR2_X1 U614 ( .A(n159), .B(n575), .ZN(n142) );
  XNOR2_X1 U615 ( .A(n315), .B(n261), .ZN(n575) );
  XNOR2_X1 U616 ( .A(n597), .B(n580), .ZN(n336) );
  NAND2_X1 U617 ( .A1(n427), .A2(n37), .ZN(n39) );
  XOR2_X1 U618 ( .A(n597), .B(a[12]), .Z(n427) );
  AND2_X1 U619 ( .A1(n581), .A2(n241), .ZN(n278) );
  AND2_X1 U620 ( .A1(n581), .A2(n235), .ZN(n260) );
  OAI22_X1 U621 ( .A1(n496), .A2(n335), .B1(n37), .B2(n334), .ZN(n262) );
  AND2_X1 U622 ( .A1(n581), .A2(n243), .ZN(n288) );
  AND2_X1 U623 ( .A1(n581), .A2(n239), .ZN(n270) );
  INV_X1 U624 ( .A(n25), .ZN(n594) );
  NAND2_X1 U625 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U626 ( .A(n40), .B(a[14]), .Z(n426) );
  INV_X1 U627 ( .A(n7), .ZN(n588) );
  XNOR2_X1 U628 ( .A(n503), .B(n580), .ZN(n363) );
  AND2_X1 U629 ( .A1(n581), .A2(n247), .ZN(n314) );
  AND2_X1 U630 ( .A1(n581), .A2(n523), .ZN(n264) );
  AND2_X1 U631 ( .A1(n581), .A2(n249), .ZN(product[0]) );
  OR2_X1 U632 ( .A1(n580), .A2(n596), .ZN(n344) );
  OR2_X1 U633 ( .A1(n580), .A2(n594), .ZN(n353) );
  OR2_X1 U634 ( .A1(n580), .A2(n531), .ZN(n364) );
  OR2_X1 U635 ( .A1(n580), .A2(n533), .ZN(n377) );
  XNOR2_X1 U636 ( .A(n503), .B(b[9]), .ZN(n354) );
  OAI22_X1 U637 ( .A1(n496), .A2(n334), .B1(n37), .B2(n333), .ZN(n261) );
  XNOR2_X1 U638 ( .A(n597), .B(n422), .ZN(n333) );
  XNOR2_X1 U639 ( .A(n589), .B(b[11]), .ZN(n365) );
  XNOR2_X1 U640 ( .A(n597), .B(n424), .ZN(n335) );
  XNOR2_X1 U641 ( .A(n597), .B(n423), .ZN(n334) );
  OAI22_X1 U642 ( .A1(n42), .A2(n331), .B1(n330), .B2(n537), .ZN(n259) );
  XNOR2_X1 U643 ( .A(n40), .B(n424), .ZN(n330) );
  XNOR2_X1 U644 ( .A(n40), .B(n580), .ZN(n331) );
  XNOR2_X1 U645 ( .A(n593), .B(n418), .ZN(n345) );
  XNOR2_X1 U646 ( .A(n595), .B(n420), .ZN(n338) );
  XNOR2_X1 U647 ( .A(n587), .B(b[13]), .ZN(n378) );
  XNOR2_X1 U648 ( .A(n595), .B(n424), .ZN(n342) );
  XNOR2_X1 U649 ( .A(n593), .B(n424), .ZN(n351) );
  XNOR2_X1 U650 ( .A(n591), .B(n424), .ZN(n362) );
  XNOR2_X1 U651 ( .A(n595), .B(n423), .ZN(n341) );
  XNOR2_X1 U652 ( .A(n595), .B(n422), .ZN(n340) );
  XNOR2_X1 U653 ( .A(n595), .B(n421), .ZN(n339) );
  XNOR2_X1 U654 ( .A(n587), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U655 ( .A(n587), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U656 ( .A(n587), .B(n418), .ZN(n384) );
  XNOR2_X1 U657 ( .A(n587), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U658 ( .A(n587), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U659 ( .A(n587), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U660 ( .A(n587), .B(n419), .ZN(n385) );
  XNOR2_X1 U661 ( .A(n547), .B(b[11]), .ZN(n397) );
  XNOR2_X1 U662 ( .A(n528), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U663 ( .A(n546), .B(b[13]), .ZN(n395) );
  XNOR2_X1 U664 ( .A(n547), .B(b[14]), .ZN(n394) );
  XNOR2_X1 U665 ( .A(n589), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U666 ( .A(n589), .B(n418), .ZN(n369) );
  XNOR2_X1 U667 ( .A(n589), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U668 ( .A(n589), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U669 ( .A(n593), .B(n423), .ZN(n350) );
  XNOR2_X1 U670 ( .A(n534), .B(n423), .ZN(n361) );
  XNOR2_X1 U671 ( .A(n591), .B(n422), .ZN(n360) );
  XNOR2_X1 U672 ( .A(n593), .B(n422), .ZN(n349) );
  XNOR2_X1 U673 ( .A(n591), .B(n421), .ZN(n359) );
  XNOR2_X1 U674 ( .A(n591), .B(n420), .ZN(n358) );
  XNOR2_X1 U675 ( .A(n593), .B(n421), .ZN(n348) );
  XNOR2_X1 U676 ( .A(n593), .B(n420), .ZN(n347) );
  XNOR2_X1 U677 ( .A(n591), .B(n418), .ZN(n356) );
  XNOR2_X1 U678 ( .A(n534), .B(n419), .ZN(n357) );
  XNOR2_X1 U679 ( .A(n593), .B(n419), .ZN(n346) );
  XNOR2_X1 U680 ( .A(n591), .B(b[8]), .ZN(n355) );
  XNOR2_X1 U681 ( .A(n546), .B(b[15]), .ZN(n393) );
  BUF_X1 U682 ( .A(n43), .Z(n581) );
  NAND2_X1 U683 ( .A1(n328), .A2(n314), .ZN(n119) );
  XNOR2_X1 U684 ( .A(n84), .B(n50), .ZN(product[11]) );
  INV_X1 U685 ( .A(n19), .ZN(n592) );
  XNOR2_X1 U686 ( .A(n70), .B(n47), .ZN(product[14]) );
  OAI22_X1 U687 ( .A1(n543), .A2(n339), .B1(n338), .B2(n530), .ZN(n265) );
  OAI22_X1 U688 ( .A1(n543), .A2(n340), .B1(n339), .B2(n530), .ZN(n266) );
  OAI22_X1 U689 ( .A1(n543), .A2(n341), .B1(n340), .B2(n530), .ZN(n267) );
  OAI22_X1 U690 ( .A1(n543), .A2(n342), .B1(n341), .B2(n530), .ZN(n268) );
  OAI22_X1 U691 ( .A1(n34), .A2(n343), .B1(n342), .B2(n498), .ZN(n269) );
  INV_X1 U692 ( .A(n32), .ZN(n239) );
  OAI22_X1 U693 ( .A1(n34), .A2(n596), .B1(n344), .B2(n498), .ZN(n253) );
  NAND2_X1 U694 ( .A1(n204), .A2(n211), .ZN(n90) );
  NOR2_X1 U695 ( .A1(n204), .A2(n211), .ZN(n89) );
  OAI22_X1 U696 ( .A1(n29), .A2(n346), .B1(n345), .B2(n494), .ZN(n271) );
  OAI22_X1 U697 ( .A1(n29), .A2(n350), .B1(n349), .B2(n494), .ZN(n275) );
  OAI22_X1 U698 ( .A1(n29), .A2(n347), .B1(n346), .B2(n494), .ZN(n272) );
  OAI22_X1 U699 ( .A1(n29), .A2(n348), .B1(n347), .B2(n548), .ZN(n273) );
  OAI22_X1 U700 ( .A1(n29), .A2(n349), .B1(n348), .B2(n548), .ZN(n274) );
  INV_X1 U701 ( .A(n27), .ZN(n241) );
  OAI22_X1 U702 ( .A1(n29), .A2(n594), .B1(n353), .B2(n494), .ZN(n254) );
  OAI22_X1 U703 ( .A1(n29), .A2(n351), .B1(n350), .B2(n548), .ZN(n276) );
  OAI22_X1 U704 ( .A1(n29), .A2(n352), .B1(n351), .B2(n548), .ZN(n277) );
  INV_X1 U705 ( .A(n88), .ZN(n87) );
  NAND2_X1 U706 ( .A1(n151), .A2(n139), .ZN(n62) );
  INV_X1 U707 ( .A(n585), .ZN(n583) );
  INV_X1 U708 ( .A(n1), .ZN(n585) );
  OR2_X1 U709 ( .A1(n580), .A2(n527), .ZN(n409) );
  XNOR2_X1 U710 ( .A(n77), .B(n48), .ZN(product[13]) );
  OAI22_X1 U711 ( .A1(n544), .A2(n358), .B1(n357), .B2(n577), .ZN(n282) );
  OAI22_X1 U712 ( .A1(n545), .A2(n356), .B1(n355), .B2(n577), .ZN(n280) );
  OAI22_X1 U713 ( .A1(n544), .A2(n362), .B1(n361), .B2(n577), .ZN(n286) );
  OAI22_X1 U714 ( .A1(n544), .A2(n357), .B1(n356), .B2(n577), .ZN(n281) );
  OAI22_X1 U715 ( .A1(n544), .A2(n360), .B1(n359), .B2(n577), .ZN(n284) );
  OAI22_X1 U716 ( .A1(n545), .A2(n361), .B1(n360), .B2(n577), .ZN(n285) );
  OAI22_X1 U717 ( .A1(n545), .A2(n531), .B1(n364), .B2(n577), .ZN(n255) );
  OAI22_X1 U718 ( .A1(n544), .A2(n363), .B1(n362), .B2(n577), .ZN(n287) );
  OAI22_X1 U719 ( .A1(n545), .A2(n355), .B1(n354), .B2(n577), .ZN(n279) );
  XNOR2_X1 U720 ( .A(n589), .B(n421), .ZN(n372) );
  OAI22_X1 U721 ( .A1(n359), .A2(n23), .B1(n358), .B2(n577), .ZN(n283) );
  XNOR2_X1 U722 ( .A(n589), .B(n423), .ZN(n374) );
  XNOR2_X1 U723 ( .A(n589), .B(n424), .ZN(n375) );
  XNOR2_X1 U724 ( .A(n501), .B(n422), .ZN(n373) );
  XNOR2_X1 U725 ( .A(n501), .B(n419), .ZN(n370) );
  XNOR2_X1 U726 ( .A(n501), .B(n420), .ZN(n371) );
  INV_X1 U727 ( .A(n577), .ZN(n243) );
  OAI21_X1 U728 ( .B1(n99), .B2(n97), .A(n98), .ZN(n96) );
  OAI22_X1 U729 ( .A1(n18), .A2(n370), .B1(n369), .B2(n16), .ZN(n293) );
  OAI22_X1 U730 ( .A1(n18), .A2(n367), .B1(n366), .B2(n16), .ZN(n290) );
  OAI22_X1 U731 ( .A1(n18), .A2(n368), .B1(n367), .B2(n16), .ZN(n291) );
  OAI22_X1 U732 ( .A1(n18), .A2(n375), .B1(n374), .B2(n16), .ZN(n298) );
  OAI22_X1 U733 ( .A1(n18), .A2(n371), .B1(n370), .B2(n16), .ZN(n294) );
  OAI22_X1 U734 ( .A1(n18), .A2(n373), .B1(n372), .B2(n16), .ZN(n296) );
  OAI22_X1 U735 ( .A1(n18), .A2(n369), .B1(n368), .B2(n16), .ZN(n292) );
  OAI22_X1 U736 ( .A1(n18), .A2(n533), .B1(n377), .B2(n16), .ZN(n256) );
  OAI22_X1 U737 ( .A1(n18), .A2(n372), .B1(n371), .B2(n16), .ZN(n295) );
  OAI22_X1 U738 ( .A1(n18), .A2(n376), .B1(n375), .B2(n16), .ZN(n299) );
  OAI22_X1 U739 ( .A1(n18), .A2(n374), .B1(n373), .B2(n16), .ZN(n297) );
  OAI22_X1 U740 ( .A1(n18), .A2(n366), .B1(n365), .B2(n16), .ZN(n289) );
  XNOR2_X1 U741 ( .A(n586), .B(n420), .ZN(n386) );
  XNOR2_X1 U742 ( .A(n587), .B(n580), .ZN(n391) );
  XNOR2_X1 U743 ( .A(n586), .B(n424), .ZN(n390) );
  XNOR2_X1 U744 ( .A(n586), .B(n422), .ZN(n388) );
  XNOR2_X1 U745 ( .A(n586), .B(n423), .ZN(n389) );
  XNOR2_X1 U746 ( .A(n586), .B(n421), .ZN(n387) );
  XOR2_X1 U747 ( .A(n497), .B(n52), .Z(product[9]) );
  XNOR2_X1 U748 ( .A(n96), .B(n53), .ZN(product[8]) );
  OAI21_X1 U749 ( .B1(n64), .B2(n490), .A(n65), .ZN(n63) );
  OAI21_X1 U750 ( .B1(n540), .B2(n78), .A(n79), .ZN(n77) );
  OAI21_X1 U751 ( .B1(n540), .B2(n526), .A(n72), .ZN(n70) );
  XNOR2_X1 U752 ( .A(n528), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U753 ( .A(n529), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U754 ( .A(n528), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U755 ( .A(n528), .B(n418), .ZN(n401) );
  XNOR2_X1 U756 ( .A(n547), .B(n580), .ZN(n408) );
  XNOR2_X1 U757 ( .A(n529), .B(n420), .ZN(n403) );
  XNOR2_X1 U758 ( .A(n547), .B(n422), .ZN(n405) );
  XNOR2_X1 U759 ( .A(n546), .B(n419), .ZN(n402) );
  XNOR2_X1 U760 ( .A(n529), .B(n421), .ZN(n404) );
  XNOR2_X1 U761 ( .A(n529), .B(n424), .ZN(n407) );
  XNOR2_X1 U762 ( .A(n547), .B(n423), .ZN(n406) );
  OAI21_X1 U763 ( .B1(n107), .B2(n105), .A(n106), .ZN(n104) );
  XOR2_X1 U764 ( .A(n56), .B(n550), .Z(product[5]) );
  XOR2_X1 U765 ( .A(n58), .B(n115), .Z(product[3]) );
  OAI22_X1 U766 ( .A1(n525), .A2(n395), .B1(n394), .B2(n541), .ZN(n316) );
  OAI22_X1 U767 ( .A1(n524), .A2(n394), .B1(n393), .B2(n541), .ZN(n315) );
  OAI22_X1 U768 ( .A1(n524), .A2(n396), .B1(n395), .B2(n541), .ZN(n317) );
  OAI22_X1 U769 ( .A1(n525), .A2(n397), .B1(n396), .B2(n541), .ZN(n318) );
  OAI22_X1 U770 ( .A1(n524), .A2(n398), .B1(n397), .B2(n541), .ZN(n319) );
  OAI22_X1 U771 ( .A1(n524), .A2(n400), .B1(n399), .B2(n541), .ZN(n321) );
  OAI22_X1 U772 ( .A1(n525), .A2(n399), .B1(n398), .B2(n541), .ZN(n320) );
  OAI22_X1 U773 ( .A1(n401), .A2(n525), .B1(n400), .B2(n541), .ZN(n322) );
  OAI22_X1 U774 ( .A1(n6), .A2(n402), .B1(n401), .B2(n541), .ZN(n323) );
  NAND2_X1 U775 ( .A1(n329), .A2(n258), .ZN(n122) );
  OAI22_X1 U776 ( .A1(n6), .A2(n404), .B1(n403), .B2(n541), .ZN(n325) );
  OAI22_X1 U777 ( .A1(n524), .A2(n403), .B1(n402), .B2(n541), .ZN(n324) );
  OAI22_X1 U778 ( .A1(n524), .A2(n406), .B1(n405), .B2(n541), .ZN(n327) );
  OAI22_X1 U779 ( .A1(n6), .A2(n405), .B1(n404), .B2(n541), .ZN(n326) );
  OAI22_X1 U780 ( .A1(n525), .A2(n407), .B1(n406), .B2(n541), .ZN(n328) );
  OAI22_X1 U781 ( .A1(n525), .A2(n408), .B1(n407), .B2(n541), .ZN(n329) );
  OAI22_X1 U782 ( .A1(n524), .A2(n527), .B1(n409), .B2(n541), .ZN(n258) );
  OAI22_X1 U783 ( .A1(n12), .A2(n379), .B1(n378), .B2(n579), .ZN(n301) );
  OAI22_X1 U784 ( .A1(n499), .A2(n380), .B1(n379), .B2(n579), .ZN(n302) );
  OAI22_X1 U785 ( .A1(n561), .A2(n385), .B1(n384), .B2(n578), .ZN(n307) );
  OAI22_X1 U786 ( .A1(n561), .A2(n382), .B1(n381), .B2(n579), .ZN(n304) );
  OAI22_X1 U787 ( .A1(n12), .A2(n381), .B1(n380), .B2(n579), .ZN(n303) );
  NAND2_X1 U788 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U789 ( .A1(n532), .A2(n383), .B1(n382), .B2(n579), .ZN(n305) );
  OAI22_X1 U790 ( .A1(n499), .A2(n384), .B1(n383), .B2(n579), .ZN(n306) );
  OAI22_X1 U791 ( .A1(n561), .A2(n386), .B1(n385), .B2(n579), .ZN(n308) );
  OAI22_X1 U792 ( .A1(n562), .A2(n387), .B1(n386), .B2(n579), .ZN(n309) );
  OAI22_X1 U793 ( .A1(n562), .A2(n500), .B1(n392), .B2(n579), .ZN(n257) );
  OAI22_X1 U794 ( .A1(n532), .A2(n389), .B1(n388), .B2(n579), .ZN(n311) );
  OAI22_X1 U795 ( .A1(n12), .A2(n388), .B1(n387), .B2(n579), .ZN(n310) );
  OAI22_X1 U796 ( .A1(n499), .A2(n390), .B1(n389), .B2(n579), .ZN(n312) );
  INV_X1 U797 ( .A(n579), .ZN(n247) );
  OAI22_X1 U798 ( .A1(n562), .A2(n391), .B1(n390), .B2(n579), .ZN(n313) );
  INV_X1 U799 ( .A(n590), .ZN(n589) );
  INV_X1 U800 ( .A(n31), .ZN(n596) );
  INV_X1 U801 ( .A(n36), .ZN(n598) );
  INV_X1 U802 ( .A(n40), .ZN(n599) );
  XOR2_X1 U803 ( .A(n259), .B(n251), .Z(n148) );
  XOR2_X1 U804 ( .A(n149), .B(n147), .Z(n144) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_3_DW01_add_2 ( A, B, CI, SUM, 
        CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n19, n20, n21, n26, n27, n28, n34, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n49, n51, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n69, n71, n72, n73, n74, n75, n77, n79, n80,
         n81, n82, n83, n85, n87, n88, n90, n94, n99, n100, n102, n104, n161,
         n162, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189;

  OR2_X1 U126 ( .A1(A[14]), .A2(B[14]), .ZN(n161) );
  OR2_X1 U127 ( .A1(A[14]), .A2(B[14]), .ZN(n186) );
  OR2_X1 U128 ( .A1(A[8]), .A2(B[8]), .ZN(n162) );
  AND2_X1 U129 ( .A1(n180), .A2(n90), .ZN(SUM[0]) );
  XNOR2_X1 U130 ( .A(n41), .B(n164), .ZN(SUM[11]) );
  AND2_X1 U131 ( .A1(n189), .A2(n174), .ZN(n164) );
  AND2_X1 U132 ( .A1(A[14]), .A2(B[14]), .ZN(n165) );
  OR2_X1 U133 ( .A1(A[13]), .A2(B[13]), .ZN(n166) );
  AND2_X1 U134 ( .A1(A[13]), .A2(B[13]), .ZN(n167) );
  CLKBUF_X1 U135 ( .A(n28), .Z(n168) );
  OAI21_X1 U136 ( .B1(n36), .B2(n40), .A(n37), .ZN(n169) );
  INV_X1 U137 ( .A(n165), .ZN(n170) );
  INV_X1 U138 ( .A(n189), .ZN(n171) );
  AOI21_X1 U139 ( .B1(n34), .B2(n42), .A(n169), .ZN(n172) );
  NOR2_X1 U140 ( .A1(A[8]), .A2(B[8]), .ZN(n173) );
  NAND2_X1 U141 ( .A1(A[11]), .A2(B[11]), .ZN(n174) );
  NAND2_X1 U142 ( .A1(A[11]), .A2(B[11]), .ZN(n175) );
  NAND2_X1 U143 ( .A1(A[10]), .A2(B[10]), .ZN(n176) );
  AOI21_X1 U144 ( .B1(n42), .B2(n34), .A(n169), .ZN(n177) );
  OR2_X1 U145 ( .A1(A[10]), .A2(B[10]), .ZN(n178) );
  OR2_X1 U146 ( .A1(A[10]), .A2(B[10]), .ZN(n187) );
  NOR2_X1 U147 ( .A1(A[12]), .A2(B[12]), .ZN(n179) );
  NOR2_X1 U148 ( .A1(A[12]), .A2(B[12]), .ZN(n36) );
  OR2_X1 U149 ( .A1(A[0]), .A2(B[0]), .ZN(n180) );
  INV_X1 U150 ( .A(n64), .ZN(n63) );
  INV_X1 U151 ( .A(n55), .ZN(n54) );
  INV_X1 U152 ( .A(n42), .ZN(n41) );
  AOI21_X1 U153 ( .B1(n183), .B2(n72), .A(n69), .ZN(n67) );
  INV_X1 U154 ( .A(n71), .ZN(n69) );
  OAI21_X1 U155 ( .B1(n75), .B2(n73), .A(n74), .ZN(n72) );
  OAI21_X1 U156 ( .B1(n83), .B2(n81), .A(n82), .ZN(n80) );
  OAI21_X1 U157 ( .B1(n67), .B2(n65), .A(n66), .ZN(n64) );
  AOI21_X1 U158 ( .B1(n186), .B2(n167), .A(n165), .ZN(n21) );
  AOI21_X1 U159 ( .B1(n56), .B2(n64), .A(n57), .ZN(n55) );
  AOI21_X1 U160 ( .B1(n54), .B2(n181), .A(n51), .ZN(n49) );
  NAND2_X1 U161 ( .A1(n162), .A2(n59), .ZN(n8) );
  INV_X1 U162 ( .A(n90), .ZN(n88) );
  OAI21_X1 U163 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  INV_X1 U164 ( .A(n53), .ZN(n51) );
  AOI21_X1 U165 ( .B1(n182), .B2(n80), .A(n77), .ZN(n75) );
  INV_X1 U166 ( .A(n79), .ZN(n77) );
  AOI21_X1 U167 ( .B1(n184), .B2(n88), .A(n85), .ZN(n83) );
  INV_X1 U168 ( .A(n87), .ZN(n85) );
  NAND2_X1 U169 ( .A1(n100), .A2(n66), .ZN(n10) );
  INV_X1 U170 ( .A(n65), .ZN(n100) );
  NAND2_X1 U171 ( .A1(n102), .A2(n74), .ZN(n12) );
  INV_X1 U172 ( .A(n73), .ZN(n102) );
  NAND2_X1 U173 ( .A1(n181), .A2(n53), .ZN(n7) );
  NAND2_X1 U174 ( .A1(n99), .A2(n62), .ZN(n9) );
  INV_X1 U175 ( .A(n61), .ZN(n99) );
  NAND2_X1 U176 ( .A1(n104), .A2(n82), .ZN(n14) );
  INV_X1 U177 ( .A(n81), .ZN(n104) );
  NAND2_X1 U178 ( .A1(n183), .A2(n71), .ZN(n11) );
  NAND2_X1 U179 ( .A1(n182), .A2(n79), .ZN(n13) );
  NAND2_X1 U180 ( .A1(n184), .A2(n87), .ZN(n15) );
  XOR2_X1 U181 ( .A(n10), .B(n67), .Z(SUM[6]) );
  XNOR2_X1 U182 ( .A(n11), .B(n72), .ZN(SUM[5]) );
  XOR2_X1 U183 ( .A(n12), .B(n75), .Z(SUM[4]) );
  XOR2_X1 U184 ( .A(n14), .B(n83), .Z(SUM[2]) );
  XNOR2_X1 U185 ( .A(n15), .B(n88), .ZN(SUM[1]) );
  NAND2_X1 U186 ( .A1(n166), .A2(n28), .ZN(n3) );
  NOR2_X1 U187 ( .A1(A[7]), .A2(B[7]), .ZN(n61) );
  NOR2_X1 U188 ( .A1(A[8]), .A2(B[8]), .ZN(n58) );
  OR2_X1 U189 ( .A1(A[9]), .A2(B[9]), .ZN(n181) );
  NOR2_X1 U190 ( .A1(A[6]), .A2(B[6]), .ZN(n65) );
  NOR2_X1 U191 ( .A1(A[4]), .A2(B[4]), .ZN(n73) );
  NOR2_X1 U192 ( .A1(A[2]), .A2(B[2]), .ZN(n81) );
  NAND2_X1 U193 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  XOR2_X1 U194 ( .A(n49), .B(n6), .Z(SUM[10]) );
  NAND2_X1 U195 ( .A1(A[11]), .A2(B[11]), .ZN(n40) );
  OR2_X1 U196 ( .A1(A[3]), .A2(B[3]), .ZN(n182) );
  OR2_X1 U197 ( .A1(A[5]), .A2(B[5]), .ZN(n183) );
  OR2_X1 U198 ( .A1(A[1]), .A2(B[1]), .ZN(n184) );
  OR2_X1 U199 ( .A1(n17), .A2(n185), .ZN(n1) );
  AND2_X1 U200 ( .A1(A[15]), .A2(B[15]), .ZN(n185) );
  XNOR2_X1 U201 ( .A(n60), .B(n8), .ZN(SUM[8]) );
  XNOR2_X1 U202 ( .A(n54), .B(n7), .ZN(SUM[9]) );
  XNOR2_X1 U203 ( .A(n13), .B(n80), .ZN(SUM[3]) );
  NAND2_X1 U204 ( .A1(A[7]), .A2(B[7]), .ZN(n62) );
  NAND2_X1 U205 ( .A1(A[4]), .A2(B[4]), .ZN(n74) );
  NAND2_X1 U206 ( .A1(A[6]), .A2(B[6]), .ZN(n66) );
  NAND2_X1 U207 ( .A1(A[2]), .A2(B[2]), .ZN(n82) );
  NAND2_X1 U208 ( .A1(A[3]), .A2(B[3]), .ZN(n79) );
  NAND2_X1 U209 ( .A1(A[5]), .A2(B[5]), .ZN(n71) );
  NAND2_X1 U210 ( .A1(A[1]), .A2(B[1]), .ZN(n87) );
  NAND2_X1 U211 ( .A1(A[0]), .A2(B[0]), .ZN(n90) );
  XOR2_X1 U212 ( .A(n63), .B(n9), .Z(SUM[7]) );
  NAND2_X1 U213 ( .A1(n94), .A2(n37), .ZN(n4) );
  INV_X1 U214 ( .A(n179), .ZN(n94) );
  AND2_X1 U215 ( .A1(A[10]), .A2(B[10]), .ZN(n188) );
  OR2_X1 U216 ( .A1(A[11]), .A2(B[11]), .ZN(n189) );
  NOR2_X1 U217 ( .A1(A[11]), .A2(B[11]), .ZN(n39) );
  NOR2_X1 U218 ( .A1(n173), .A2(n61), .ZN(n56) );
  OAI21_X1 U219 ( .B1(n58), .B2(n62), .A(n59), .ZN(n57) );
  NAND2_X1 U220 ( .A1(A[8]), .A2(B[8]), .ZN(n59) );
  NAND2_X1 U221 ( .A1(n161), .A2(n170), .ZN(n2) );
  NAND2_X1 U222 ( .A1(A[12]), .A2(B[12]), .ZN(n37) );
  NAND2_X1 U223 ( .A1(A[9]), .A2(B[9]), .ZN(n53) );
  XNOR2_X1 U224 ( .A(n19), .B(n1), .ZN(SUM[15]) );
  OAI21_X1 U225 ( .B1(n41), .B2(n171), .A(n175), .ZN(n38) );
  NOR2_X1 U226 ( .A1(A[13]), .A2(B[13]), .ZN(n27) );
  NOR2_X1 U227 ( .A1(n179), .A2(n39), .ZN(n34) );
  NOR2_X1 U228 ( .A1(A[15]), .A2(B[15]), .ZN(n17) );
  NAND2_X1 U229 ( .A1(n178), .A2(n176), .ZN(n6) );
  OAI21_X1 U230 ( .B1(n43), .B2(n55), .A(n44), .ZN(n42) );
  NAND2_X1 U231 ( .A1(n178), .A2(n181), .ZN(n43) );
  AOI21_X1 U232 ( .B1(n187), .B2(n51), .A(n188), .ZN(n44) );
  XNOR2_X1 U233 ( .A(n38), .B(n4), .ZN(SUM[12]) );
  NAND2_X1 U234 ( .A1(n161), .A2(n166), .ZN(n20) );
  XNOR2_X1 U235 ( .A(n26), .B(n2), .ZN(SUM[14]) );
  XOR2_X1 U236 ( .A(n172), .B(n3), .Z(SUM[13]) );
  OAI21_X1 U237 ( .B1(n177), .B2(n27), .A(n168), .ZN(n26) );
  OAI21_X1 U238 ( .B1(n172), .B2(n20), .A(n21), .ZN(n19) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_3 ( clk, clear_acc, 
        data_out_x, data_out, data_out_w, data_out_b, wr_en_y, m_valid, 
        m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [3:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N27, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, n1, n2, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n87, n104, n113, n114, n115, n116, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n15), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n221), .CK(clk), .Q(n20) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n222), .CK(clk), .Q(n21) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n223), .CK(clk), .Q(n22) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n224), .CK(clk), .Q(n23) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n225), .CK(clk), .Q(n24) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n226), .CK(clk), .Q(n25) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n227), .CK(clk), .Q(n26) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n228), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n229), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n230), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n231), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n232), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n233), .CK(clk), .Q(n34) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n234), .CK(clk), .Q(n35) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n235), .CK(clk), .Q(n36) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n236), .CK(clk), .Q(n38) );
  DFF_X1 \f_reg[7]  ( .D(n81), .CK(clk), .Q(f[7]), .QN(n213) );
  DFF_X1 \f_reg[8]  ( .D(n80), .CK(clk), .Q(f[8]), .QN(n214) );
  DFF_X1 \f_reg[9]  ( .D(n79), .CK(clk), .Q(f[9]), .QN(n215) );
  DFF_X1 \f_reg[10]  ( .D(n78), .CK(clk), .Q(n49), .QN(n216) );
  DFF_X1 \f_reg[11]  ( .D(n77), .CK(clk), .Q(n47), .QN(n217) );
  DFF_X1 \f_reg[12]  ( .D(n76), .CK(clk), .Q(n45), .QN(n218) );
  DFF_X1 \f_reg[14]  ( .D(n5), .CK(clk), .Q(n43), .QN(n220) );
  DFF_X1 \f_reg[15]  ( .D(n75), .CK(clk), .Q(f[15]), .QN(n73) );
  DFF_X1 \data_out_reg[15]  ( .D(n114), .CK(clk), .Q(data_out[15]), .QN(n193)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n115), .CK(clk), .Q(data_out[14]), .QN(n192)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n116), .CK(clk), .Q(data_out[13]), .QN(n191)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n165), .CK(clk), .Q(data_out[12]), .QN(n190)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n166), .CK(clk), .Q(data_out[11]), .QN(n189)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n167), .CK(clk), .Q(data_out[10]), .QN(n188)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n168), .CK(clk), .Q(data_out[9]), .QN(n187) );
  DFF_X1 \data_out_reg[8]  ( .D(n169), .CK(clk), .Q(data_out[8]), .QN(n186) );
  DFF_X1 \data_out_reg[7]  ( .D(n170), .CK(clk), .Q(data_out[7]), .QN(n185) );
  DFF_X1 \data_out_reg[6]  ( .D(n171), .CK(clk), .Q(data_out[6]), .QN(n184) );
  DFF_X1 \data_out_reg[5]  ( .D(n172), .CK(clk), .Q(data_out[5]), .QN(n183) );
  DFF_X1 \data_out_reg[4]  ( .D(n173), .CK(clk), .Q(data_out[4]), .QN(n182) );
  DFF_X1 \data_out_reg[3]  ( .D(n174), .CK(clk), .Q(data_out[3]), .QN(n181) );
  DFF_X1 \data_out_reg[2]  ( .D(n175), .CK(clk), .Q(data_out[2]), .QN(n180) );
  DFF_X1 \data_out_reg[1]  ( .D(n176), .CK(clk), .Q(data_out[1]), .QN(n179) );
  DFF_X1 \data_out_reg[0]  ( .D(n177), .CK(clk), .Q(data_out[0]), .QN(n178) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_3_DW_mult_tc_1 mult_960 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_3_DW01_add_2 add_961 ( .A({n200, 
        n199, n198, n197, n196, n195, n209, n208, n207, n206, n205, n204, n203, 
        n202, n201, n194}), .B({f[15], n43, n44, n45, n47, n49, f[9:3], n57, 
        n59, n61}), .CI(1'b0), .SUM(adder) );
  DFF_X2 delay_reg ( .D(N27), .CK(clk), .Q(n12), .QN(n237) );
  DFF_X1 \f_reg[3]  ( .D(n85), .CK(clk), .Q(f[3]), .QN(n65) );
  DFF_X1 \f_reg[4]  ( .D(n84), .CK(clk), .Q(f[4]), .QN(n66) );
  DFF_X1 \f_reg[2]  ( .D(n87), .CK(clk), .Q(n57), .QN(n212) );
  DFF_X1 \f_reg[1]  ( .D(n104), .CK(clk), .Q(n59), .QN(n211) );
  DFF_X1 \f_reg[0]  ( .D(n113), .CK(clk), .Q(n61), .QN(n210) );
  DFF_X1 \f_reg[5]  ( .D(n83), .CK(clk), .Q(f[5]), .QN(n67) );
  DFF_X1 \f_reg[6]  ( .D(n82), .CK(clk), .Q(f[6]), .QN(n68) );
  DFF_X2 \f_reg[13]  ( .D(n4), .CK(clk), .Q(n44), .QN(n219) );
  AND2_X2 U3 ( .A1(n41), .A2(n16), .ZN(n13) );
  AND2_X1 U4 ( .A1(n63), .A2(f[15]), .ZN(n1) );
  AND2_X1 U5 ( .A1(data_out_b[15]), .A2(n15), .ZN(n2) );
  NAND3_X1 U6 ( .A1(n7), .A2(n6), .A3(n8), .ZN(n4) );
  NAND3_X1 U8 ( .A1(n10), .A2(n9), .A3(n11), .ZN(n5) );
  MUX2_X2 U9 ( .A(N43), .B(n21), .S(n12), .Z(n199) );
  MUX2_X2 U10 ( .A(n27), .B(N37), .S(n237), .Z(n208) );
  MUX2_X2 U11 ( .A(n26), .B(N38), .S(n237), .Z(n209) );
  NAND2_X1 U12 ( .A1(data_out_b[13]), .A2(n15), .ZN(n6) );
  NAND2_X1 U13 ( .A1(adder[13]), .A2(n13), .ZN(n7) );
  NAND2_X1 U14 ( .A1(n63), .A2(n44), .ZN(n8) );
  AOI211_X1 U15 ( .C1(adder[15]), .C2(n13), .A(n1), .B(n2), .ZN(n42) );
  MUX2_X2 U16 ( .A(n24), .B(N40), .S(n237), .Z(n196) );
  MUX2_X2 U17 ( .A(n22), .B(N42), .S(n237), .Z(n198) );
  NAND2_X1 U18 ( .A1(data_out_b[14]), .A2(n15), .ZN(n9) );
  NAND2_X1 U19 ( .A1(adder[14]), .A2(n13), .ZN(n10) );
  NAND2_X1 U20 ( .A1(n63), .A2(n43), .ZN(n11) );
  INV_X2 U21 ( .A(n41), .ZN(n63) );
  MUX2_X2 U22 ( .A(N39), .B(n25), .S(n12), .Z(n195) );
  MUX2_X2 U23 ( .A(n23), .B(N41), .S(n237), .Z(n197) );
  INV_X1 U24 ( .A(n16), .ZN(n15) );
  INV_X1 U25 ( .A(clear_acc), .ZN(n16) );
  NAND2_X1 U26 ( .A1(n14), .A2(N27), .ZN(n239) );
  INV_X1 U27 ( .A(n19), .ZN(n37) );
  OAI22_X1 U28 ( .A1(n181), .A2(n239), .B1(n65), .B2(n238), .ZN(n174) );
  OAI22_X1 U29 ( .A1(n182), .A2(n239), .B1(n66), .B2(n238), .ZN(n173) );
  OAI22_X1 U30 ( .A1(n183), .A2(n239), .B1(n67), .B2(n238), .ZN(n172) );
  OAI22_X1 U31 ( .A1(n184), .A2(n239), .B1(n68), .B2(n238), .ZN(n171) );
  OAI22_X1 U32 ( .A1(n185), .A2(n239), .B1(n213), .B2(n238), .ZN(n170) );
  OAI22_X1 U33 ( .A1(n186), .A2(n239), .B1(n214), .B2(n238), .ZN(n169) );
  OAI22_X1 U34 ( .A1(n187), .A2(n239), .B1(n215), .B2(n238), .ZN(n168) );
  MUX2_X1 U35 ( .A(n20), .B(N44), .S(n237), .Z(n200) );
  INV_X1 U36 ( .A(wr_en_y), .ZN(n14) );
  AND2_X1 U37 ( .A1(sel[0]), .A2(sel[1]), .ZN(n18) );
  INV_X1 U38 ( .A(m_ready), .ZN(n17) );
  NAND2_X1 U39 ( .A1(m_valid), .A2(n17), .ZN(n39) );
  OAI211_X1 U40 ( .C1(sel[2]), .C2(n18), .A(sel[3]), .B(n39), .ZN(N27) );
  NAND2_X1 U41 ( .A1(clear_acc_delay), .A2(n237), .ZN(n19) );
  MUX2_X1 U42 ( .A(n20), .B(N44), .S(n37), .Z(n221) );
  MUX2_X1 U43 ( .A(n21), .B(N43), .S(n37), .Z(n222) );
  MUX2_X1 U44 ( .A(n22), .B(N42), .S(n37), .Z(n223) );
  MUX2_X1 U45 ( .A(n23), .B(N41), .S(n37), .Z(n224) );
  MUX2_X1 U46 ( .A(n24), .B(N40), .S(n37), .Z(n225) );
  MUX2_X1 U47 ( .A(n25), .B(N39), .S(n37), .Z(n226) );
  MUX2_X1 U48 ( .A(n26), .B(N38), .S(n37), .Z(n227) );
  MUX2_X1 U49 ( .A(n27), .B(N37), .S(n37), .Z(n228) );
  MUX2_X1 U50 ( .A(n28), .B(N36), .S(n37), .Z(n229) );
  MUX2_X1 U51 ( .A(n28), .B(N36), .S(n237), .Z(n207) );
  MUX2_X1 U52 ( .A(n29), .B(N35), .S(n37), .Z(n230) );
  MUX2_X1 U53 ( .A(n29), .B(N35), .S(n237), .Z(n206) );
  MUX2_X1 U54 ( .A(n32), .B(N34), .S(n37), .Z(n231) );
  MUX2_X1 U55 ( .A(n32), .B(N34), .S(n237), .Z(n205) );
  MUX2_X1 U56 ( .A(n33), .B(N33), .S(n37), .Z(n232) );
  MUX2_X1 U57 ( .A(n33), .B(N33), .S(n237), .Z(n204) );
  MUX2_X1 U58 ( .A(n34), .B(N32), .S(n37), .Z(n233) );
  MUX2_X1 U59 ( .A(n34), .B(N32), .S(n237), .Z(n203) );
  MUX2_X1 U60 ( .A(n35), .B(N31), .S(n37), .Z(n234) );
  MUX2_X1 U61 ( .A(n35), .B(N31), .S(n237), .Z(n202) );
  MUX2_X1 U62 ( .A(n36), .B(N30), .S(n37), .Z(n235) );
  MUX2_X1 U63 ( .A(n36), .B(N30), .S(n237), .Z(n201) );
  MUX2_X1 U64 ( .A(n38), .B(N29), .S(n37), .Z(n236) );
  MUX2_X1 U65 ( .A(n38), .B(N29), .S(n237), .Z(n194) );
  INV_X1 U66 ( .A(n39), .ZN(n40) );
  OAI21_X1 U67 ( .B1(n40), .B2(n12), .A(n16), .ZN(n41) );
  INV_X1 U68 ( .A(n42), .ZN(n75) );
  AOI222_X1 U69 ( .A1(data_out_b[12]), .A2(n15), .B1(adder[12]), .B2(n13), 
        .C1(n63), .C2(n45), .ZN(n46) );
  INV_X1 U70 ( .A(n46), .ZN(n76) );
  AOI222_X1 U71 ( .A1(data_out_b[11]), .A2(n15), .B1(adder[11]), .B2(n13), 
        .C1(n63), .C2(n47), .ZN(n48) );
  INV_X1 U72 ( .A(n48), .ZN(n77) );
  AOI222_X1 U73 ( .A1(data_out_b[10]), .A2(n15), .B1(adder[10]), .B2(n13), 
        .C1(n63), .C2(n49), .ZN(n50) );
  INV_X1 U74 ( .A(n50), .ZN(n78) );
  AOI222_X1 U75 ( .A1(data_out_b[8]), .A2(n15), .B1(adder[8]), .B2(n13), .C1(
        n63), .C2(f[8]), .ZN(n51) );
  INV_X1 U76 ( .A(n51), .ZN(n80) );
  AOI222_X1 U77 ( .A1(data_out_b[7]), .A2(n15), .B1(adder[7]), .B2(n13), .C1(
        n63), .C2(f[7]), .ZN(n52) );
  INV_X1 U78 ( .A(n52), .ZN(n81) );
  AOI222_X1 U79 ( .A1(data_out_b[6]), .A2(n15), .B1(adder[6]), .B2(n13), .C1(
        n63), .C2(f[6]), .ZN(n53) );
  INV_X1 U80 ( .A(n53), .ZN(n82) );
  AOI222_X1 U81 ( .A1(data_out_b[5]), .A2(n15), .B1(adder[5]), .B2(n13), .C1(
        n63), .C2(f[5]), .ZN(n54) );
  INV_X1 U82 ( .A(n54), .ZN(n83) );
  AOI222_X1 U83 ( .A1(data_out_b[4]), .A2(n15), .B1(adder[4]), .B2(n13), .C1(
        n63), .C2(f[4]), .ZN(n55) );
  INV_X1 U84 ( .A(n55), .ZN(n84) );
  AOI222_X1 U85 ( .A1(data_out_b[3]), .A2(n15), .B1(adder[3]), .B2(n13), .C1(
        n63), .C2(f[3]), .ZN(n56) );
  INV_X1 U86 ( .A(n56), .ZN(n85) );
  AOI222_X1 U87 ( .A1(data_out_b[2]), .A2(n15), .B1(adder[2]), .B2(n13), .C1(
        n63), .C2(n57), .ZN(n58) );
  INV_X1 U88 ( .A(n58), .ZN(n87) );
  AOI222_X1 U89 ( .A1(data_out_b[1]), .A2(n15), .B1(adder[1]), .B2(n13), .C1(
        n63), .C2(n59), .ZN(n60) );
  INV_X1 U90 ( .A(n60), .ZN(n104) );
  AOI222_X1 U91 ( .A1(data_out_b[0]), .A2(n15), .B1(adder[0]), .B2(n13), .C1(
        n63), .C2(n61), .ZN(n62) );
  INV_X1 U92 ( .A(n62), .ZN(n113) );
  AOI222_X1 U93 ( .A1(data_out_b[9]), .A2(n15), .B1(adder[9]), .B2(n13), .C1(
        n63), .C2(f[9]), .ZN(n64) );
  INV_X1 U94 ( .A(n64), .ZN(n79) );
  NOR4_X1 U95 ( .A1(n47), .A2(n45), .A3(n44), .A4(n43), .ZN(n72) );
  NOR4_X1 U96 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n49), .ZN(n71) );
  NAND4_X1 U97 ( .A1(n68), .A2(n67), .A3(n66), .A4(n65), .ZN(n69) );
  NOR4_X1 U98 ( .A1(n69), .A2(n61), .A3(n59), .A4(n57), .ZN(n70) );
  NAND3_X1 U99 ( .A1(n72), .A2(n71), .A3(n70), .ZN(n74) );
  NAND3_X1 U100 ( .A1(wr_en_y), .A2(n74), .A3(n73), .ZN(n238) );
  OAI22_X1 U101 ( .A1(n178), .A2(n239), .B1(n210), .B2(n238), .ZN(n177) );
  OAI22_X1 U102 ( .A1(n179), .A2(n239), .B1(n211), .B2(n238), .ZN(n176) );
  OAI22_X1 U103 ( .A1(n180), .A2(n239), .B1(n212), .B2(n238), .ZN(n175) );
  OAI22_X1 U104 ( .A1(n188), .A2(n239), .B1(n216), .B2(n238), .ZN(n167) );
  OAI22_X1 U105 ( .A1(n189), .A2(n239), .B1(n217), .B2(n238), .ZN(n166) );
  OAI22_X1 U106 ( .A1(n190), .A2(n239), .B1(n218), .B2(n238), .ZN(n165) );
  OAI22_X1 U107 ( .A1(n191), .A2(n239), .B1(n219), .B2(n238), .ZN(n116) );
  OAI22_X1 U108 ( .A1(n192), .A2(n239), .B1(n220), .B2(n238), .ZN(n115) );
  OAI22_X1 U109 ( .A1(n193), .A2(n239), .B1(n73), .B2(n238), .ZN(n114) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_2_DW_mult_tc_1 ( a, b, 
        product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n9, n12, n13, n16, n18, n19, n23, n25, n29, n31, n32, n34,
         n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n50, n53, n54,
         n55, n56, n57, n58, n59, n62, n63, n64, n65, n67, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n95, n96, n97, n98, n99, n101, n103, n104,
         n105, n106, n107, n111, n112, n113, n114, n115, n117, n119, n120,
         n122, n125, n127, n131, n133, n135, n139, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n247, n249, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n418, n419,
         n420, n421, n422, n423, n424, n426, n427, n429, n432, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U148 ( .A(n265), .B(n144), .Z(n145) );
  XOR2_X1 U150 ( .A(n271), .B(n146), .Z(n147) );
  XOR2_X1 U152 ( .A(n301), .B(n148), .Z(n149) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U161 ( .A(n177), .B(n168), .CI(n166), .CO(n163), .S(n164) );
  FA_X1 U162 ( .A(n170), .B(n172), .CI(n179), .CO(n165), .S(n166) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n263), .CI(n291), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n317), .B(n252), .CO(n173), .S(n174) );
  FA_X1 U167 ( .A(n180), .B(n187), .CI(n178), .CO(n175), .S(n176) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U169 ( .A(n193), .B(n282), .CI(n191), .CO(n179), .S(n180) );
  FA_X1 U170 ( .A(n268), .B(n292), .CI(n274), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U172 ( .A(n197), .B(n190), .CI(n188), .CO(n185), .S(n186) );
  FA_X1 U173 ( .A(n199), .B(n201), .CI(n192), .CO(n187), .S(n188) );
  FA_X1 U174 ( .A(n293), .B(n275), .CI(n194), .CO(n189), .S(n190) );
  FA_X1 U175 ( .A(n253), .B(n283), .CI(n305), .CO(n191), .S(n192) );
  HA_X1 U176 ( .A(n319), .B(n269), .CO(n193), .S(n194) );
  FA_X1 U177 ( .A(n205), .B(n200), .CI(n198), .CO(n195), .S(n196) );
  FA_X1 U178 ( .A(n209), .B(n207), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U179 ( .A(n276), .B(n284), .CI(n294), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n320), .B(n270), .CI(n306), .CO(n201), .S(n202) );
  FA_X1 U182 ( .A(n210), .B(n307), .CI(n215), .CO(n205), .S(n206) );
  FA_X1 U183 ( .A(n285), .B(n254), .CI(n295), .CO(n207), .S(n208) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U185 ( .A(n216), .B(n219), .CI(n214), .CO(n211), .S(n212) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n322), .B(n278), .CI(n308), .CO(n215), .S(n216) );
  FA_X1 U188 ( .A(n225), .B(n222), .CI(n220), .CO(n217), .S(n218) );
  FA_X1 U189 ( .A(n255), .B(n309), .CI(n297), .CO(n219), .S(n220) );
  HA_X1 U190 ( .A(n287), .B(n323), .CO(n221), .S(n222) );
  FA_X1 U192 ( .A(n324), .B(n288), .CI(n310), .CO(n225), .S(n226) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  HA_X1 U194 ( .A(n311), .B(n325), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n312), .B(n300), .CI(n326), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  BUF_X1 U414 ( .A(n498), .Z(n508) );
  AND2_X1 U415 ( .A1(n212), .A2(n217), .ZN(n490) );
  BUF_X2 U416 ( .A(n570), .Z(n512) );
  BUF_X1 U417 ( .A(n570), .Z(n511) );
  CLKBUF_X3 U418 ( .A(n9), .Z(n567) );
  BUF_X1 U419 ( .A(n509), .Z(n491) );
  BUF_X1 U420 ( .A(n498), .Z(n509) );
  XOR2_X1 U421 ( .A(n526), .B(a[8]), .Z(n492) );
  OR2_X1 U422 ( .A1(n329), .A2(n258), .ZN(n493) );
  OR2_X1 U423 ( .A1(n529), .A2(n548), .ZN(n18) );
  INV_X1 U424 ( .A(n548), .ZN(n16) );
  INV_X1 U425 ( .A(n577), .ZN(n576) );
  BUF_X1 U426 ( .A(n23), .Z(n506) );
  XOR2_X1 U427 ( .A(n577), .B(a[4]), .Z(n529) );
  OR2_X2 U428 ( .A1(n527), .A2(n555), .ZN(n497) );
  BUF_X2 U429 ( .A(n570), .Z(n513) );
  OR2_X2 U430 ( .A1(n538), .A2(n249), .ZN(n539) );
  XOR2_X1 U431 ( .A(n578), .B(a[8]), .Z(n494) );
  XNOR2_X1 U432 ( .A(n580), .B(a[8]), .ZN(n429) );
  INV_X1 U433 ( .A(n573), .ZN(n495) );
  OR2_X1 U434 ( .A1(n527), .A2(n555), .ZN(n496) );
  OR2_X1 U435 ( .A1(n527), .A2(n555), .ZN(n23) );
  XOR2_X1 U436 ( .A(n577), .B(a[6]), .Z(n498) );
  CLKBUF_X1 U437 ( .A(n96), .Z(n499) );
  INV_X1 U438 ( .A(n576), .ZN(n500) );
  CLKBUF_X1 U439 ( .A(n505), .Z(n541) );
  XNOR2_X1 U440 ( .A(n45), .B(n501), .ZN(product[12]) );
  AND2_X1 U441 ( .A1(n504), .A2(n79), .ZN(n501) );
  NAND2_X1 U442 ( .A1(n429), .A2(n507), .ZN(n502) );
  XNOR2_X1 U443 ( .A(n541), .B(n503), .ZN(product[9]) );
  AND2_X1 U444 ( .A1(n537), .A2(n90), .ZN(n503) );
  OR2_X1 U445 ( .A1(n176), .A2(n185), .ZN(n504) );
  AOI21_X1 U446 ( .B1(n96), .B2(n557), .A(n490), .ZN(n505) );
  AOI21_X1 U447 ( .B1(n96), .B2(n557), .A(n490), .ZN(n91) );
  INV_X2 U448 ( .A(n584), .ZN(n583) );
  BUF_X4 U449 ( .A(n19), .Z(n526) );
  OR2_X2 U450 ( .A1(n529), .A2(n548), .ZN(n530) );
  XOR2_X1 U451 ( .A(n571), .B(a[2]), .Z(n9) );
  XNOR2_X1 U452 ( .A(n526), .B(a[8]), .ZN(n507) );
  INV_X2 U453 ( .A(n574), .ZN(n572) );
  INV_X1 U454 ( .A(n519), .ZN(n37) );
  BUF_X1 U455 ( .A(n498), .Z(n510) );
  INV_X1 U456 ( .A(n571), .ZN(n570) );
  NOR2_X1 U457 ( .A1(n164), .A2(n175), .ZN(n514) );
  NOR2_X1 U458 ( .A1(n164), .A2(n175), .ZN(n75) );
  NAND2_X1 U459 ( .A1(n432), .A2(n566), .ZN(n515) );
  CLKBUF_X1 U460 ( .A(n104), .Z(n516) );
  OAI21_X1 U461 ( .B1(n105), .B2(n107), .A(n106), .ZN(n104) );
  NAND2_X1 U462 ( .A1(n196), .A2(n203), .ZN(n517) );
  OAI21_X1 U463 ( .B1(n505), .B2(n89), .A(n90), .ZN(n518) );
  OAI21_X1 U464 ( .B1(n91), .B2(n89), .A(n90), .ZN(n88) );
  XNOR2_X1 U465 ( .A(n582), .B(a[12]), .ZN(n519) );
  INV_X1 U466 ( .A(n582), .ZN(n581) );
  CLKBUF_X1 U467 ( .A(n105), .Z(n520) );
  NOR2_X1 U468 ( .A1(n186), .A2(n195), .ZN(n521) );
  NOR2_X1 U469 ( .A1(n186), .A2(n195), .ZN(n82) );
  XOR2_X1 U470 ( .A(n582), .B(a[10]), .Z(n523) );
  BUF_X2 U471 ( .A(n9), .Z(n566) );
  XNOR2_X1 U472 ( .A(n518), .B(n522), .ZN(product[10]) );
  NAND2_X1 U473 ( .A1(n525), .A2(n517), .ZN(n522) );
  OR2_X2 U474 ( .A1(n523), .A2(n540), .ZN(n34) );
  INV_X1 U475 ( .A(n492), .ZN(n524) );
  OR2_X1 U476 ( .A1(n196), .A2(n203), .ZN(n525) );
  XOR2_X1 U477 ( .A(n578), .B(a[6]), .Z(n527) );
  NAND2_X1 U478 ( .A1(n429), .A2(n507), .ZN(n29) );
  AOI21_X1 U479 ( .B1(n80), .B2(n518), .A(n81), .ZN(n528) );
  AOI21_X1 U480 ( .B1(n80), .B2(n88), .A(n81), .ZN(n45) );
  CLKBUF_X1 U481 ( .A(n112), .Z(n531) );
  INV_X1 U482 ( .A(n532), .ZN(n111) );
  AND2_X1 U483 ( .A1(n232), .A2(n233), .ZN(n532) );
  XOR2_X1 U484 ( .A(n208), .B(n213), .Z(n533) );
  XOR2_X1 U485 ( .A(n206), .B(n533), .Z(n204) );
  NAND2_X1 U486 ( .A1(n206), .A2(n208), .ZN(n534) );
  NAND2_X1 U487 ( .A1(n206), .A2(n213), .ZN(n535) );
  NAND2_X1 U488 ( .A1(n208), .A2(n213), .ZN(n536) );
  NAND3_X1 U489 ( .A1(n534), .A2(n535), .A3(n536), .ZN(n203) );
  XNOR2_X1 U490 ( .A(n574), .B(a[2]), .ZN(n432) );
  OR2_X1 U491 ( .A1(n204), .A2(n211), .ZN(n537) );
  OR2_X1 U492 ( .A1(n538), .A2(n249), .ZN(n6) );
  XNOR2_X1 U493 ( .A(n1), .B(n249), .ZN(n538) );
  INV_X1 U494 ( .A(n540), .ZN(n32) );
  XNOR2_X1 U495 ( .A(n580), .B(a[10]), .ZN(n540) );
  NAND2_X1 U496 ( .A1(n432), .A2(n566), .ZN(n542) );
  NAND2_X1 U497 ( .A1(n432), .A2(n566), .ZN(n543) );
  NAND2_X1 U498 ( .A1(n432), .A2(n566), .ZN(n12) );
  AOI21_X1 U499 ( .B1(n558), .B2(n516), .A(n101), .ZN(n544) );
  CLKBUF_X1 U500 ( .A(n107), .Z(n545) );
  INV_X1 U501 ( .A(n249), .ZN(n546) );
  INV_X1 U502 ( .A(n249), .ZN(n547) );
  XNOR2_X1 U503 ( .A(n574), .B(a[4]), .ZN(n548) );
  XNOR2_X1 U504 ( .A(n226), .B(n549), .ZN(n224) );
  XNOR2_X1 U505 ( .A(n229), .B(n298), .ZN(n549) );
  NAND2_X1 U506 ( .A1(n226), .A2(n229), .ZN(n550) );
  NAND2_X1 U507 ( .A1(n226), .A2(n298), .ZN(n551) );
  NAND2_X1 U508 ( .A1(n229), .A2(n298), .ZN(n552) );
  NAND3_X1 U509 ( .A1(n550), .A2(n551), .A3(n552), .ZN(n223) );
  OR2_X1 U510 ( .A1(n6), .A2(n403), .ZN(n553) );
  OR2_X1 U511 ( .A1(n402), .A2(n547), .ZN(n554) );
  NAND2_X1 U512 ( .A1(n553), .A2(n554), .ZN(n324) );
  INV_X2 U513 ( .A(n580), .ZN(n579) );
  XNOR2_X1 U514 ( .A(n577), .B(a[6]), .ZN(n555) );
  NAND2_X1 U515 ( .A1(n556), .A2(n69), .ZN(n47) );
  INV_X1 U516 ( .A(n73), .ZN(n71) );
  AOI21_X1 U517 ( .B1(n556), .B2(n74), .A(n67), .ZN(n65) );
  INV_X1 U518 ( .A(n69), .ZN(n67) );
  INV_X1 U519 ( .A(n74), .ZN(n72) );
  NOR2_X1 U520 ( .A1(n75), .A2(n78), .ZN(n73) );
  XNOR2_X1 U521 ( .A(n84), .B(n50), .ZN(product[11]) );
  NAND2_X1 U522 ( .A1(n127), .A2(n83), .ZN(n50) );
  OR2_X1 U523 ( .A1(n152), .A2(n163), .ZN(n556) );
  OAI21_X1 U524 ( .B1(n514), .B2(n79), .A(n76), .ZN(n74) );
  NAND2_X1 U525 ( .A1(n125), .A2(n76), .ZN(n48) );
  INV_X1 U526 ( .A(n75), .ZN(n125) );
  NAND2_X1 U527 ( .A1(n152), .A2(n163), .ZN(n69) );
  NAND2_X1 U528 ( .A1(n557), .A2(n95), .ZN(n53) );
  INV_X1 U529 ( .A(n103), .ZN(n101) );
  OAI21_X1 U530 ( .B1(n115), .B2(n113), .A(n114), .ZN(n112) );
  NAND2_X1 U531 ( .A1(n133), .A2(n106), .ZN(n56) );
  INV_X1 U532 ( .A(n520), .ZN(n133) );
  NAND2_X1 U533 ( .A1(n131), .A2(n98), .ZN(n54) );
  INV_X1 U534 ( .A(n97), .ZN(n131) );
  AOI21_X1 U535 ( .B1(n560), .B2(n120), .A(n117), .ZN(n115) );
  INV_X1 U536 ( .A(n119), .ZN(n117) );
  XOR2_X1 U537 ( .A(n58), .B(n115), .Z(product[3]) );
  INV_X1 U538 ( .A(n113), .ZN(n135) );
  NOR2_X1 U539 ( .A1(n196), .A2(n203), .ZN(n85) );
  XNOR2_X1 U540 ( .A(n55), .B(n516), .ZN(product[6]) );
  NAND2_X1 U541 ( .A1(n558), .A2(n103), .ZN(n55) );
  XNOR2_X1 U542 ( .A(n57), .B(n531), .ZN(product[4]) );
  NAND2_X1 U543 ( .A1(n559), .A2(n111), .ZN(n57) );
  NAND2_X1 U544 ( .A1(n186), .A2(n195), .ZN(n83) );
  NAND2_X1 U545 ( .A1(n176), .A2(n185), .ZN(n79) );
  NAND2_X1 U546 ( .A1(n164), .A2(n175), .ZN(n76) );
  NAND2_X1 U547 ( .A1(n196), .A2(n203), .ZN(n86) );
  NAND2_X1 U548 ( .A1(n212), .A2(n217), .ZN(n95) );
  OR2_X1 U549 ( .A1(n212), .A2(n217), .ZN(n557) );
  XNOR2_X1 U550 ( .A(n59), .B(n120), .ZN(product[2]) );
  NAND2_X1 U551 ( .A1(n560), .A2(n119), .ZN(n59) );
  NAND2_X1 U552 ( .A1(n561), .A2(n62), .ZN(n46) );
  NAND2_X1 U553 ( .A1(n73), .A2(n556), .ZN(n64) );
  INV_X1 U554 ( .A(n577), .ZN(n575) );
  NAND2_X1 U555 ( .A1(n328), .A2(n314), .ZN(n119) );
  OR2_X1 U556 ( .A1(n224), .A2(n227), .ZN(n558) );
  OR2_X1 U557 ( .A1(n233), .A2(n232), .ZN(n559) );
  OR2_X1 U558 ( .A1(n328), .A2(n314), .ZN(n560) );
  OR2_X1 U559 ( .A1(n151), .A2(n139), .ZN(n561) );
  NOR2_X1 U560 ( .A1(n218), .A2(n223), .ZN(n97) );
  NAND2_X1 U561 ( .A1(n218), .A2(n223), .ZN(n98) );
  NAND2_X1 U562 ( .A1(n228), .A2(n231), .ZN(n106) );
  INV_X1 U563 ( .A(n41), .ZN(n235) );
  AND2_X1 U564 ( .A1(n493), .A2(n122), .ZN(product[1]) );
  XNOR2_X1 U565 ( .A(n583), .B(a[14]), .ZN(n41) );
  OR2_X1 U566 ( .A1(n569), .A2(n495), .ZN(n392) );
  XNOR2_X1 U567 ( .A(n526), .B(n43), .ZN(n363) );
  AND2_X1 U568 ( .A1(n569), .A2(n548), .ZN(n300) );
  AND2_X1 U569 ( .A1(n569), .A2(n492), .ZN(n278) );
  AND2_X1 U570 ( .A1(n569), .A2(n540), .ZN(n270) );
  XNOR2_X1 U571 ( .A(n155), .B(n563), .ZN(n139) );
  XNOR2_X1 U572 ( .A(n153), .B(n141), .ZN(n563) );
  XNOR2_X1 U573 ( .A(n157), .B(n564), .ZN(n141) );
  XNOR2_X1 U574 ( .A(n145), .B(n143), .ZN(n564) );
  OAI22_X1 U575 ( .A1(n39), .A2(n584), .B1(n337), .B2(n37), .ZN(n252) );
  OR2_X1 U576 ( .A1(n569), .A2(n584), .ZN(n337) );
  OAI22_X1 U577 ( .A1(n42), .A2(n586), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U578 ( .A1(n43), .A2(n586), .ZN(n332) );
  XNOR2_X1 U579 ( .A(n159), .B(n565), .ZN(n142) );
  XNOR2_X1 U580 ( .A(n315), .B(n261), .ZN(n565) );
  XNOR2_X1 U581 ( .A(n576), .B(n43), .ZN(n376) );
  XNOR2_X1 U582 ( .A(n583), .B(n43), .ZN(n336) );
  AND2_X1 U583 ( .A1(n569), .A2(n247), .ZN(n314) );
  OAI22_X1 U584 ( .A1(n39), .A2(n336), .B1(n37), .B2(n335), .ZN(n263) );
  AND2_X1 U585 ( .A1(n569), .A2(n519), .ZN(n264) );
  AND2_X1 U586 ( .A1(n569), .A2(n555), .ZN(n288) );
  AND2_X1 U587 ( .A1(n569), .A2(n235), .ZN(n260) );
  OAI22_X1 U588 ( .A1(n39), .A2(n335), .B1(n37), .B2(n334), .ZN(n262) );
  NAND2_X1 U589 ( .A1(n427), .A2(n37), .ZN(n39) );
  XOR2_X1 U590 ( .A(n583), .B(a[12]), .Z(n427) );
  INV_X1 U591 ( .A(n25), .ZN(n580) );
  XNOR2_X1 U592 ( .A(n579), .B(n43), .ZN(n352) );
  NAND2_X1 U593 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U594 ( .A(n585), .B(a[14]), .Z(n426) );
  INV_X1 U595 ( .A(n7), .ZN(n574) );
  AND2_X1 U596 ( .A1(n569), .A2(n249), .ZN(product[0]) );
  OR2_X1 U597 ( .A1(n43), .A2(n582), .ZN(n344) );
  OR2_X1 U598 ( .A1(n43), .A2(n580), .ZN(n353) );
  OR2_X1 U599 ( .A1(n43), .A2(n578), .ZN(n364) );
  OR2_X1 U600 ( .A1(n569), .A2(n500), .ZN(n377) );
  XNOR2_X1 U601 ( .A(n526), .B(b[9]), .ZN(n354) );
  XNOR2_X1 U602 ( .A(n576), .B(b[11]), .ZN(n365) );
  OAI22_X1 U603 ( .A1(n39), .A2(n334), .B1(n37), .B2(n333), .ZN(n261) );
  XNOR2_X1 U604 ( .A(n583), .B(n422), .ZN(n333) );
  XNOR2_X1 U605 ( .A(n583), .B(n424), .ZN(n335) );
  XNOR2_X1 U606 ( .A(n583), .B(n423), .ZN(n334) );
  OAI22_X1 U607 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U608 ( .A(n585), .B(n424), .ZN(n330) );
  XNOR2_X1 U609 ( .A(n585), .B(n43), .ZN(n331) );
  XNOR2_X1 U610 ( .A(n573), .B(b[13]), .ZN(n378) );
  XNOR2_X1 U611 ( .A(n579), .B(n418), .ZN(n345) );
  XNOR2_X1 U612 ( .A(n581), .B(n420), .ZN(n338) );
  XNOR2_X1 U613 ( .A(n572), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U614 ( .A(n572), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U615 ( .A(n573), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U616 ( .A(n572), .B(n418), .ZN(n384) );
  XNOR2_X1 U617 ( .A(n572), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U618 ( .A(n573), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U619 ( .A(n573), .B(n419), .ZN(n385) );
  XNOR2_X1 U620 ( .A(n526), .B(n424), .ZN(n362) );
  XNOR2_X1 U621 ( .A(n579), .B(n424), .ZN(n351) );
  XNOR2_X1 U622 ( .A(n576), .B(n418), .ZN(n369) );
  XNOR2_X1 U623 ( .A(n576), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U624 ( .A(n576), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U625 ( .A(n576), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U626 ( .A(n526), .B(n423), .ZN(n361) );
  XNOR2_X1 U627 ( .A(n579), .B(n423), .ZN(n350) );
  XNOR2_X1 U628 ( .A(n512), .B(b[11]), .ZN(n397) );
  XNOR2_X1 U629 ( .A(n511), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U630 ( .A(n512), .B(b[13]), .ZN(n395) );
  XNOR2_X1 U631 ( .A(n512), .B(b[14]), .ZN(n394) );
  XNOR2_X1 U632 ( .A(n579), .B(n422), .ZN(n349) );
  XNOR2_X1 U633 ( .A(n526), .B(n422), .ZN(n360) );
  XNOR2_X1 U634 ( .A(n526), .B(n421), .ZN(n359) );
  XNOR2_X1 U635 ( .A(n526), .B(n420), .ZN(n358) );
  XNOR2_X1 U636 ( .A(n579), .B(n421), .ZN(n348) );
  XNOR2_X1 U637 ( .A(n579), .B(n420), .ZN(n347) );
  XNOR2_X1 U638 ( .A(n581), .B(n421), .ZN(n339) );
  XNOR2_X1 U639 ( .A(n526), .B(n418), .ZN(n356) );
  XNOR2_X1 U640 ( .A(n526), .B(n419), .ZN(n357) );
  XNOR2_X1 U641 ( .A(n579), .B(n419), .ZN(n346) );
  XNOR2_X1 U642 ( .A(n526), .B(b[8]), .ZN(n355) );
  XNOR2_X1 U643 ( .A(n511), .B(b[15]), .ZN(n393) );
  BUF_X1 U644 ( .A(n43), .Z(n569) );
  XNOR2_X1 U645 ( .A(n581), .B(n422), .ZN(n340) );
  XNOR2_X1 U646 ( .A(n581), .B(n424), .ZN(n342) );
  XNOR2_X1 U647 ( .A(n581), .B(n423), .ZN(n341) );
  XNOR2_X1 U648 ( .A(n581), .B(n43), .ZN(n343) );
  XNOR2_X1 U649 ( .A(n575), .B(n419), .ZN(n370) );
  XNOR2_X1 U650 ( .A(n576), .B(n424), .ZN(n375) );
  XNOR2_X1 U651 ( .A(n575), .B(n420), .ZN(n371) );
  XNOR2_X1 U652 ( .A(n575), .B(n423), .ZN(n374) );
  XNOR2_X1 U653 ( .A(n575), .B(n422), .ZN(n373) );
  XNOR2_X1 U654 ( .A(n575), .B(n421), .ZN(n372) );
  INV_X1 U655 ( .A(n521), .ZN(n127) );
  NOR2_X1 U656 ( .A1(n521), .A2(n85), .ZN(n80) );
  OAI21_X1 U657 ( .B1(n82), .B2(n86), .A(n83), .ZN(n81) );
  OAI22_X1 U658 ( .A1(n34), .A2(n339), .B1(n338), .B2(n32), .ZN(n265) );
  OAI22_X1 U659 ( .A1(n34), .A2(n340), .B1(n339), .B2(n32), .ZN(n266) );
  OAI22_X1 U660 ( .A1(n34), .A2(n341), .B1(n340), .B2(n32), .ZN(n267) );
  OAI22_X1 U661 ( .A1(n34), .A2(n342), .B1(n341), .B2(n32), .ZN(n268) );
  OAI22_X1 U662 ( .A1(n34), .A2(n343), .B1(n342), .B2(n32), .ZN(n269) );
  OAI22_X1 U663 ( .A1(n34), .A2(n582), .B1(n344), .B2(n32), .ZN(n253) );
  NOR2_X1 U664 ( .A1(n234), .A2(n257), .ZN(n113) );
  OAI22_X1 U665 ( .A1(n539), .A2(n394), .B1(n393), .B2(n546), .ZN(n315) );
  OAI22_X1 U666 ( .A1(n539), .A2(n395), .B1(n394), .B2(n547), .ZN(n316) );
  OAI22_X1 U667 ( .A1(n539), .A2(n400), .B1(n399), .B2(n546), .ZN(n321) );
  OAI22_X1 U668 ( .A1(n539), .A2(n398), .B1(n397), .B2(n547), .ZN(n319) );
  OAI22_X1 U669 ( .A1(n539), .A2(n401), .B1(n400), .B2(n546), .ZN(n322) );
  OAI22_X1 U670 ( .A1(n539), .A2(n397), .B1(n396), .B2(n547), .ZN(n318) );
  OAI22_X1 U671 ( .A1(n539), .A2(n396), .B1(n395), .B2(n546), .ZN(n317) );
  OAI22_X1 U672 ( .A1(n539), .A2(n399), .B1(n398), .B2(n546), .ZN(n320) );
  OAI22_X1 U673 ( .A1(n6), .A2(n404), .B1(n403), .B2(n546), .ZN(n325) );
  OAI22_X1 U674 ( .A1(n539), .A2(n405), .B1(n404), .B2(n547), .ZN(n326) );
  OAI22_X1 U675 ( .A1(n539), .A2(n406), .B1(n405), .B2(n547), .ZN(n327) );
  OAI22_X1 U676 ( .A1(n539), .A2(n402), .B1(n401), .B2(n547), .ZN(n323) );
  OAI22_X1 U677 ( .A1(n539), .A2(n407), .B1(n406), .B2(n547), .ZN(n328) );
  OAI22_X1 U678 ( .A1(n539), .A2(n408), .B1(n407), .B2(n546), .ZN(n329) );
  NOR2_X1 U679 ( .A1(n228), .A2(n231), .ZN(n105) );
  OAI21_X1 U680 ( .B1(n87), .B2(n85), .A(n517), .ZN(n84) );
  XNOR2_X1 U681 ( .A(n63), .B(n46), .ZN(product[15]) );
  INV_X1 U682 ( .A(n19), .ZN(n578) );
  NAND2_X1 U683 ( .A1(n204), .A2(n211), .ZN(n90) );
  NOR2_X1 U684 ( .A1(n204), .A2(n211), .ZN(n89) );
  OAI22_X1 U685 ( .A1(n29), .A2(n350), .B1(n349), .B2(n494), .ZN(n275) );
  OAI22_X1 U686 ( .A1(n29), .A2(n346), .B1(n345), .B2(n494), .ZN(n271) );
  OAI22_X1 U687 ( .A1(n502), .A2(n348), .B1(n347), .B2(n524), .ZN(n273) );
  OAI22_X1 U688 ( .A1(n502), .A2(n347), .B1(n346), .B2(n524), .ZN(n272) );
  OAI22_X1 U689 ( .A1(n29), .A2(n351), .B1(n350), .B2(n507), .ZN(n276) );
  OAI22_X1 U690 ( .A1(n502), .A2(n349), .B1(n348), .B2(n494), .ZN(n274) );
  OAI22_X1 U691 ( .A1(n29), .A2(n580), .B1(n353), .B2(n494), .ZN(n254) );
  OAI22_X1 U692 ( .A1(n502), .A2(n352), .B1(n351), .B2(n524), .ZN(n277) );
  XNOR2_X1 U693 ( .A(n77), .B(n48), .ZN(product[13]) );
  INV_X1 U694 ( .A(n88), .ZN(n87) );
  XNOR2_X1 U695 ( .A(n70), .B(n47), .ZN(product[14]) );
  INV_X1 U696 ( .A(n13), .ZN(n577) );
  INV_X1 U697 ( .A(n512), .ZN(n568) );
  OAI21_X1 U698 ( .B1(n99), .B2(n97), .A(n98), .ZN(n96) );
  NOR2_X1 U699 ( .A1(n176), .A2(n185), .ZN(n78) );
  XNOR2_X1 U700 ( .A(n572), .B(n420), .ZN(n386) );
  XNOR2_X1 U701 ( .A(n572), .B(n43), .ZN(n391) );
  XNOR2_X1 U702 ( .A(n572), .B(n424), .ZN(n390) );
  XNOR2_X1 U703 ( .A(n572), .B(n422), .ZN(n388) );
  XNOR2_X1 U704 ( .A(n572), .B(n421), .ZN(n387) );
  XNOR2_X1 U705 ( .A(n572), .B(n423), .ZN(n389) );
  INV_X1 U706 ( .A(n1), .ZN(n571) );
  OR2_X1 U707 ( .A1(n43), .A2(n568), .ZN(n409) );
  NAND2_X1 U708 ( .A1(n224), .A2(n227), .ZN(n103) );
  AOI21_X1 U709 ( .B1(n559), .B2(n112), .A(n532), .ZN(n107) );
  OAI21_X1 U710 ( .B1(n64), .B2(n528), .A(n65), .ZN(n63) );
  OAI22_X1 U711 ( .A1(n506), .A2(n358), .B1(n357), .B2(n510), .ZN(n282) );
  OAI22_X1 U712 ( .A1(n506), .A2(n356), .B1(n355), .B2(n491), .ZN(n280) );
  OAI22_X1 U713 ( .A1(n506), .A2(n362), .B1(n361), .B2(n491), .ZN(n286) );
  OAI22_X1 U714 ( .A1(n496), .A2(n578), .B1(n364), .B2(n510), .ZN(n255) );
  OAI22_X1 U715 ( .A1(n496), .A2(n357), .B1(n356), .B2(n510), .ZN(n281) );
  OAI22_X1 U716 ( .A1(n497), .A2(n355), .B1(n354), .B2(n510), .ZN(n279) );
  OAI22_X1 U717 ( .A1(n497), .A2(n363), .B1(n362), .B2(n509), .ZN(n287) );
  OAI22_X1 U718 ( .A1(n497), .A2(n361), .B1(n360), .B2(n510), .ZN(n285) );
  OAI22_X1 U719 ( .A1(n496), .A2(n360), .B1(n359), .B2(n509), .ZN(n284) );
  OAI22_X1 U720 ( .A1(n23), .A2(n359), .B1(n358), .B2(n508), .ZN(n283) );
  XOR2_X1 U721 ( .A(n56), .B(n545), .Z(product[5]) );
  NAND2_X1 U722 ( .A1(n151), .A2(n139), .ZN(n62) );
  OAI22_X1 U723 ( .A1(n530), .A2(n370), .B1(n369), .B2(n16), .ZN(n293) );
  OAI22_X1 U724 ( .A1(n530), .A2(n367), .B1(n366), .B2(n16), .ZN(n290) );
  OAI22_X1 U725 ( .A1(n530), .A2(n375), .B1(n374), .B2(n16), .ZN(n298) );
  OAI22_X1 U726 ( .A1(n18), .A2(n374), .B1(n373), .B2(n16), .ZN(n297) );
  OAI22_X1 U727 ( .A1(n530), .A2(n368), .B1(n367), .B2(n16), .ZN(n291) );
  OAI22_X1 U728 ( .A1(n18), .A2(n372), .B1(n371), .B2(n16), .ZN(n295) );
  OAI22_X1 U729 ( .A1(n530), .A2(n373), .B1(n372), .B2(n16), .ZN(n296) );
  OAI22_X1 U730 ( .A1(n18), .A2(n369), .B1(n368), .B2(n16), .ZN(n292) );
  OAI22_X1 U731 ( .A1(n530), .A2(n371), .B1(n370), .B2(n16), .ZN(n294) );
  OAI22_X1 U732 ( .A1(n530), .A2(n376), .B1(n375), .B2(n16), .ZN(n299) );
  OAI22_X1 U733 ( .A1(n18), .A2(n500), .B1(n377), .B2(n16), .ZN(n256) );
  OAI22_X1 U734 ( .A1(n18), .A2(n366), .B1(n365), .B2(n16), .ZN(n289) );
  NAND2_X1 U735 ( .A1(n135), .A2(n114), .ZN(n58) );
  XNOR2_X1 U736 ( .A(n512), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U737 ( .A(n513), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U738 ( .A(n513), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U739 ( .A(n513), .B(n418), .ZN(n401) );
  XNOR2_X1 U740 ( .A(n513), .B(n419), .ZN(n402) );
  XNOR2_X1 U741 ( .A(n513), .B(n420), .ZN(n403) );
  XNOR2_X1 U742 ( .A(n513), .B(n421), .ZN(n404) );
  XNOR2_X1 U743 ( .A(n512), .B(n422), .ZN(n405) );
  XNOR2_X1 U744 ( .A(n512), .B(n43), .ZN(n408) );
  XNOR2_X1 U745 ( .A(n511), .B(n423), .ZN(n406) );
  XNOR2_X1 U746 ( .A(n511), .B(n424), .ZN(n407) );
  OAI21_X1 U747 ( .B1(n528), .B2(n71), .A(n72), .ZN(n70) );
  OAI21_X1 U748 ( .B1(n45), .B2(n78), .A(n79), .ZN(n77) );
  XNOR2_X1 U749 ( .A(n499), .B(n53), .ZN(product[8]) );
  INV_X1 U750 ( .A(n122), .ZN(n120) );
  NAND2_X1 U751 ( .A1(n329), .A2(n258), .ZN(n122) );
  AOI21_X1 U752 ( .B1(n104), .B2(n558), .A(n101), .ZN(n99) );
  OAI22_X1 U753 ( .A1(n6), .A2(n568), .B1(n409), .B2(n546), .ZN(n258) );
  XOR2_X1 U754 ( .A(n544), .B(n54), .Z(product[7]) );
  OAI22_X1 U755 ( .A1(n515), .A2(n379), .B1(n378), .B2(n567), .ZN(n301) );
  OAI22_X1 U756 ( .A1(n12), .A2(n380), .B1(n379), .B2(n567), .ZN(n302) );
  OAI22_X1 U757 ( .A1(n543), .A2(n385), .B1(n384), .B2(n567), .ZN(n307) );
  OAI22_X1 U758 ( .A1(n12), .A2(n382), .B1(n381), .B2(n567), .ZN(n304) );
  OAI22_X1 U759 ( .A1(n542), .A2(n381), .B1(n380), .B2(n567), .ZN(n303) );
  NAND2_X1 U760 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U761 ( .A1(n542), .A2(n383), .B1(n567), .B2(n382), .ZN(n305) );
  OAI22_X1 U762 ( .A1(n543), .A2(n384), .B1(n383), .B2(n567), .ZN(n306) );
  OAI22_X1 U763 ( .A1(n543), .A2(n386), .B1(n385), .B2(n567), .ZN(n308) );
  OAI22_X1 U764 ( .A1(n542), .A2(n387), .B1(n386), .B2(n567), .ZN(n309) );
  OAI22_X1 U765 ( .A1(n542), .A2(n495), .B1(n392), .B2(n567), .ZN(n257) );
  OAI22_X1 U766 ( .A1(n12), .A2(n389), .B1(n567), .B2(n388), .ZN(n311) );
  OAI22_X1 U767 ( .A1(n543), .A2(n388), .B1(n387), .B2(n567), .ZN(n310) );
  OAI22_X1 U768 ( .A1(n515), .A2(n390), .B1(n389), .B2(n567), .ZN(n312) );
  INV_X1 U769 ( .A(n567), .ZN(n247) );
  OAI22_X1 U770 ( .A1(n515), .A2(n391), .B1(n390), .B2(n567), .ZN(n313) );
  INV_X1 U771 ( .A(n574), .ZN(n573) );
  INV_X1 U772 ( .A(n31), .ZN(n582) );
  INV_X1 U773 ( .A(n36), .ZN(n584) );
  INV_X1 U774 ( .A(n586), .ZN(n585) );
  INV_X1 U775 ( .A(n40), .ZN(n586) );
  XOR2_X1 U776 ( .A(n259), .B(n251), .Z(n148) );
  XOR2_X1 U777 ( .A(n289), .B(n279), .Z(n146) );
  XOR2_X1 U778 ( .A(n149), .B(n147), .Z(n144) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_2_DW01_add_2 ( A, B, CI, SUM, 
        CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n4, n7, n8, n9, n10, n11, n12, n13, n14, n15, n18, n19, n20,
         n21, n23, n25, n26, n27, n28, n30, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n48, n49, n51, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n71, n72, n73, n74,
         n75, n77, n79, n80, n81, n82, n83, n85, n87, n88, n90, n93, n94, n99,
         n100, n102, n104, n161, n162, n163, n164, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184;

  AOI21_X1 U126 ( .B1(n56), .B2(n64), .A(n57), .ZN(n161) );
  OR2_X1 U127 ( .A1(A[11]), .A2(B[11]), .ZN(n162) );
  OR2_X1 U128 ( .A1(A[10]), .A2(B[10]), .ZN(n163) );
  OR2_X1 U129 ( .A1(A[10]), .A2(B[10]), .ZN(n183) );
  OR2_X1 U130 ( .A1(A[8]), .A2(B[8]), .ZN(n164) );
  AND2_X1 U131 ( .A1(n178), .A2(n90), .ZN(SUM[0]) );
  OR2_X1 U132 ( .A1(A[15]), .A2(B[15]), .ZN(n166) );
  XNOR2_X1 U133 ( .A(n49), .B(n167), .ZN(SUM[10]) );
  AND2_X1 U134 ( .A1(n163), .A2(n48), .ZN(n167) );
  XNOR2_X1 U135 ( .A(n41), .B(n168), .ZN(SUM[11]) );
  AND2_X1 U136 ( .A1(n162), .A2(n40), .ZN(n168) );
  XNOR2_X1 U137 ( .A(n33), .B(n169), .ZN(SUM[13]) );
  AND2_X1 U138 ( .A1(n93), .A2(n28), .ZN(n169) );
  BUF_X1 U139 ( .A(n34), .Z(n172) );
  INV_X1 U140 ( .A(n162), .ZN(n170) );
  NOR2_X1 U141 ( .A1(A[8]), .A2(B[8]), .ZN(n171) );
  BUF_X1 U142 ( .A(n35), .Z(n173) );
  NOR2_X1 U143 ( .A1(A[12]), .A2(B[12]), .ZN(n174) );
  NOR2_X1 U144 ( .A1(A[12]), .A2(B[12]), .ZN(n36) );
  CLKBUF_X1 U145 ( .A(n42), .Z(n175) );
  INV_X1 U146 ( .A(n176), .ZN(n48) );
  AND2_X1 U147 ( .A1(A[10]), .A2(B[10]), .ZN(n176) );
  AOI21_X1 U148 ( .B1(n42), .B2(n34), .A(n35), .ZN(n177) );
  OR2_X1 U149 ( .A1(A[0]), .A2(B[0]), .ZN(n178) );
  INV_X1 U150 ( .A(n161), .ZN(n54) );
  INV_X1 U151 ( .A(n42), .ZN(n41) );
  AOI21_X1 U152 ( .B1(n175), .B2(n172), .A(n173), .ZN(n33) );
  AOI21_X1 U153 ( .B1(n181), .B2(n80), .A(n77), .ZN(n75) );
  INV_X1 U154 ( .A(n79), .ZN(n77) );
  AOI21_X1 U155 ( .B1(n182), .B2(n88), .A(n85), .ZN(n83) );
  INV_X1 U156 ( .A(n87), .ZN(n85) );
  AOI21_X1 U157 ( .B1(n56), .B2(n64), .A(n57), .ZN(n55) );
  OAI21_X1 U158 ( .B1(n83), .B2(n81), .A(n82), .ZN(n80) );
  AOI21_X1 U159 ( .B1(n184), .B2(n72), .A(n69), .ZN(n67) );
  INV_X1 U160 ( .A(n71), .ZN(n69) );
  NAND2_X1 U161 ( .A1(n179), .A2(n93), .ZN(n20) );
  AOI21_X1 U162 ( .B1(n179), .B2(n30), .A(n23), .ZN(n21) );
  OAI21_X1 U163 ( .B1(n75), .B2(n73), .A(n74), .ZN(n72) );
  AOI21_X1 U164 ( .B1(n54), .B2(n180), .A(n51), .ZN(n49) );
  NAND2_X1 U165 ( .A1(n164), .A2(n59), .ZN(n8) );
  INV_X1 U166 ( .A(n90), .ZN(n88) );
  OAI21_X1 U167 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  INV_X1 U168 ( .A(n53), .ZN(n51) );
  INV_X1 U169 ( .A(n27), .ZN(n93) );
  INV_X1 U170 ( .A(n25), .ZN(n23) );
  NAND2_X1 U171 ( .A1(n102), .A2(n74), .ZN(n12) );
  INV_X1 U172 ( .A(n73), .ZN(n102) );
  INV_X1 U173 ( .A(n174), .ZN(n94) );
  NAND2_X1 U174 ( .A1(n180), .A2(n53), .ZN(n7) );
  NAND2_X1 U175 ( .A1(n99), .A2(n62), .ZN(n9) );
  INV_X1 U176 ( .A(n61), .ZN(n99) );
  NAND2_X1 U177 ( .A1(n104), .A2(n82), .ZN(n14) );
  INV_X1 U178 ( .A(n81), .ZN(n104) );
  NAND2_X1 U179 ( .A1(n184), .A2(n71), .ZN(n11) );
  NAND2_X1 U180 ( .A1(n181), .A2(n79), .ZN(n13) );
  NAND2_X1 U181 ( .A1(n182), .A2(n87), .ZN(n15) );
  NAND2_X1 U182 ( .A1(n100), .A2(n66), .ZN(n10) );
  INV_X1 U183 ( .A(n65), .ZN(n100) );
  XNOR2_X1 U184 ( .A(n11), .B(n72), .ZN(SUM[5]) );
  XOR2_X1 U185 ( .A(n12), .B(n75), .Z(SUM[4]) );
  XNOR2_X1 U186 ( .A(n13), .B(n80), .ZN(SUM[3]) );
  XNOR2_X1 U187 ( .A(n15), .B(n88), .ZN(SUM[1]) );
  NAND2_X1 U188 ( .A1(n94), .A2(n37), .ZN(n4) );
  OR2_X1 U189 ( .A1(A[14]), .A2(B[14]), .ZN(n179) );
  NOR2_X1 U190 ( .A1(A[7]), .A2(B[7]), .ZN(n61) );
  OR2_X1 U191 ( .A1(A[9]), .A2(B[9]), .ZN(n180) );
  NOR2_X1 U192 ( .A1(A[2]), .A2(B[2]), .ZN(n81) );
  NOR2_X1 U193 ( .A1(A[4]), .A2(B[4]), .ZN(n73) );
  NAND2_X1 U194 ( .A1(n179), .A2(n25), .ZN(n2) );
  OR2_X1 U195 ( .A1(A[3]), .A2(B[3]), .ZN(n181) );
  OR2_X1 U196 ( .A1(A[1]), .A2(B[1]), .ZN(n182) );
  NOR2_X1 U197 ( .A1(A[8]), .A2(B[8]), .ZN(n58) );
  XNOR2_X1 U198 ( .A(n60), .B(n8), .ZN(SUM[8]) );
  NOR2_X1 U199 ( .A1(A[6]), .A2(B[6]), .ZN(n65) );
  NAND2_X1 U200 ( .A1(A[7]), .A2(B[7]), .ZN(n62) );
  OR2_X1 U201 ( .A1(A[5]), .A2(B[5]), .ZN(n184) );
  NAND2_X1 U202 ( .A1(A[2]), .A2(B[2]), .ZN(n82) );
  NAND2_X1 U203 ( .A1(A[4]), .A2(B[4]), .ZN(n74) );
  NAND2_X1 U204 ( .A1(A[3]), .A2(B[3]), .ZN(n79) );
  NAND2_X1 U205 ( .A1(A[1]), .A2(B[1]), .ZN(n87) );
  NAND2_X1 U206 ( .A1(A[5]), .A2(B[5]), .ZN(n71) );
  NAND2_X1 U207 ( .A1(A[0]), .A2(B[0]), .ZN(n90) );
  NAND2_X1 U208 ( .A1(A[11]), .A2(B[11]), .ZN(n40) );
  NAND2_X1 U209 ( .A1(A[8]), .A2(B[8]), .ZN(n59) );
  NAND2_X1 U210 ( .A1(A[6]), .A2(B[6]), .ZN(n66) );
  XNOR2_X1 U211 ( .A(n54), .B(n7), .ZN(SUM[9]) );
  XOR2_X1 U212 ( .A(n63), .B(n9), .Z(SUM[7]) );
  XOR2_X1 U213 ( .A(n14), .B(n83), .Z(SUM[2]) );
  NAND2_X1 U214 ( .A1(n166), .A2(n18), .ZN(n1) );
  NAND2_X1 U215 ( .A1(A[15]), .A2(B[15]), .ZN(n18) );
  NOR2_X1 U216 ( .A1(n171), .A2(n61), .ZN(n56) );
  OAI21_X1 U217 ( .B1(n58), .B2(n62), .A(n59), .ZN(n57) );
  NAND2_X1 U218 ( .A1(A[12]), .A2(B[12]), .ZN(n37) );
  INV_X1 U219 ( .A(n28), .ZN(n30) );
  INV_X1 U220 ( .A(n64), .ZN(n63) );
  NAND2_X1 U221 ( .A1(A[9]), .A2(B[9]), .ZN(n53) );
  NAND2_X1 U222 ( .A1(A[14]), .A2(B[14]), .ZN(n25) );
  NAND2_X1 U223 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  NOR2_X1 U224 ( .A1(A[13]), .A2(B[13]), .ZN(n27) );
  XOR2_X1 U225 ( .A(n67), .B(n10), .Z(SUM[6]) );
  OAI21_X1 U226 ( .B1(n67), .B2(n65), .A(n66), .ZN(n64) );
  OAI21_X1 U227 ( .B1(n36), .B2(n40), .A(n37), .ZN(n35) );
  AOI21_X1 U228 ( .B1(n183), .B2(n51), .A(n176), .ZN(n44) );
  OAI21_X1 U229 ( .B1(n41), .B2(n170), .A(n40), .ZN(n38) );
  NOR2_X1 U230 ( .A1(n174), .A2(n39), .ZN(n34) );
  NOR2_X1 U231 ( .A1(A[11]), .A2(B[11]), .ZN(n39) );
  OAI21_X1 U232 ( .B1(n43), .B2(n55), .A(n44), .ZN(n42) );
  NAND2_X1 U233 ( .A1(n163), .A2(n180), .ZN(n43) );
  XNOR2_X1 U234 ( .A(n38), .B(n4), .ZN(SUM[12]) );
  XNOR2_X1 U235 ( .A(n19), .B(n1), .ZN(SUM[15]) );
  XNOR2_X1 U236 ( .A(n26), .B(n2), .ZN(SUM[14]) );
  OAI21_X1 U237 ( .B1(n177), .B2(n27), .A(n28), .ZN(n26) );
  OAI21_X1 U238 ( .B1(n177), .B2(n20), .A(n21), .ZN(n19) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_2 ( clk, clear_acc, 
        data_out_x, data_out, data_out_w, data_out_b, wr_en_y, m_valid, 
        m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [3:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N27, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, n1, n2, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n87, n104, n113, n114, n115, n116, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n22), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n227), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n228), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n229), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n230), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n231), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n232), .CK(clk), .Q(n34) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n233), .CK(clk), .Q(n35) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n234), .CK(clk), .Q(n36) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n235), .CK(clk), .Q(n37) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n236), .CK(clk), .Q(n38) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n237), .CK(clk), .Q(n39) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n238), .CK(clk), .Q(n40) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n239), .CK(clk), .Q(n41) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n240), .CK(clk), .Q(n42) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n241), .CK(clk), .Q(n43) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n242), .CK(clk), .Q(n45) );
  DFF_X1 \f_reg[7]  ( .D(n84), .CK(clk), .Q(f[7]), .QN(n219) );
  DFF_X1 \f_reg[8]  ( .D(n83), .CK(clk), .Q(f[8]), .QN(n220) );
  DFF_X1 \f_reg[9]  ( .D(n82), .CK(clk), .Q(f[9]), .QN(n221) );
  DFF_X1 \f_reg[10]  ( .D(n81), .CK(clk), .Q(n54), .QN(n222) );
  DFF_X1 \f_reg[11]  ( .D(n80), .CK(clk), .Q(n52), .QN(n223) );
  DFF_X1 \f_reg[12]  ( .D(n2), .CK(clk), .Q(n51), .QN(n224) );
  DFF_X1 \f_reg[13]  ( .D(n7), .CK(clk), .Q(n50), .QN(n225) );
  DFF_X1 \f_reg[14]  ( .D(n1), .CK(clk), .Q(n49), .QN(n226) );
  DFF_X1 \f_reg[15]  ( .D(n11), .CK(clk), .Q(f[15]), .QN(n78) );
  DFF_X1 \data_out_reg[15]  ( .D(n168), .CK(clk), .Q(data_out[15]), .QN(n199)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n169), .CK(clk), .Q(data_out[14]), .QN(n198)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n170), .CK(clk), .Q(data_out[13]), .QN(n197)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n171), .CK(clk), .Q(data_out[12]), .QN(n196)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n172), .CK(clk), .Q(data_out[11]), .QN(n195)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n173), .CK(clk), .Q(data_out[10]), .QN(n194)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n174), .CK(clk), .Q(data_out[9]), .QN(n193) );
  DFF_X1 \data_out_reg[8]  ( .D(n175), .CK(clk), .Q(data_out[8]), .QN(n192) );
  DFF_X1 \data_out_reg[7]  ( .D(n176), .CK(clk), .Q(data_out[7]), .QN(n191) );
  DFF_X1 \data_out_reg[6]  ( .D(n177), .CK(clk), .Q(data_out[6]), .QN(n190) );
  DFF_X1 \data_out_reg[5]  ( .D(n178), .CK(clk), .Q(data_out[5]), .QN(n189) );
  DFF_X1 \data_out_reg[4]  ( .D(n179), .CK(clk), .Q(data_out[4]), .QN(n188) );
  DFF_X1 \data_out_reg[3]  ( .D(n180), .CK(clk), .Q(data_out[3]), .QN(n187) );
  DFF_X1 \data_out_reg[2]  ( .D(n181), .CK(clk), .Q(data_out[2]), .QN(n186) );
  DFF_X1 \data_out_reg[1]  ( .D(n182), .CK(clk), .Q(data_out[1]), .QN(n185) );
  DFF_X1 \data_out_reg[0]  ( .D(n183), .CK(clk), .Q(data_out[0]), .QN(n184) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_2_DW_mult_tc_1 mult_960 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_2_DW01_add_2 add_961 ( .A({n206, 
        n205, n204, n203, n202, n201, n215, n214, n213, n212, n211, n210, n209, 
        n208, n207, n200}), .B({f[15], n49, n50, n51, n52, n54, f[9:3], n62, 
        n64, n66}), .CI(1'b0), .SUM(adder) );
  DFF_X2 delay_reg ( .D(N27), .CK(clk), .Q(n19), .QN(n243) );
  DFF_X1 \f_reg[2]  ( .D(n114), .CK(clk), .Q(n62), .QN(n218) );
  DFF_X1 \f_reg[3]  ( .D(n113), .CK(clk), .Q(f[3]), .QN(n70) );
  DFF_X1 \f_reg[1]  ( .D(n115), .CK(clk), .Q(n64), .QN(n217) );
  DFF_X1 \f_reg[0]  ( .D(n116), .CK(clk), .Q(n66), .QN(n216) );
  DFF_X1 \f_reg[4]  ( .D(n104), .CK(clk), .Q(f[4]), .QN(n71) );
  DFF_X1 \f_reg[5]  ( .D(n87), .CK(clk), .Q(f[5]), .QN(n72) );
  DFF_X1 \f_reg[6]  ( .D(n85), .CK(clk), .Q(f[6]), .QN(n73) );
  MUX2_X2 U3 ( .A(n33), .B(N40), .S(n243), .Z(n202) );
  AND2_X2 U4 ( .A1(n48), .A2(n23), .ZN(n20) );
  NAND3_X1 U5 ( .A1(n17), .A2(n16), .A3(n18), .ZN(n1) );
  NAND3_X1 U6 ( .A1(n5), .A2(n4), .A3(n6), .ZN(n2) );
  MUX2_X2 U8 ( .A(n36), .B(N37), .S(n243), .Z(n214) );
  NAND2_X1 U9 ( .A1(data_out_b[12]), .A2(n22), .ZN(n4) );
  NAND2_X1 U10 ( .A1(adder[12]), .A2(n20), .ZN(n5) );
  NAND2_X1 U11 ( .A1(n68), .A2(n51), .ZN(n6) );
  NAND3_X1 U12 ( .A1(n9), .A2(n8), .A3(n10), .ZN(n7) );
  NAND2_X1 U13 ( .A1(data_out_b[13]), .A2(n22), .ZN(n8) );
  NAND2_X1 U14 ( .A1(adder[13]), .A2(n20), .ZN(n9) );
  NAND2_X1 U15 ( .A1(n68), .A2(n50), .ZN(n10) );
  NAND3_X1 U16 ( .A1(n13), .A2(n12), .A3(n14), .ZN(n11) );
  MUX2_X2 U17 ( .A(N42), .B(n29), .S(n19), .Z(n204) );
  MUX2_X2 U18 ( .A(N43), .B(n28), .S(n19), .Z(n205) );
  MUX2_X1 U19 ( .A(N39), .B(n34), .S(n19), .Z(n201) );
  NAND2_X1 U20 ( .A1(data_out_b[15]), .A2(n22), .ZN(n12) );
  NAND2_X1 U21 ( .A1(adder[15]), .A2(n20), .ZN(n13) );
  NAND2_X1 U22 ( .A1(n68), .A2(f[15]), .ZN(n14) );
  CLKBUF_X1 U23 ( .A(N39), .Z(n15) );
  NAND2_X1 U24 ( .A1(data_out_b[14]), .A2(n22), .ZN(n16) );
  NAND2_X1 U25 ( .A1(adder[14]), .A2(n20), .ZN(n17) );
  NAND2_X1 U26 ( .A1(n68), .A2(n49), .ZN(n18) );
  INV_X2 U27 ( .A(n48), .ZN(n68) );
  MUX2_X2 U28 ( .A(n32), .B(N41), .S(n243), .Z(n203) );
  INV_X1 U29 ( .A(n23), .ZN(n22) );
  INV_X1 U30 ( .A(clear_acc), .ZN(n23) );
  NAND2_X1 U31 ( .A1(n21), .A2(N27), .ZN(n245) );
  OAI22_X1 U32 ( .A1(n187), .A2(n245), .B1(n70), .B2(n244), .ZN(n180) );
  OAI22_X1 U33 ( .A1(n188), .A2(n245), .B1(n71), .B2(n244), .ZN(n179) );
  OAI22_X1 U34 ( .A1(n189), .A2(n245), .B1(n72), .B2(n244), .ZN(n178) );
  OAI22_X1 U35 ( .A1(n190), .A2(n245), .B1(n73), .B2(n244), .ZN(n177) );
  OAI22_X1 U36 ( .A1(n191), .A2(n245), .B1(n219), .B2(n244), .ZN(n176) );
  OAI22_X1 U37 ( .A1(n192), .A2(n245), .B1(n220), .B2(n244), .ZN(n175) );
  OAI22_X1 U38 ( .A1(n193), .A2(n245), .B1(n221), .B2(n244), .ZN(n174) );
  INV_X1 U39 ( .A(n26), .ZN(n44) );
  INV_X1 U40 ( .A(wr_en_y), .ZN(n21) );
  AND2_X1 U41 ( .A1(sel[0]), .A2(sel[1]), .ZN(n25) );
  INV_X1 U42 ( .A(m_ready), .ZN(n24) );
  NAND2_X1 U43 ( .A1(m_valid), .A2(n24), .ZN(n46) );
  OAI211_X1 U44 ( .C1(sel[2]), .C2(n25), .A(sel[3]), .B(n46), .ZN(N27) );
  NAND2_X1 U45 ( .A1(clear_acc_delay), .A2(n243), .ZN(n26) );
  MUX2_X1 U46 ( .A(n27), .B(N44), .S(n44), .Z(n227) );
  MUX2_X1 U47 ( .A(n27), .B(N44), .S(n243), .Z(n206) );
  MUX2_X1 U48 ( .A(n28), .B(N43), .S(n44), .Z(n228) );
  MUX2_X1 U49 ( .A(n29), .B(N42), .S(n44), .Z(n229) );
  MUX2_X1 U50 ( .A(n32), .B(N41), .S(n44), .Z(n230) );
  MUX2_X1 U51 ( .A(n33), .B(N40), .S(n44), .Z(n231) );
  MUX2_X1 U52 ( .A(n34), .B(n15), .S(n44), .Z(n232) );
  MUX2_X1 U53 ( .A(n35), .B(N38), .S(n44), .Z(n233) );
  MUX2_X1 U54 ( .A(n35), .B(N38), .S(n243), .Z(n215) );
  MUX2_X1 U55 ( .A(n36), .B(N37), .S(n44), .Z(n234) );
  MUX2_X1 U56 ( .A(n37), .B(N36), .S(n44), .Z(n235) );
  MUX2_X1 U57 ( .A(n37), .B(N36), .S(n243), .Z(n213) );
  MUX2_X1 U58 ( .A(n38), .B(N35), .S(n44), .Z(n236) );
  MUX2_X1 U59 ( .A(n38), .B(N35), .S(n243), .Z(n212) );
  MUX2_X1 U60 ( .A(n39), .B(N34), .S(n44), .Z(n237) );
  MUX2_X1 U61 ( .A(n39), .B(N34), .S(n243), .Z(n211) );
  MUX2_X1 U62 ( .A(n40), .B(N33), .S(n44), .Z(n238) );
  MUX2_X1 U63 ( .A(n40), .B(N33), .S(n243), .Z(n210) );
  MUX2_X1 U64 ( .A(n41), .B(N32), .S(n44), .Z(n239) );
  MUX2_X1 U65 ( .A(n41), .B(N32), .S(n243), .Z(n209) );
  MUX2_X1 U66 ( .A(n42), .B(N31), .S(n44), .Z(n240) );
  MUX2_X1 U67 ( .A(n42), .B(N31), .S(n243), .Z(n208) );
  MUX2_X1 U68 ( .A(n43), .B(N30), .S(n44), .Z(n241) );
  MUX2_X1 U69 ( .A(n43), .B(N30), .S(n243), .Z(n207) );
  MUX2_X1 U70 ( .A(n45), .B(N29), .S(n44), .Z(n242) );
  MUX2_X1 U71 ( .A(n45), .B(N29), .S(n243), .Z(n200) );
  INV_X1 U72 ( .A(n46), .ZN(n47) );
  OAI21_X1 U73 ( .B1(n47), .B2(n19), .A(n23), .ZN(n48) );
  AOI222_X1 U74 ( .A1(data_out_b[11]), .A2(n22), .B1(adder[11]), .B2(n20), 
        .C1(n68), .C2(n52), .ZN(n53) );
  INV_X1 U75 ( .A(n53), .ZN(n80) );
  AOI222_X1 U76 ( .A1(data_out_b[10]), .A2(n22), .B1(adder[10]), .B2(n20), 
        .C1(n68), .C2(n54), .ZN(n55) );
  INV_X1 U77 ( .A(n55), .ZN(n81) );
  AOI222_X1 U78 ( .A1(data_out_b[8]), .A2(n22), .B1(adder[8]), .B2(n20), .C1(
        n68), .C2(f[8]), .ZN(n56) );
  INV_X1 U79 ( .A(n56), .ZN(n83) );
  AOI222_X1 U80 ( .A1(data_out_b[7]), .A2(n22), .B1(adder[7]), .B2(n20), .C1(
        n68), .C2(f[7]), .ZN(n57) );
  INV_X1 U81 ( .A(n57), .ZN(n84) );
  AOI222_X1 U82 ( .A1(data_out_b[6]), .A2(n22), .B1(adder[6]), .B2(n20), .C1(
        n68), .C2(f[6]), .ZN(n58) );
  INV_X1 U83 ( .A(n58), .ZN(n85) );
  AOI222_X1 U84 ( .A1(data_out_b[5]), .A2(n22), .B1(adder[5]), .B2(n20), .C1(
        n68), .C2(f[5]), .ZN(n59) );
  INV_X1 U85 ( .A(n59), .ZN(n87) );
  AOI222_X1 U86 ( .A1(data_out_b[4]), .A2(n22), .B1(adder[4]), .B2(n20), .C1(
        n68), .C2(f[4]), .ZN(n60) );
  INV_X1 U87 ( .A(n60), .ZN(n104) );
  AOI222_X1 U88 ( .A1(data_out_b[3]), .A2(n22), .B1(adder[3]), .B2(n20), .C1(
        n68), .C2(f[3]), .ZN(n61) );
  INV_X1 U89 ( .A(n61), .ZN(n113) );
  AOI222_X1 U90 ( .A1(data_out_b[2]), .A2(n22), .B1(adder[2]), .B2(n20), .C1(
        n68), .C2(n62), .ZN(n63) );
  INV_X1 U91 ( .A(n63), .ZN(n114) );
  AOI222_X1 U92 ( .A1(data_out_b[1]), .A2(n22), .B1(adder[1]), .B2(n20), .C1(
        n68), .C2(n64), .ZN(n65) );
  INV_X1 U93 ( .A(n65), .ZN(n115) );
  AOI222_X1 U94 ( .A1(data_out_b[0]), .A2(n22), .B1(adder[0]), .B2(n20), .C1(
        n68), .C2(n66), .ZN(n67) );
  INV_X1 U95 ( .A(n67), .ZN(n116) );
  AOI222_X1 U96 ( .A1(data_out_b[9]), .A2(n22), .B1(adder[9]), .B2(n20), .C1(
        n68), .C2(f[9]), .ZN(n69) );
  INV_X1 U97 ( .A(n69), .ZN(n82) );
  NOR4_X1 U98 ( .A1(n52), .A2(n51), .A3(n50), .A4(n49), .ZN(n77) );
  NOR4_X1 U99 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n54), .ZN(n76) );
  NAND4_X1 U100 ( .A1(n73), .A2(n72), .A3(n71), .A4(n70), .ZN(n74) );
  NOR4_X1 U101 ( .A1(n74), .A2(n66), .A3(n64), .A4(n62), .ZN(n75) );
  NAND3_X1 U102 ( .A1(n77), .A2(n76), .A3(n75), .ZN(n79) );
  NAND3_X1 U103 ( .A1(wr_en_y), .A2(n79), .A3(n78), .ZN(n244) );
  OAI22_X1 U104 ( .A1(n184), .A2(n245), .B1(n216), .B2(n244), .ZN(n183) );
  OAI22_X1 U105 ( .A1(n185), .A2(n245), .B1(n217), .B2(n244), .ZN(n182) );
  OAI22_X1 U106 ( .A1(n186), .A2(n245), .B1(n218), .B2(n244), .ZN(n181) );
  OAI22_X1 U107 ( .A1(n194), .A2(n245), .B1(n222), .B2(n244), .ZN(n173) );
  OAI22_X1 U108 ( .A1(n195), .A2(n245), .B1(n223), .B2(n244), .ZN(n172) );
  OAI22_X1 U109 ( .A1(n196), .A2(n245), .B1(n224), .B2(n244), .ZN(n171) );
  OAI22_X1 U110 ( .A1(n197), .A2(n245), .B1(n225), .B2(n244), .ZN(n170) );
  OAI22_X1 U111 ( .A1(n198), .A2(n245), .B1(n226), .B2(n244), .ZN(n169) );
  OAI22_X1 U112 ( .A1(n199), .A2(n245), .B1(n78), .B2(n244), .ZN(n168) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_1_DW_mult_tc_1 ( a, b, 
        product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n9, n12, n13, n16, n18, n19, n21, n23, n25, n27, n29, n31,
         n32, n34, n36, n37, n39, n40, n41, n42, n43, n46, n47, n48, n49, n50,
         n52, n53, n54, n55, n56, n57, n58, n59, n62, n63, n64, n65, n67, n69,
         n70, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n93, n95, n96, n97, n98, n99, n103,
         n104, n105, n106, n107, n109, n111, n112, n113, n114, n115, n117,
         n119, n120, n122, n125, n126, n131, n135, n139, n141, n142, n143,
         n144, n145, n147, n148, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n237, n247, n249, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n418, n419,
         n420, n421, n422, n423, n424, n426, n427, n429, n431, n433, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U148 ( .A(n265), .B(n144), .Z(n145) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U161 ( .A(n177), .B(n168), .CI(n166), .CO(n163), .S(n164) );
  FA_X1 U162 ( .A(n170), .B(n172), .CI(n179), .CO(n165), .S(n166) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n273), .CI(n281), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n291), .CI(n263), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n317), .B(n252), .CO(n173), .S(n174) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U170 ( .A(n268), .B(n292), .CI(n274), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U173 ( .A(n199), .B(n201), .CI(n192), .CO(n187), .S(n188) );
  FA_X1 U174 ( .A(n275), .B(n293), .CI(n194), .CO(n189), .S(n190) );
  HA_X1 U176 ( .A(n269), .B(n319), .CO(n193), .S(n194) );
  FA_X1 U177 ( .A(n205), .B(n200), .CI(n198), .CO(n195), .S(n196) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U179 ( .A(n276), .B(n294), .CI(n284), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n320), .B(n270), .CI(n306), .CO(n201), .S(n202) );
  FA_X1 U181 ( .A(n208), .B(n213), .CI(n206), .CO(n203), .S(n204) );
  FA_X1 U182 ( .A(n210), .B(n307), .CI(n215), .CO(n205), .S(n206) );
  FA_X1 U183 ( .A(n254), .B(n285), .CI(n295), .CO(n207), .S(n208) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U185 ( .A(n216), .B(n219), .CI(n214), .CO(n211), .S(n212) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n322), .B(n278), .CI(n308), .CO(n215), .S(n216) );
  FA_X1 U189 ( .A(n255), .B(n309), .CI(n297), .CO(n219), .S(n220) );
  HA_X1 U190 ( .A(n323), .B(n287), .CO(n221), .S(n222) );
  FA_X1 U192 ( .A(n310), .B(n288), .CI(n324), .CO(n225), .S(n226) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  HA_X1 U194 ( .A(n311), .B(n325), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n326), .B(n300), .CI(n312), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  BUF_X1 U414 ( .A(n9), .Z(n589) );
  CLKBUF_X3 U415 ( .A(n9), .Z(n588) );
  OR2_X1 U416 ( .A1(n329), .A2(n258), .ZN(n490) );
  XNOR2_X1 U417 ( .A(n491), .B(n305), .ZN(n192) );
  XNOR2_X1 U418 ( .A(n253), .B(n283), .ZN(n491) );
  CLKBUF_X1 U419 ( .A(n86), .Z(n492) );
  INV_X1 U420 ( .A(n1), .ZN(n598) );
  XNOR2_X1 U421 ( .A(n88), .B(n493), .ZN(product[10]) );
  NAND2_X1 U422 ( .A1(n521), .A2(n86), .ZN(n493) );
  AOI21_X1 U423 ( .B1(n96), .B2(n579), .A(n93), .ZN(n494) );
  AOI21_X1 U424 ( .B1(n96), .B2(n579), .A(n93), .ZN(n91) );
  AOI21_X1 U425 ( .B1(n583), .B2(n112), .A(n109), .ZN(n495) );
  INV_X1 U426 ( .A(n600), .ZN(n496) );
  XNOR2_X1 U427 ( .A(n542), .B(a[8]), .ZN(n497) );
  OR2_X1 U428 ( .A1(n228), .A2(n231), .ZN(n498) );
  XNOR2_X1 U429 ( .A(n271), .B(n499), .ZN(n147) );
  XNOR2_X1 U430 ( .A(n289), .B(n279), .ZN(n499) );
  OAI21_X1 U431 ( .B1(n105), .B2(n495), .A(n106), .ZN(n500) );
  XOR2_X1 U432 ( .A(n7), .B(a[4]), .Z(n571) );
  INV_X1 U433 ( .A(n7), .ZN(n601) );
  XOR2_X1 U434 ( .A(n187), .B(n180), .Z(n501) );
  XOR2_X1 U435 ( .A(n178), .B(n501), .Z(n176) );
  NAND2_X1 U436 ( .A1(n178), .A2(n187), .ZN(n502) );
  NAND2_X1 U437 ( .A1(n178), .A2(n180), .ZN(n503) );
  NAND2_X1 U438 ( .A1(n187), .A2(n180), .ZN(n504) );
  NAND3_X1 U439 ( .A1(n502), .A2(n503), .A3(n504), .ZN(n175) );
  XNOR2_X1 U440 ( .A(n188), .B(n505), .ZN(n186) );
  XNOR2_X1 U441 ( .A(n197), .B(n190), .ZN(n505) );
  XOR2_X1 U442 ( .A(n225), .B(n222), .Z(n506) );
  XOR2_X1 U443 ( .A(n220), .B(n506), .Z(n218) );
  NAND2_X1 U444 ( .A1(n220), .A2(n225), .ZN(n507) );
  NAND2_X1 U445 ( .A1(n220), .A2(n222), .ZN(n508) );
  NAND2_X1 U446 ( .A1(n225), .A2(n222), .ZN(n509) );
  NAND3_X1 U447 ( .A1(n507), .A2(n508), .A3(n509), .ZN(n217) );
  NOR2_X2 U448 ( .A1(n218), .A2(n223), .ZN(n97) );
  XNOR2_X1 U449 ( .A(n510), .B(n147), .ZN(n144) );
  XNOR2_X1 U450 ( .A(n301), .B(n148), .ZN(n510) );
  NAND2_X1 U451 ( .A1(n253), .A2(n283), .ZN(n511) );
  NAND2_X1 U452 ( .A1(n253), .A2(n305), .ZN(n512) );
  NAND2_X1 U453 ( .A1(n283), .A2(n305), .ZN(n513) );
  NAND3_X1 U454 ( .A1(n511), .A2(n512), .A3(n513), .ZN(n191) );
  XOR2_X1 U455 ( .A(n193), .B(n282), .Z(n514) );
  XOR2_X1 U456 ( .A(n514), .B(n191), .Z(n180) );
  NAND2_X1 U457 ( .A1(n193), .A2(n282), .ZN(n515) );
  NAND2_X1 U458 ( .A1(n193), .A2(n191), .ZN(n516) );
  NAND2_X1 U459 ( .A1(n282), .A2(n191), .ZN(n517) );
  NAND3_X1 U460 ( .A1(n515), .A2(n516), .A3(n517), .ZN(n179) );
  INV_X1 U461 ( .A(n571), .ZN(n538) );
  NAND2_X1 U462 ( .A1(n188), .A2(n197), .ZN(n518) );
  NAND2_X1 U463 ( .A1(n188), .A2(n190), .ZN(n519) );
  NAND2_X1 U464 ( .A1(n197), .A2(n190), .ZN(n520) );
  NAND3_X1 U465 ( .A1(n518), .A2(n519), .A3(n520), .ZN(n185) );
  INV_X2 U466 ( .A(n541), .ZN(n555) );
  XOR2_X1 U467 ( .A(n541), .B(a[6]), .Z(n563) );
  OR2_X1 U468 ( .A1(n196), .A2(n203), .ZN(n521) );
  INV_X2 U469 ( .A(n497), .ZN(n522) );
  INV_X1 U470 ( .A(n561), .ZN(n27) );
  OR2_X1 U471 ( .A1(n75), .A2(n78), .ZN(n523) );
  INV_X1 U472 ( .A(n523), .ZN(n73) );
  INV_X2 U473 ( .A(n609), .ZN(n608) );
  OR2_X1 U474 ( .A1(n186), .A2(n195), .ZN(n524) );
  INV_X1 U475 ( .A(n601), .ZN(n525) );
  INV_X1 U476 ( .A(n601), .ZN(n600) );
  AOI21_X1 U477 ( .B1(n532), .B2(n80), .A(n81), .ZN(n526) );
  AOI21_X1 U478 ( .B1(n532), .B2(n80), .A(n81), .ZN(n527) );
  NOR2_X1 U479 ( .A1(n164), .A2(n175), .ZN(n528) );
  NOR2_X1 U480 ( .A1(n164), .A2(n175), .ZN(n75) );
  XNOR2_X1 U481 ( .A(n596), .B(a[2]), .ZN(n529) );
  INV_X1 U482 ( .A(n535), .ZN(n530) );
  XOR2_X1 U483 ( .A(n598), .B(a[2]), .Z(n9) );
  CLKBUF_X1 U484 ( .A(n21), .Z(n531) );
  OAI21_X1 U485 ( .B1(n494), .B2(n89), .A(n90), .ZN(n532) );
  BUF_X2 U486 ( .A(n595), .Z(n533) );
  BUF_X2 U487 ( .A(n23), .Z(n534) );
  INV_X1 U488 ( .A(n607), .ZN(n535) );
  NAND2_X1 U489 ( .A1(n577), .A2(n529), .ZN(n536) );
  NAND2_X1 U490 ( .A1(n577), .A2(n529), .ZN(n537) );
  NAND2_X1 U491 ( .A1(n577), .A2(n540), .ZN(n570) );
  INV_X1 U492 ( .A(n571), .ZN(n16) );
  CLKBUF_X1 U493 ( .A(n74), .Z(n539) );
  XNOR2_X1 U494 ( .A(n605), .B(a[8]), .ZN(n429) );
  XNOR2_X1 U495 ( .A(n601), .B(a[2]), .ZN(n577) );
  XNOR2_X1 U496 ( .A(n596), .B(a[2]), .ZN(n540) );
  INV_X1 U497 ( .A(n19), .ZN(n541) );
  INV_X1 U498 ( .A(n19), .ZN(n542) );
  INV_X1 U499 ( .A(n602), .ZN(n543) );
  INV_X2 U500 ( .A(n603), .ZN(n602) );
  CLKBUF_X1 U501 ( .A(n21), .Z(n544) );
  XNOR2_X1 U502 ( .A(n603), .B(a[4]), .ZN(n431) );
  NOR2_X1 U503 ( .A1(n186), .A2(n195), .ZN(n545) );
  INV_X1 U504 ( .A(n607), .ZN(n546) );
  NOR2_X1 U505 ( .A1(n186), .A2(n195), .ZN(n82) );
  INV_X1 U506 ( .A(n607), .ZN(n606) );
  AOI21_X1 U507 ( .B1(n500), .B2(n580), .A(n558), .ZN(n547) );
  BUF_X1 U508 ( .A(n37), .Z(n548) );
  OR2_X2 U509 ( .A1(n549), .A2(n565), .ZN(n34) );
  XNOR2_X1 U510 ( .A(n606), .B(a[10]), .ZN(n549) );
  INV_X1 U511 ( .A(n565), .ZN(n32) );
  XOR2_X1 U512 ( .A(n298), .B(n229), .Z(n550) );
  XOR2_X1 U513 ( .A(n226), .B(n550), .Z(n224) );
  NAND2_X1 U514 ( .A1(n298), .A2(n226), .ZN(n551) );
  NAND2_X1 U515 ( .A1(n226), .A2(n229), .ZN(n552) );
  NAND2_X1 U516 ( .A1(n298), .A2(n229), .ZN(n553) );
  NAND3_X1 U517 ( .A1(n551), .A2(n552), .A3(n553), .ZN(n223) );
  INV_X1 U518 ( .A(n542), .ZN(n554) );
  OR2_X1 U519 ( .A1(n23), .A2(n359), .ZN(n556) );
  OR2_X1 U520 ( .A1(n21), .A2(n358), .ZN(n557) );
  NAND2_X1 U521 ( .A1(n556), .A2(n557), .ZN(n283) );
  INV_X1 U522 ( .A(n558), .ZN(n103) );
  AND2_X1 U523 ( .A1(n224), .A2(n227), .ZN(n558) );
  XNOR2_X1 U524 ( .A(n598), .B(n249), .ZN(n433) );
  NAND2_X1 U525 ( .A1(n431), .A2(n16), .ZN(n559) );
  NAND2_X1 U526 ( .A1(n431), .A2(n16), .ZN(n560) );
  NAND2_X1 U527 ( .A1(n431), .A2(n538), .ZN(n18) );
  XNOR2_X1 U528 ( .A(n542), .B(a[8]), .ZN(n561) );
  INV_X1 U529 ( .A(n575), .ZN(n562) );
  INV_X1 U530 ( .A(n601), .ZN(n599) );
  OR2_X2 U531 ( .A1(n563), .A2(n576), .ZN(n23) );
  INV_X1 U532 ( .A(n576), .ZN(n21) );
  CLKBUF_X1 U533 ( .A(n115), .Z(n564) );
  XNOR2_X1 U534 ( .A(n605), .B(a[10]), .ZN(n565) );
  CLKBUF_X1 U535 ( .A(n107), .Z(n566) );
  OR2_X1 U536 ( .A1(n204), .A2(n211), .ZN(n567) );
  NAND2_X1 U537 ( .A1(n27), .A2(n429), .ZN(n568) );
  NAND2_X1 U538 ( .A1(n429), .A2(n27), .ZN(n569) );
  NAND2_X1 U539 ( .A1(n429), .A2(n522), .ZN(n29) );
  NAND2_X1 U540 ( .A1(n577), .A2(n540), .ZN(n12) );
  INV_X2 U541 ( .A(n605), .ZN(n604) );
  OAI21_X1 U542 ( .B1(n547), .B2(n97), .A(n98), .ZN(n572) );
  NAND2_X1 U543 ( .A1(n433), .A2(n562), .ZN(n573) );
  NAND2_X1 U544 ( .A1(n433), .A2(n562), .ZN(n574) );
  CLKBUF_X1 U545 ( .A(n249), .Z(n575) );
  NAND2_X1 U546 ( .A1(n562), .A2(n433), .ZN(n6) );
  XNOR2_X1 U547 ( .A(n603), .B(a[6]), .ZN(n576) );
  BUF_X1 U548 ( .A(n43), .Z(n593) );
  NAND2_X1 U549 ( .A1(n578), .A2(n69), .ZN(n47) );
  AOI21_X1 U550 ( .B1(n539), .B2(n578), .A(n67), .ZN(n65) );
  INV_X1 U551 ( .A(n69), .ZN(n67) );
  INV_X1 U552 ( .A(n74), .ZN(n72) );
  INV_X1 U553 ( .A(n95), .ZN(n93) );
  XNOR2_X1 U554 ( .A(n84), .B(n50), .ZN(product[11]) );
  NAND2_X1 U555 ( .A1(n524), .A2(n83), .ZN(n50) );
  NAND2_X1 U556 ( .A1(n126), .A2(n79), .ZN(n49) );
  INV_X1 U557 ( .A(n78), .ZN(n126) );
  NAND2_X1 U558 ( .A1(n567), .A2(n90), .ZN(n52) );
  OR2_X1 U559 ( .A1(n152), .A2(n163), .ZN(n578) );
  NAND2_X1 U560 ( .A1(n125), .A2(n76), .ZN(n48) );
  NAND2_X1 U561 ( .A1(n152), .A2(n163), .ZN(n69) );
  NAND2_X1 U562 ( .A1(n579), .A2(n95), .ZN(n53) );
  OAI21_X1 U563 ( .B1(n113), .B2(n115), .A(n114), .ZN(n112) );
  AOI21_X1 U564 ( .B1(n583), .B2(n112), .A(n109), .ZN(n107) );
  AOI21_X1 U565 ( .B1(n580), .B2(n104), .A(n558), .ZN(n99) );
  OAI21_X1 U566 ( .B1(n105), .B2(n107), .A(n106), .ZN(n104) );
  NAND2_X1 U567 ( .A1(n498), .A2(n106), .ZN(n56) );
  NAND2_X1 U568 ( .A1(n131), .A2(n98), .ZN(n54) );
  INV_X1 U569 ( .A(n97), .ZN(n131) );
  AOI21_X1 U570 ( .B1(n581), .B2(n120), .A(n117), .ZN(n115) );
  INV_X1 U571 ( .A(n119), .ZN(n117) );
  NAND2_X1 U572 ( .A1(n580), .A2(n103), .ZN(n55) );
  OAI21_X1 U573 ( .B1(n99), .B2(n97), .A(n98), .ZN(n96) );
  XOR2_X1 U574 ( .A(n58), .B(n564), .Z(product[3]) );
  NAND2_X1 U575 ( .A1(n135), .A2(n114), .ZN(n58) );
  INV_X1 U576 ( .A(n113), .ZN(n135) );
  NOR2_X1 U577 ( .A1(n176), .A2(n185), .ZN(n78) );
  INV_X1 U578 ( .A(n122), .ZN(n120) );
  NOR2_X1 U579 ( .A1(n196), .A2(n203), .ZN(n85) );
  XNOR2_X1 U580 ( .A(n57), .B(n112), .ZN(product[4]) );
  NAND2_X1 U581 ( .A1(n583), .A2(n111), .ZN(n57) );
  NAND2_X1 U582 ( .A1(n176), .A2(n185), .ZN(n79) );
  NAND2_X1 U583 ( .A1(n196), .A2(n203), .ZN(n86) );
  NAND2_X1 U584 ( .A1(n186), .A2(n195), .ZN(n83) );
  NAND2_X1 U585 ( .A1(n212), .A2(n217), .ZN(n95) );
  OR2_X1 U586 ( .A1(n212), .A2(n217), .ZN(n579) );
  XNOR2_X1 U587 ( .A(n59), .B(n120), .ZN(product[2]) );
  NAND2_X1 U588 ( .A1(n581), .A2(n119), .ZN(n59) );
  NAND2_X1 U589 ( .A1(n582), .A2(n62), .ZN(n46) );
  NAND2_X1 U590 ( .A1(n73), .A2(n578), .ZN(n64) );
  OR2_X1 U591 ( .A1(n224), .A2(n227), .ZN(n580) );
  NAND2_X1 U592 ( .A1(n328), .A2(n314), .ZN(n119) );
  OR2_X1 U593 ( .A1(n328), .A2(n314), .ZN(n581) );
  NOR2_X1 U594 ( .A1(n228), .A2(n231), .ZN(n105) );
  OR2_X1 U595 ( .A1(n151), .A2(n139), .ZN(n582) );
  NAND2_X1 U596 ( .A1(n218), .A2(n223), .ZN(n98) );
  NAND2_X1 U597 ( .A1(n228), .A2(n231), .ZN(n106) );
  OR2_X1 U598 ( .A1(n232), .A2(n233), .ZN(n583) );
  INV_X1 U599 ( .A(n37), .ZN(n237) );
  NAND2_X1 U600 ( .A1(n232), .A2(n233), .ZN(n111) );
  INV_X1 U601 ( .A(n41), .ZN(n235) );
  AND2_X1 U602 ( .A1(n490), .A2(n122), .ZN(product[1]) );
  XNOR2_X1 U603 ( .A(n606), .B(a[12]), .ZN(n37) );
  XNOR2_X1 U604 ( .A(n608), .B(a[14]), .ZN(n41) );
  INV_X1 U605 ( .A(n249), .ZN(n595) );
  OR2_X1 U606 ( .A1(n593), .A2(n496), .ZN(n392) );
  OAI22_X1 U607 ( .A1(n39), .A2(n336), .B1(n548), .B2(n335), .ZN(n263) );
  AND2_X1 U608 ( .A1(n594), .A2(n565), .ZN(n270) );
  AND2_X1 U609 ( .A1(n594), .A2(n571), .ZN(n300) );
  XNOR2_X1 U610 ( .A(n602), .B(n593), .ZN(n376) );
  XNOR2_X1 U611 ( .A(n599), .B(n593), .ZN(n391) );
  OAI22_X1 U612 ( .A1(n39), .A2(n609), .B1(n337), .B2(n548), .ZN(n252) );
  OR2_X1 U613 ( .A1(n593), .A2(n609), .ZN(n337) );
  OAI22_X1 U614 ( .A1(n42), .A2(n611), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U615 ( .A1(n593), .A2(n611), .ZN(n332) );
  XNOR2_X1 U616 ( .A(n155), .B(n585), .ZN(n139) );
  XNOR2_X1 U617 ( .A(n153), .B(n141), .ZN(n585) );
  XNOR2_X1 U618 ( .A(n157), .B(n586), .ZN(n141) );
  XNOR2_X1 U619 ( .A(n145), .B(n143), .ZN(n586) );
  XNOR2_X1 U620 ( .A(n159), .B(n587), .ZN(n142) );
  XNOR2_X1 U621 ( .A(n315), .B(n261), .ZN(n587) );
  XNOR2_X1 U622 ( .A(n608), .B(n593), .ZN(n336) );
  AND2_X1 U623 ( .A1(n594), .A2(n247), .ZN(n314) );
  AND2_X1 U624 ( .A1(n594), .A2(n561), .ZN(n278) );
  AND2_X1 U625 ( .A1(n594), .A2(n237), .ZN(n264) );
  AND2_X1 U626 ( .A1(n594), .A2(n576), .ZN(n288) );
  AND2_X1 U627 ( .A1(n594), .A2(n235), .ZN(n260) );
  OAI22_X1 U628 ( .A1(n39), .A2(n335), .B1(n548), .B2(n334), .ZN(n262) );
  NAND2_X1 U629 ( .A1(n427), .A2(n37), .ZN(n39) );
  XOR2_X1 U630 ( .A(n608), .B(a[12]), .Z(n427) );
  INV_X1 U631 ( .A(n25), .ZN(n605) );
  INV_X1 U632 ( .A(n13), .ZN(n603) );
  XNOR2_X1 U633 ( .A(n604), .B(n593), .ZN(n352) );
  NAND2_X1 U634 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U635 ( .A(n610), .B(a[14]), .Z(n426) );
  XNOR2_X1 U636 ( .A(n554), .B(n593), .ZN(n363) );
  AND2_X1 U637 ( .A1(n594), .A2(n575), .ZN(product[0]) );
  OR2_X1 U638 ( .A1(n593), .A2(n605), .ZN(n353) );
  OR2_X1 U639 ( .A1(n593), .A2(n541), .ZN(n364) );
  OR2_X1 U640 ( .A1(n593), .A2(n530), .ZN(n344) );
  OR2_X1 U641 ( .A1(n593), .A2(n543), .ZN(n377) );
  XNOR2_X1 U642 ( .A(n554), .B(b[9]), .ZN(n354) );
  XNOR2_X1 U643 ( .A(n602), .B(b[11]), .ZN(n365) );
  OAI22_X1 U644 ( .A1(n39), .A2(n334), .B1(n548), .B2(n333), .ZN(n261) );
  XNOR2_X1 U645 ( .A(n608), .B(n422), .ZN(n333) );
  XNOR2_X1 U646 ( .A(n608), .B(n423), .ZN(n334) );
  XNOR2_X1 U647 ( .A(n608), .B(n424), .ZN(n335) );
  OAI22_X1 U648 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U649 ( .A(n610), .B(n424), .ZN(n330) );
  XNOR2_X1 U650 ( .A(n610), .B(n593), .ZN(n331) );
  XNOR2_X1 U651 ( .A(n599), .B(b[13]), .ZN(n378) );
  XNOR2_X1 U652 ( .A(n604), .B(n418), .ZN(n345) );
  XNOR2_X1 U653 ( .A(n546), .B(n420), .ZN(n338) );
  XNOR2_X1 U654 ( .A(n599), .B(n424), .ZN(n390) );
  XNOR2_X1 U655 ( .A(n554), .B(n424), .ZN(n362) );
  XNOR2_X1 U656 ( .A(n604), .B(n424), .ZN(n351) );
  XNOR2_X1 U657 ( .A(n525), .B(n418), .ZN(n384) );
  XNOR2_X1 U658 ( .A(n600), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U659 ( .A(n599), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U660 ( .A(n599), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U661 ( .A(n525), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U662 ( .A(n599), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U663 ( .A(n525), .B(n419), .ZN(n385) );
  XNOR2_X1 U664 ( .A(n602), .B(n418), .ZN(n369) );
  XNOR2_X1 U665 ( .A(n602), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U666 ( .A(n602), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U667 ( .A(n602), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U668 ( .A(n600), .B(n423), .ZN(n389) );
  XNOR2_X1 U669 ( .A(n555), .B(n423), .ZN(n361) );
  XNOR2_X1 U670 ( .A(n604), .B(n423), .ZN(n350) );
  XNOR2_X1 U671 ( .A(n525), .B(n421), .ZN(n387) );
  XNOR2_X1 U672 ( .A(n555), .B(n421), .ZN(n359) );
  XNOR2_X1 U673 ( .A(n604), .B(n421), .ZN(n348) );
  XNOR2_X1 U674 ( .A(n555), .B(n420), .ZN(n358) );
  XNOR2_X1 U675 ( .A(n525), .B(n420), .ZN(n386) );
  XNOR2_X1 U676 ( .A(n604), .B(n420), .ZN(n347) );
  XNOR2_X1 U677 ( .A(n555), .B(n418), .ZN(n356) );
  XNOR2_X1 U678 ( .A(n604), .B(n419), .ZN(n346) );
  XNOR2_X1 U679 ( .A(n554), .B(n419), .ZN(n357) );
  XNOR2_X1 U680 ( .A(n597), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U681 ( .A(n600), .B(n422), .ZN(n388) );
  XNOR2_X1 U682 ( .A(n592), .B(b[13]), .ZN(n395) );
  XNOR2_X1 U683 ( .A(n555), .B(b[8]), .ZN(n355) );
  XNOR2_X1 U684 ( .A(n591), .B(b[11]), .ZN(n397) );
  XNOR2_X1 U685 ( .A(n591), .B(b[14]), .ZN(n394) );
  XNOR2_X1 U686 ( .A(n554), .B(n422), .ZN(n360) );
  XNOR2_X1 U687 ( .A(n604), .B(n422), .ZN(n349) );
  XNOR2_X1 U688 ( .A(n546), .B(n422), .ZN(n340) );
  BUF_X1 U689 ( .A(n43), .Z(n594) );
  XNOR2_X1 U690 ( .A(n597), .B(b[15]), .ZN(n393) );
  XNOR2_X1 U691 ( .A(n535), .B(n424), .ZN(n342) );
  XNOR2_X1 U692 ( .A(n535), .B(n423), .ZN(n341) );
  XNOR2_X1 U693 ( .A(n546), .B(n593), .ZN(n343) );
  XNOR2_X1 U694 ( .A(n546), .B(n421), .ZN(n339) );
  INV_X1 U695 ( .A(n597), .ZN(n590) );
  INV_X1 U696 ( .A(n75), .ZN(n125) );
  OAI21_X1 U697 ( .B1(n528), .B2(n79), .A(n76), .ZN(n74) );
  NAND2_X1 U698 ( .A1(n164), .A2(n175), .ZN(n76) );
  OAI22_X1 U699 ( .A1(n34), .A2(n339), .B1(n338), .B2(n32), .ZN(n265) );
  OAI22_X1 U700 ( .A1(n34), .A2(n340), .B1(n339), .B2(n32), .ZN(n266) );
  OAI22_X1 U701 ( .A1(n34), .A2(n342), .B1(n341), .B2(n32), .ZN(n268) );
  OAI22_X1 U702 ( .A1(n34), .A2(n343), .B1(n342), .B2(n32), .ZN(n269) );
  OAI22_X1 U703 ( .A1(n34), .A2(n341), .B1(n340), .B2(n32), .ZN(n267) );
  OAI22_X1 U704 ( .A1(n34), .A2(n530), .B1(n344), .B2(n32), .ZN(n253) );
  OAI22_X1 U705 ( .A1(n573), .A2(n394), .B1(n393), .B2(n533), .ZN(n315) );
  OAI22_X1 U706 ( .A1(n574), .A2(n395), .B1(n394), .B2(n533), .ZN(n316) );
  OAI22_X1 U707 ( .A1(n573), .A2(n400), .B1(n399), .B2(n533), .ZN(n321) );
  OAI22_X1 U708 ( .A1(n574), .A2(n401), .B1(n400), .B2(n533), .ZN(n322) );
  OAI22_X1 U709 ( .A1(n6), .A2(n402), .B1(n401), .B2(n533), .ZN(n323) );
  OAI22_X1 U710 ( .A1(n574), .A2(n397), .B1(n396), .B2(n533), .ZN(n318) );
  OAI22_X1 U711 ( .A1(n573), .A2(n398), .B1(n397), .B2(n533), .ZN(n319) );
  OAI22_X1 U712 ( .A1(n573), .A2(n396), .B1(n395), .B2(n533), .ZN(n317) );
  OAI22_X1 U713 ( .A1(n6), .A2(n399), .B1(n398), .B2(n533), .ZN(n320) );
  OAI22_X1 U714 ( .A1(n6), .A2(n404), .B1(n403), .B2(n533), .ZN(n325) );
  OAI22_X1 U715 ( .A1(n6), .A2(n405), .B1(n404), .B2(n533), .ZN(n326) );
  OAI22_X1 U716 ( .A1(n574), .A2(n406), .B1(n405), .B2(n533), .ZN(n327) );
  OAI22_X1 U717 ( .A1(n574), .A2(n403), .B1(n402), .B2(n533), .ZN(n324) );
  OAI22_X1 U718 ( .A1(n573), .A2(n407), .B1(n406), .B2(n533), .ZN(n328) );
  OAI22_X1 U719 ( .A1(n573), .A2(n408), .B1(n407), .B2(n533), .ZN(n329) );
  NAND2_X1 U720 ( .A1(n204), .A2(n211), .ZN(n90) );
  NOR2_X1 U721 ( .A1(n204), .A2(n211), .ZN(n89) );
  OAI22_X1 U722 ( .A1(n568), .A2(n346), .B1(n345), .B2(n522), .ZN(n271) );
  OAI22_X1 U723 ( .A1(n568), .A2(n350), .B1(n349), .B2(n522), .ZN(n275) );
  OAI22_X1 U724 ( .A1(n569), .A2(n347), .B1(n346), .B2(n522), .ZN(n272) );
  OAI22_X1 U725 ( .A1(n569), .A2(n351), .B1(n350), .B2(n522), .ZN(n276) );
  OAI22_X1 U726 ( .A1(n569), .A2(n349), .B1(n348), .B2(n522), .ZN(n274) );
  OAI22_X1 U727 ( .A1(n568), .A2(n348), .B1(n347), .B2(n522), .ZN(n273) );
  OAI22_X1 U728 ( .A1(n568), .A2(n605), .B1(n353), .B2(n522), .ZN(n254) );
  OAI22_X1 U729 ( .A1(n29), .A2(n352), .B1(n351), .B2(n522), .ZN(n277) );
  INV_X1 U730 ( .A(n598), .ZN(n591) );
  INV_X1 U731 ( .A(n598), .ZN(n592) );
  INV_X1 U732 ( .A(n598), .ZN(n596) );
  XNOR2_X1 U733 ( .A(n63), .B(n46), .ZN(product[15]) );
  XNOR2_X1 U734 ( .A(n77), .B(n48), .ZN(product[13]) );
  OR2_X1 U735 ( .A1(n593), .A2(n590), .ZN(n409) );
  INV_X1 U736 ( .A(n598), .ZN(n597) );
  XNOR2_X1 U737 ( .A(n70), .B(n47), .ZN(product[14]) );
  NOR2_X1 U738 ( .A1(n82), .A2(n85), .ZN(n80) );
  OAI21_X1 U739 ( .B1(n86), .B2(n545), .A(n83), .ZN(n81) );
  XNOR2_X1 U740 ( .A(n602), .B(n424), .ZN(n375) );
  XNOR2_X1 U741 ( .A(n602), .B(n423), .ZN(n374) );
  XNOR2_X1 U742 ( .A(n602), .B(n421), .ZN(n372) );
  XNOR2_X1 U743 ( .A(n602), .B(n422), .ZN(n373) );
  XNOR2_X1 U744 ( .A(n602), .B(n419), .ZN(n370) );
  XNOR2_X1 U745 ( .A(n602), .B(n420), .ZN(n371) );
  OAI21_X1 U746 ( .B1(n87), .B2(n85), .A(n492), .ZN(n84) );
  XNOR2_X1 U747 ( .A(n572), .B(n53), .ZN(product[8]) );
  NOR2_X1 U748 ( .A1(n234), .A2(n257), .ZN(n113) );
  OAI21_X1 U749 ( .B1(n91), .B2(n89), .A(n90), .ZN(n88) );
  XOR2_X1 U750 ( .A(n547), .B(n54), .Z(product[7]) );
  INV_X1 U751 ( .A(n88), .ZN(n87) );
  OAI22_X1 U752 ( .A1(n534), .A2(n358), .B1(n357), .B2(n544), .ZN(n282) );
  OAI22_X1 U753 ( .A1(n534), .A2(n356), .B1(n355), .B2(n544), .ZN(n280) );
  OAI22_X1 U754 ( .A1(n534), .A2(n360), .B1(n359), .B2(n531), .ZN(n284) );
  OAI22_X1 U755 ( .A1(n534), .A2(n357), .B1(n356), .B2(n531), .ZN(n281) );
  OAI22_X1 U756 ( .A1(n534), .A2(n355), .B1(n354), .B2(n531), .ZN(n279) );
  OAI22_X1 U757 ( .A1(n534), .A2(n362), .B1(n361), .B2(n544), .ZN(n286) );
  OAI22_X1 U758 ( .A1(n23), .A2(n361), .B1(n360), .B2(n21), .ZN(n285) );
  OAI22_X1 U759 ( .A1(n23), .A2(n542), .B1(n364), .B2(n21), .ZN(n255) );
  OAI22_X1 U760 ( .A1(n23), .A2(n363), .B1(n362), .B2(n21), .ZN(n287) );
  XNOR2_X1 U761 ( .A(n592), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U762 ( .A(n597), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U763 ( .A(n591), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U764 ( .A(n592), .B(n418), .ZN(n401) );
  XNOR2_X1 U765 ( .A(n597), .B(n593), .ZN(n408) );
  XNOR2_X1 U766 ( .A(n592), .B(n419), .ZN(n402) );
  XNOR2_X1 U767 ( .A(n591), .B(n420), .ZN(n403) );
  XNOR2_X1 U768 ( .A(n592), .B(n422), .ZN(n405) );
  XNOR2_X1 U769 ( .A(n592), .B(n424), .ZN(n407) );
  XNOR2_X1 U770 ( .A(n597), .B(n423), .ZN(n406) );
  XNOR2_X1 U771 ( .A(n591), .B(n421), .ZN(n404) );
  OAI21_X1 U772 ( .B1(n64), .B2(n527), .A(n65), .ZN(n63) );
  OAI21_X1 U773 ( .B1(n527), .B2(n78), .A(n79), .ZN(n77) );
  XNOR2_X1 U774 ( .A(n55), .B(n500), .ZN(product[6]) );
  NAND2_X1 U775 ( .A1(n151), .A2(n139), .ZN(n62) );
  OAI22_X1 U776 ( .A1(n559), .A2(n367), .B1(n366), .B2(n538), .ZN(n290) );
  OAI22_X1 U777 ( .A1(n560), .A2(n370), .B1(n369), .B2(n538), .ZN(n293) );
  OAI22_X1 U778 ( .A1(n559), .A2(n375), .B1(n374), .B2(n538), .ZN(n298) );
  OAI22_X1 U779 ( .A1(n559), .A2(n368), .B1(n367), .B2(n538), .ZN(n291) );
  OAI22_X1 U780 ( .A1(n560), .A2(n373), .B1(n372), .B2(n538), .ZN(n296) );
  OAI22_X1 U781 ( .A1(n559), .A2(n369), .B1(n368), .B2(n538), .ZN(n292) );
  OAI22_X1 U782 ( .A1(n18), .A2(n374), .B1(n373), .B2(n538), .ZN(n297) );
  OAI22_X1 U783 ( .A1(n560), .A2(n372), .B1(n371), .B2(n16), .ZN(n295) );
  OAI22_X1 U784 ( .A1(n559), .A2(n543), .B1(n377), .B2(n538), .ZN(n256) );
  OAI22_X1 U785 ( .A1(n560), .A2(n376), .B1(n375), .B2(n538), .ZN(n299) );
  OAI22_X1 U786 ( .A1(n18), .A2(n371), .B1(n370), .B2(n538), .ZN(n294) );
  OAI22_X1 U787 ( .A1(n560), .A2(n366), .B1(n365), .B2(n538), .ZN(n289) );
  OAI21_X1 U788 ( .B1(n527), .B2(n523), .A(n72), .ZN(n70) );
  XOR2_X1 U789 ( .A(n526), .B(n49), .Z(product[12]) );
  XOR2_X1 U790 ( .A(n494), .B(n52), .Z(product[9]) );
  XOR2_X1 U791 ( .A(n56), .B(n566), .Z(product[5]) );
  NAND2_X1 U792 ( .A1(n329), .A2(n258), .ZN(n122) );
  INV_X1 U793 ( .A(n111), .ZN(n109) );
  OAI22_X1 U794 ( .A1(n574), .A2(n590), .B1(n409), .B2(n533), .ZN(n258) );
  OAI22_X1 U795 ( .A1(n12), .A2(n379), .B1(n378), .B2(n588), .ZN(n301) );
  OAI22_X1 U796 ( .A1(n12), .A2(n380), .B1(n379), .B2(n588), .ZN(n302) );
  OAI22_X1 U797 ( .A1(n536), .A2(n385), .B1(n384), .B2(n588), .ZN(n307) );
  OAI22_X1 U798 ( .A1(n537), .A2(n382), .B1(n381), .B2(n588), .ZN(n304) );
  OAI22_X1 U799 ( .A1(n12), .A2(n381), .B1(n380), .B2(n588), .ZN(n303) );
  NAND2_X1 U800 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U801 ( .A1(n570), .A2(n383), .B1(n382), .B2(n588), .ZN(n305) );
  OAI22_X1 U802 ( .A1(n570), .A2(n384), .B1(n383), .B2(n589), .ZN(n306) );
  OAI22_X1 U803 ( .A1(n536), .A2(n386), .B1(n385), .B2(n588), .ZN(n308) );
  OAI22_X1 U804 ( .A1(n537), .A2(n387), .B1(n386), .B2(n588), .ZN(n309) );
  OAI22_X1 U805 ( .A1(n537), .A2(n496), .B1(n392), .B2(n588), .ZN(n257) );
  OAI22_X1 U806 ( .A1(n570), .A2(n389), .B1(n388), .B2(n589), .ZN(n311) );
  OAI22_X1 U807 ( .A1(n536), .A2(n388), .B1(n387), .B2(n589), .ZN(n310) );
  OAI22_X1 U808 ( .A1(n536), .A2(n390), .B1(n389), .B2(n589), .ZN(n312) );
  INV_X1 U809 ( .A(n588), .ZN(n247) );
  OAI22_X1 U810 ( .A1(n12), .A2(n391), .B1(n390), .B2(n589), .ZN(n313) );
  INV_X1 U811 ( .A(n31), .ZN(n607) );
  INV_X1 U812 ( .A(n36), .ZN(n609) );
  INV_X1 U813 ( .A(n611), .ZN(n610) );
  INV_X1 U814 ( .A(n40), .ZN(n611) );
  XOR2_X1 U815 ( .A(n259), .B(n251), .Z(n148) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_1_DW01_add_2 ( A, B, CI, SUM, 
        CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n18,
         n19, n20, n21, n23, n25, n26, n27, n28, n30, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n48, n49, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n71, n72, n73,
         n74, n75, n77, n79, n80, n81, n82, n83, n85, n87, n88, n90, n93, n94,
         n95, n99, n100, n102, n104, n161, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180;

  OR2_X1 U126 ( .A1(A[8]), .A2(B[8]), .ZN(n161) );
  AND2_X1 U127 ( .A1(n174), .A2(n90), .ZN(SUM[0]) );
  OR2_X1 U128 ( .A1(A[15]), .A2(B[15]), .ZN(n163) );
  BUF_X1 U129 ( .A(n171), .Z(n164) );
  OR2_X1 U130 ( .A1(A[10]), .A2(B[10]), .ZN(n165) );
  OR2_X1 U131 ( .A1(A[10]), .A2(B[10]), .ZN(n166) );
  OR2_X1 U132 ( .A1(A[10]), .A2(B[10]), .ZN(n180) );
  AND2_X1 U133 ( .A1(A[9]), .A2(B[9]), .ZN(n167) );
  BUF_X1 U134 ( .A(n42), .Z(n169) );
  NOR2_X1 U135 ( .A1(A[12]), .A2(B[12]), .ZN(n168) );
  NOR2_X1 U136 ( .A1(A[12]), .A2(B[12]), .ZN(n36) );
  OAI21_X1 U137 ( .B1(n168), .B2(n40), .A(n37), .ZN(n170) );
  INV_X1 U138 ( .A(n164), .ZN(n48) );
  AND2_X1 U139 ( .A1(A[10]), .A2(B[10]), .ZN(n171) );
  AOI21_X1 U140 ( .B1(n42), .B2(n34), .A(n35), .ZN(n172) );
  AOI21_X1 U141 ( .B1(n169), .B2(n34), .A(n170), .ZN(n173) );
  OR2_X1 U142 ( .A1(A[0]), .A2(B[0]), .ZN(n174) );
  INV_X1 U143 ( .A(n64), .ZN(n63) );
  INV_X1 U144 ( .A(n55), .ZN(n54) );
  AOI21_X1 U145 ( .B1(n169), .B2(n34), .A(n170), .ZN(n33) );
  AOI21_X1 U146 ( .B1(n178), .B2(n72), .A(n69), .ZN(n67) );
  INV_X1 U147 ( .A(n71), .ZN(n69) );
  AOI21_X1 U148 ( .B1(n177), .B2(n80), .A(n77), .ZN(n75) );
  INV_X1 U149 ( .A(n79), .ZN(n77) );
  AOI21_X1 U150 ( .B1(n179), .B2(n88), .A(n85), .ZN(n83) );
  INV_X1 U151 ( .A(n87), .ZN(n85) );
  OAI21_X1 U152 ( .B1(n75), .B2(n73), .A(n74), .ZN(n72) );
  OAI21_X1 U153 ( .B1(n83), .B2(n81), .A(n82), .ZN(n80) );
  OAI21_X1 U154 ( .B1(n67), .B2(n65), .A(n66), .ZN(n64) );
  NAND2_X1 U155 ( .A1(n175), .A2(n93), .ZN(n20) );
  AOI21_X1 U156 ( .B1(n175), .B2(n30), .A(n23), .ZN(n21) );
  AOI21_X1 U157 ( .B1(n54), .B2(n176), .A(n167), .ZN(n49) );
  AOI21_X1 U158 ( .B1(n56), .B2(n64), .A(n57), .ZN(n55) );
  NOR2_X1 U159 ( .A1(n58), .A2(n61), .ZN(n56) );
  OAI21_X1 U160 ( .B1(n58), .B2(n62), .A(n59), .ZN(n57) );
  INV_X1 U161 ( .A(n90), .ZN(n88) );
  OAI21_X1 U162 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  INV_X1 U163 ( .A(n25), .ZN(n23) );
  NAND2_X1 U164 ( .A1(n161), .A2(n59), .ZN(n8) );
  NAND2_X1 U165 ( .A1(n100), .A2(n66), .ZN(n10) );
  INV_X1 U166 ( .A(n65), .ZN(n100) );
  NAND2_X1 U167 ( .A1(n102), .A2(n74), .ZN(n12) );
  INV_X1 U168 ( .A(n73), .ZN(n102) );
  INV_X1 U169 ( .A(n168), .ZN(n94) );
  NAND2_X1 U170 ( .A1(n176), .A2(n53), .ZN(n7) );
  NAND2_X1 U171 ( .A1(n99), .A2(n62), .ZN(n9) );
  INV_X1 U172 ( .A(n61), .ZN(n99) );
  NAND2_X1 U173 ( .A1(n104), .A2(n82), .ZN(n14) );
  INV_X1 U174 ( .A(n81), .ZN(n104) );
  NAND2_X1 U175 ( .A1(n178), .A2(n71), .ZN(n11) );
  NAND2_X1 U176 ( .A1(n177), .A2(n79), .ZN(n13) );
  NAND2_X1 U177 ( .A1(n179), .A2(n87), .ZN(n15) );
  XNOR2_X1 U178 ( .A(n13), .B(n80), .ZN(SUM[3]) );
  NAND2_X1 U179 ( .A1(n94), .A2(n37), .ZN(n4) );
  NOR2_X1 U180 ( .A1(A[7]), .A2(B[7]), .ZN(n61) );
  NOR2_X1 U181 ( .A1(A[8]), .A2(B[8]), .ZN(n58) );
  OR2_X1 U182 ( .A1(A[14]), .A2(B[14]), .ZN(n175) );
  OR2_X1 U183 ( .A1(A[9]), .A2(B[9]), .ZN(n176) );
  NOR2_X1 U184 ( .A1(A[2]), .A2(B[2]), .ZN(n81) );
  NOR2_X1 U185 ( .A1(A[4]), .A2(B[4]), .ZN(n73) );
  NOR2_X1 U186 ( .A1(A[6]), .A2(B[6]), .ZN(n65) );
  NAND2_X1 U187 ( .A1(n175), .A2(n25), .ZN(n2) );
  XOR2_X1 U188 ( .A(n49), .B(n6), .Z(SUM[10]) );
  OR2_X1 U189 ( .A1(A[3]), .A2(B[3]), .ZN(n177) );
  OR2_X1 U190 ( .A1(A[5]), .A2(B[5]), .ZN(n178) );
  OR2_X1 U191 ( .A1(A[1]), .A2(B[1]), .ZN(n179) );
  NAND2_X1 U192 ( .A1(A[7]), .A2(B[7]), .ZN(n62) );
  XNOR2_X1 U193 ( .A(n54), .B(n7), .ZN(SUM[9]) );
  XNOR2_X1 U194 ( .A(n11), .B(n72), .ZN(SUM[5]) );
  NAND2_X1 U195 ( .A1(A[8]), .A2(B[8]), .ZN(n59) );
  NAND2_X1 U196 ( .A1(A[2]), .A2(B[2]), .ZN(n82) );
  NAND2_X1 U197 ( .A1(A[4]), .A2(B[4]), .ZN(n74) );
  NAND2_X1 U198 ( .A1(A[6]), .A2(B[6]), .ZN(n66) );
  NAND2_X1 U199 ( .A1(A[3]), .A2(B[3]), .ZN(n79) );
  NAND2_X1 U200 ( .A1(A[5]), .A2(B[5]), .ZN(n71) );
  NAND2_X1 U201 ( .A1(A[1]), .A2(B[1]), .ZN(n87) );
  NAND2_X1 U202 ( .A1(A[0]), .A2(B[0]), .ZN(n90) );
  NAND2_X1 U203 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  NAND2_X1 U204 ( .A1(A[12]), .A2(B[12]), .ZN(n37) );
  XNOR2_X1 U205 ( .A(n60), .B(n8), .ZN(SUM[8]) );
  XOR2_X1 U206 ( .A(n63), .B(n9), .Z(SUM[7]) );
  XOR2_X1 U207 ( .A(n10), .B(n67), .Z(SUM[6]) );
  XOR2_X1 U208 ( .A(n12), .B(n75), .Z(SUM[4]) );
  XOR2_X1 U209 ( .A(n14), .B(n83), .Z(SUM[2]) );
  XNOR2_X1 U210 ( .A(n15), .B(n88), .ZN(SUM[1]) );
  NAND2_X1 U211 ( .A1(n163), .A2(n18), .ZN(n1) );
  NAND2_X1 U212 ( .A1(A[15]), .A2(B[15]), .ZN(n18) );
  NAND2_X1 U213 ( .A1(A[9]), .A2(B[9]), .ZN(n53) );
  NAND2_X1 U214 ( .A1(n93), .A2(n28), .ZN(n3) );
  INV_X1 U215 ( .A(n28), .ZN(n30) );
  INV_X1 U216 ( .A(n27), .ZN(n93) );
  OAI21_X1 U217 ( .B1(n36), .B2(n40), .A(n37), .ZN(n35) );
  NAND2_X1 U218 ( .A1(n95), .A2(n40), .ZN(n5) );
  NAND2_X1 U219 ( .A1(A[11]), .A2(B[11]), .ZN(n40) );
  NOR2_X1 U220 ( .A1(n36), .A2(n39), .ZN(n34) );
  INV_X1 U221 ( .A(n39), .ZN(n95) );
  NOR2_X1 U222 ( .A1(A[11]), .A2(B[11]), .ZN(n39) );
  NAND2_X1 U223 ( .A1(A[14]), .A2(B[14]), .ZN(n25) );
  AOI21_X1 U224 ( .B1(n165), .B2(n167), .A(n171), .ZN(n44) );
  NAND2_X1 U225 ( .A1(n180), .A2(n176), .ZN(n43) );
  NAND2_X1 U226 ( .A1(n166), .A2(n48), .ZN(n6) );
  XOR2_X1 U227 ( .A(n41), .B(n5), .Z(SUM[11]) );
  OAI21_X1 U228 ( .B1(n41), .B2(n39), .A(n40), .ZN(n38) );
  XNOR2_X1 U229 ( .A(n26), .B(n2), .ZN(SUM[14]) );
  INV_X1 U230 ( .A(n42), .ZN(n41) );
  XNOR2_X1 U231 ( .A(n19), .B(n1), .ZN(SUM[15]) );
  NOR2_X1 U232 ( .A1(A[13]), .A2(B[13]), .ZN(n27) );
  XNOR2_X1 U233 ( .A(n38), .B(n4), .ZN(SUM[12]) );
  XOR2_X1 U234 ( .A(n33), .B(n3), .Z(SUM[13]) );
  OAI21_X1 U235 ( .B1(n172), .B2(n27), .A(n28), .ZN(n26) );
  OAI21_X1 U236 ( .B1(n173), .B2(n20), .A(n21), .ZN(n19) );
  OAI21_X1 U237 ( .B1(n43), .B2(n55), .A(n44), .ZN(n42) );
endmodule


module layer2_12_8_12_16_datapath_M12_N8_T16_P12_1 ( clk, clear_acc, 
        data_out_x, data_out, data_out_w, data_out_b, wr_en_y, m_valid, 
        m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [3:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N27, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, n1, n2, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n87, n104, n113, n114, n115, n116, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n13), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n217), .CK(clk), .Q(n18) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n218), .CK(clk), .Q(n19) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n219), .CK(clk), .Q(n20) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n220), .CK(clk), .Q(n21) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n221), .CK(clk), .Q(n22) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n222), .CK(clk), .Q(n23) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n223), .CK(clk), .Q(n24) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n224), .CK(clk), .Q(n25) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n225), .CK(clk), .Q(n26) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n226), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n227), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n228), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n229), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n230), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n231), .CK(clk), .Q(n34) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n232), .CK(clk), .Q(n36) );
  DFF_X1 \f_reg[8]  ( .D(n78), .CK(clk), .Q(f[8]), .QN(n210) );
  DFF_X1 \f_reg[9]  ( .D(n77), .CK(clk), .Q(f[9]), .QN(n211) );
  DFF_X1 \f_reg[10]  ( .D(n76), .CK(clk), .Q(n47), .QN(n212) );
  DFF_X1 \f_reg[11]  ( .D(n75), .CK(clk), .Q(n45), .QN(n213) );
  DFF_X1 \f_reg[12]  ( .D(n74), .CK(clk), .Q(n43), .QN(n214) );
  DFF_X1 \f_reg[13]  ( .D(n73), .CK(clk), .Q(n41), .QN(n215) );
  DFF_X1 \f_reg[14]  ( .D(n1), .CK(clk), .Q(n40), .QN(n216) );
  DFF_X1 \f_reg[15]  ( .D(n2), .CK(clk), .Q(f[15]), .QN(n71) );
  DFF_X1 \data_out_reg[15]  ( .D(n104), .CK(clk), .Q(data_out[15]), .QN(n189)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n113), .CK(clk), .Q(data_out[14]), .QN(n188)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n114), .CK(clk), .Q(data_out[13]), .QN(n187)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n115), .CK(clk), .Q(data_out[12]), .QN(n186)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n116), .CK(clk), .Q(data_out[11]), .QN(n185)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n163), .CK(clk), .Q(data_out[10]), .QN(n184)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n164), .CK(clk), .Q(data_out[9]), .QN(n183) );
  DFF_X1 \data_out_reg[8]  ( .D(n165), .CK(clk), .Q(data_out[8]), .QN(n182) );
  DFF_X1 \data_out_reg[7]  ( .D(n166), .CK(clk), .Q(data_out[7]), .QN(n181) );
  DFF_X1 \data_out_reg[6]  ( .D(n167), .CK(clk), .Q(data_out[6]), .QN(n180) );
  DFF_X1 \data_out_reg[5]  ( .D(n168), .CK(clk), .Q(data_out[5]), .QN(n179) );
  DFF_X1 \data_out_reg[4]  ( .D(n169), .CK(clk), .Q(data_out[4]), .QN(n178) );
  DFF_X1 \data_out_reg[3]  ( .D(n170), .CK(clk), .Q(data_out[3]), .QN(n177) );
  DFF_X1 \data_out_reg[2]  ( .D(n171), .CK(clk), .Q(data_out[2]), .QN(n176) );
  DFF_X1 \data_out_reg[1]  ( .D(n172), .CK(clk), .Q(data_out[1]), .QN(n175) );
  DFF_X1 \data_out_reg[0]  ( .D(n173), .CK(clk), .Q(data_out[0]), .QN(n174) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_1_DW_mult_tc_1 mult_960 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_1_DW01_add_2 add_961 ( .A({n196, 
        n195, n194, n193, n192, n191, n205, n204, n203, n202, n201, n200, n199, 
        n198, n197, n190}), .B({f[15], n40, n41, n43, n45, n47, f[9:3], n55, 
        n57, n59}), .CI(1'b0), .SUM(adder) );
  DFF_X2 delay_reg ( .D(N27), .CK(clk), .Q(n7), .QN(n233) );
  DFF_X1 \f_reg[4]  ( .D(n82), .CK(clk), .Q(f[4]), .QN(n64) );
  DFF_X1 \f_reg[2]  ( .D(n84), .CK(clk), .Q(n55), .QN(n208) );
  DFF_X1 \f_reg[1]  ( .D(n85), .CK(clk), .Q(n57), .QN(n207) );
  DFF_X1 \f_reg[3]  ( .D(n83), .CK(clk), .Q(f[3]), .QN(n63) );
  DFF_X1 \f_reg[0]  ( .D(n87), .CK(clk), .Q(n59), .QN(n206) );
  DFF_X1 \f_reg[5]  ( .D(n81), .CK(clk), .Q(f[5]), .QN(n65) );
  DFF_X1 \f_reg[6]  ( .D(n80), .CK(clk), .Q(f[6]), .QN(n66) );
  DFF_X1 \f_reg[7]  ( .D(n79), .CK(clk), .Q(f[7]), .QN(n209) );
  MUX2_X2 U3 ( .A(N39), .B(n23), .S(n7), .Z(n191) );
  MUX2_X2 U4 ( .A(n25), .B(N37), .S(n233), .Z(n204) );
  MUX2_X1 U5 ( .A(N42), .B(n20), .S(n7), .Z(n194) );
  AND2_X2 U6 ( .A1(n39), .A2(n14), .ZN(n11) );
  NAND3_X1 U8 ( .A1(n5), .A2(n4), .A3(n6), .ZN(n1) );
  NAND3_X1 U9 ( .A1(n9), .A2(n8), .A3(n10), .ZN(n2) );
  NAND2_X1 U10 ( .A1(data_out_b[14]), .A2(n13), .ZN(n4) );
  NAND2_X1 U11 ( .A1(adder[14]), .A2(n11), .ZN(n5) );
  NAND2_X1 U12 ( .A1(n61), .A2(n40), .ZN(n6) );
  MUX2_X2 U13 ( .A(n21), .B(N41), .S(n233), .Z(n193) );
  NAND2_X1 U14 ( .A1(data_out_b[15]), .A2(n13), .ZN(n8) );
  NAND2_X1 U15 ( .A1(adder[15]), .A2(n11), .ZN(n9) );
  NAND2_X1 U16 ( .A1(n61), .A2(f[15]), .ZN(n10) );
  INV_X2 U17 ( .A(n39), .ZN(n61) );
  INV_X1 U18 ( .A(n14), .ZN(n13) );
  INV_X1 U19 ( .A(clear_acc), .ZN(n14) );
  NAND2_X1 U20 ( .A1(n12), .A2(N27), .ZN(n235) );
  OAI22_X1 U21 ( .A1(n177), .A2(n235), .B1(n63), .B2(n234), .ZN(n170) );
  OAI22_X1 U22 ( .A1(n178), .A2(n235), .B1(n64), .B2(n234), .ZN(n169) );
  OAI22_X1 U23 ( .A1(n179), .A2(n235), .B1(n65), .B2(n234), .ZN(n168) );
  OAI22_X1 U24 ( .A1(n180), .A2(n235), .B1(n66), .B2(n234), .ZN(n167) );
  OAI22_X1 U25 ( .A1(n181), .A2(n235), .B1(n209), .B2(n234), .ZN(n166) );
  OAI22_X1 U26 ( .A1(n182), .A2(n235), .B1(n210), .B2(n234), .ZN(n165) );
  OAI22_X1 U27 ( .A1(n183), .A2(n235), .B1(n211), .B2(n234), .ZN(n164) );
  INV_X1 U28 ( .A(n17), .ZN(n35) );
  INV_X1 U29 ( .A(wr_en_y), .ZN(n12) );
  AND2_X1 U30 ( .A1(sel[0]), .A2(sel[1]), .ZN(n16) );
  INV_X1 U31 ( .A(m_ready), .ZN(n15) );
  NAND2_X1 U32 ( .A1(m_valid), .A2(n15), .ZN(n37) );
  OAI211_X1 U33 ( .C1(sel[2]), .C2(n16), .A(sel[3]), .B(n37), .ZN(N27) );
  NAND2_X1 U34 ( .A1(clear_acc_delay), .A2(n233), .ZN(n17) );
  MUX2_X1 U35 ( .A(n18), .B(N44), .S(n35), .Z(n217) );
  MUX2_X1 U36 ( .A(n18), .B(N44), .S(n233), .Z(n196) );
  MUX2_X1 U37 ( .A(n19), .B(N43), .S(n35), .Z(n218) );
  MUX2_X1 U38 ( .A(n19), .B(N43), .S(n233), .Z(n195) );
  MUX2_X1 U39 ( .A(n20), .B(N42), .S(n35), .Z(n219) );
  MUX2_X1 U40 ( .A(n21), .B(N41), .S(n35), .Z(n220) );
  MUX2_X1 U41 ( .A(n22), .B(N40), .S(n35), .Z(n221) );
  MUX2_X1 U42 ( .A(n22), .B(N40), .S(n233), .Z(n192) );
  MUX2_X1 U43 ( .A(n23), .B(N39), .S(n35), .Z(n222) );
  MUX2_X1 U44 ( .A(n24), .B(N38), .S(n35), .Z(n223) );
  MUX2_X1 U45 ( .A(n24), .B(N38), .S(n233), .Z(n205) );
  MUX2_X1 U46 ( .A(n25), .B(N37), .S(n35), .Z(n224) );
  MUX2_X1 U47 ( .A(n26), .B(N36), .S(n35), .Z(n225) );
  MUX2_X1 U48 ( .A(n26), .B(N36), .S(n233), .Z(n203) );
  MUX2_X1 U49 ( .A(n27), .B(N35), .S(n35), .Z(n226) );
  MUX2_X1 U50 ( .A(n27), .B(N35), .S(n233), .Z(n202) );
  MUX2_X1 U51 ( .A(n28), .B(N34), .S(n35), .Z(n227) );
  MUX2_X1 U52 ( .A(n28), .B(N34), .S(n233), .Z(n201) );
  MUX2_X1 U53 ( .A(n29), .B(N33), .S(n35), .Z(n228) );
  MUX2_X1 U54 ( .A(n29), .B(N33), .S(n233), .Z(n200) );
  MUX2_X1 U55 ( .A(n32), .B(N32), .S(n35), .Z(n229) );
  MUX2_X1 U56 ( .A(n32), .B(N32), .S(n233), .Z(n199) );
  MUX2_X1 U57 ( .A(n33), .B(N31), .S(n35), .Z(n230) );
  MUX2_X1 U58 ( .A(n33), .B(N31), .S(n233), .Z(n198) );
  MUX2_X1 U59 ( .A(n34), .B(N30), .S(n35), .Z(n231) );
  MUX2_X1 U60 ( .A(n34), .B(N30), .S(n233), .Z(n197) );
  MUX2_X1 U61 ( .A(n36), .B(N29), .S(n35), .Z(n232) );
  MUX2_X1 U62 ( .A(n36), .B(N29), .S(n233), .Z(n190) );
  INV_X1 U63 ( .A(n37), .ZN(n38) );
  OAI21_X1 U64 ( .B1(n38), .B2(n7), .A(n14), .ZN(n39) );
  AOI222_X1 U65 ( .A1(data_out_b[13]), .A2(n13), .B1(adder[13]), .B2(n11), 
        .C1(n61), .C2(n41), .ZN(n42) );
  INV_X1 U66 ( .A(n42), .ZN(n73) );
  AOI222_X1 U67 ( .A1(data_out_b[12]), .A2(n13), .B1(adder[12]), .B2(n11), 
        .C1(n61), .C2(n43), .ZN(n44) );
  INV_X1 U68 ( .A(n44), .ZN(n74) );
  AOI222_X1 U69 ( .A1(data_out_b[11]), .A2(n13), .B1(adder[11]), .B2(n11), 
        .C1(n61), .C2(n45), .ZN(n46) );
  INV_X1 U70 ( .A(n46), .ZN(n75) );
  AOI222_X1 U71 ( .A1(data_out_b[10]), .A2(n13), .B1(adder[10]), .B2(n11), 
        .C1(n61), .C2(n47), .ZN(n48) );
  INV_X1 U72 ( .A(n48), .ZN(n76) );
  AOI222_X1 U73 ( .A1(data_out_b[8]), .A2(n13), .B1(adder[8]), .B2(n11), .C1(
        n61), .C2(f[8]), .ZN(n49) );
  INV_X1 U74 ( .A(n49), .ZN(n78) );
  AOI222_X1 U75 ( .A1(data_out_b[7]), .A2(n13), .B1(adder[7]), .B2(n11), .C1(
        n61), .C2(f[7]), .ZN(n50) );
  INV_X1 U76 ( .A(n50), .ZN(n79) );
  AOI222_X1 U77 ( .A1(data_out_b[6]), .A2(n13), .B1(adder[6]), .B2(n11), .C1(
        n61), .C2(f[6]), .ZN(n51) );
  INV_X1 U78 ( .A(n51), .ZN(n80) );
  AOI222_X1 U79 ( .A1(data_out_b[5]), .A2(n13), .B1(adder[5]), .B2(n11), .C1(
        n61), .C2(f[5]), .ZN(n52) );
  INV_X1 U80 ( .A(n52), .ZN(n81) );
  AOI222_X1 U81 ( .A1(data_out_b[4]), .A2(n13), .B1(adder[4]), .B2(n11), .C1(
        n61), .C2(f[4]), .ZN(n53) );
  INV_X1 U82 ( .A(n53), .ZN(n82) );
  AOI222_X1 U83 ( .A1(data_out_b[3]), .A2(n13), .B1(adder[3]), .B2(n11), .C1(
        n61), .C2(f[3]), .ZN(n54) );
  INV_X1 U84 ( .A(n54), .ZN(n83) );
  AOI222_X1 U85 ( .A1(data_out_b[2]), .A2(n13), .B1(adder[2]), .B2(n11), .C1(
        n61), .C2(n55), .ZN(n56) );
  INV_X1 U86 ( .A(n56), .ZN(n84) );
  AOI222_X1 U87 ( .A1(data_out_b[1]), .A2(n13), .B1(adder[1]), .B2(n11), .C1(
        n61), .C2(n57), .ZN(n58) );
  INV_X1 U88 ( .A(n58), .ZN(n85) );
  AOI222_X1 U89 ( .A1(data_out_b[0]), .A2(n13), .B1(adder[0]), .B2(n11), .C1(
        n61), .C2(n59), .ZN(n60) );
  INV_X1 U90 ( .A(n60), .ZN(n87) );
  AOI222_X1 U91 ( .A1(data_out_b[9]), .A2(n13), .B1(adder[9]), .B2(n11), .C1(
        n61), .C2(f[9]), .ZN(n62) );
  INV_X1 U92 ( .A(n62), .ZN(n77) );
  NOR4_X1 U93 ( .A1(n45), .A2(n43), .A3(n41), .A4(n40), .ZN(n70) );
  NOR4_X1 U94 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n47), .ZN(n69) );
  NAND4_X1 U95 ( .A1(n66), .A2(n65), .A3(n64), .A4(n63), .ZN(n67) );
  NOR4_X1 U96 ( .A1(n67), .A2(n59), .A3(n57), .A4(n55), .ZN(n68) );
  NAND3_X1 U97 ( .A1(n70), .A2(n69), .A3(n68), .ZN(n72) );
  NAND3_X1 U98 ( .A1(wr_en_y), .A2(n72), .A3(n71), .ZN(n234) );
  OAI22_X1 U99 ( .A1(n174), .A2(n235), .B1(n206), .B2(n234), .ZN(n173) );
  OAI22_X1 U100 ( .A1(n175), .A2(n235), .B1(n207), .B2(n234), .ZN(n172) );
  OAI22_X1 U101 ( .A1(n176), .A2(n235), .B1(n208), .B2(n234), .ZN(n171) );
  OAI22_X1 U102 ( .A1(n184), .A2(n235), .B1(n212), .B2(n234), .ZN(n163) );
  OAI22_X1 U103 ( .A1(n185), .A2(n235), .B1(n213), .B2(n234), .ZN(n116) );
  OAI22_X1 U104 ( .A1(n186), .A2(n235), .B1(n214), .B2(n234), .ZN(n115) );
  OAI22_X1 U105 ( .A1(n187), .A2(n235), .B1(n215), .B2(n234), .ZN(n114) );
  OAI22_X1 U106 ( .A1(n188), .A2(n235), .B1(n216), .B2(n234), .ZN(n113) );
  OAI22_X1 U107 ( .A1(n189), .A2(n235), .B1(n71), .B2(n234), .ZN(n104) );
endmodule


module layer2_12_8_12_16_ctrlpath_M12_N8_T16_P12 ( clk, reset, s_valid, 
        s_ready, m_valid, m_ready, clear_acc, wr_en_x, wr_en_y, sel, addr_x, 
        addr_w_0, addr_b_0, addr_w_1, addr_b_1, addr_w_2, addr_b_2, addr_w_3, 
        addr_b_3, addr_w_4, addr_b_4, addr_w_5, addr_b_5, addr_w_6, addr_b_6, 
        addr_w_7, addr_b_7, addr_w_8, addr_b_8, addr_w_9, addr_b_9, addr_w_10, 
        addr_b_10, addr_w_11, addr_b_11 );
  output [3:0] sel;
  output [3:0] addr_x;
  output [3:0] addr_w_0;
  output [0:0] addr_b_0;
  output [3:0] addr_w_1;
  output [0:0] addr_b_1;
  output [3:0] addr_w_2;
  output [0:0] addr_b_2;
  output [3:0] addr_w_3;
  output [0:0] addr_b_3;
  output [3:0] addr_w_4;
  output [0:0] addr_b_4;
  output [3:0] addr_w_5;
  output [0:0] addr_b_5;
  output [3:0] addr_w_6;
  output [0:0] addr_b_6;
  output [3:0] addr_w_7;
  output [0:0] addr_b_7;
  output [3:0] addr_w_8;
  output [0:0] addr_b_8;
  output [3:0] addr_w_9;
  output [0:0] addr_b_9;
  output [3:0] addr_w_10;
  output [0:0] addr_b_10;
  output [3:0] addr_w_11;
  output [0:0] addr_b_11;
  input clk, reset, s_valid, m_ready;
  output s_ready, m_valid, clear_acc, wr_en_x, wr_en_y;
  wire   n108, \state[1] , N11, clear_acc_delay, N179, N180, N181, N182, N201,
         N202, N203, N204, N223, N224, N225, N226, N245, N246, N247, N248,
         N267, N268, N269, N270, N289, N290, N291, N292, N311, N312, N313,
         N314, N333, N334, N335, N336, N355, N356, N357, N358, N377, N378,
         N379, N380, N399, N400, N401, N402, N421, N422, N423, N424, N439,
         N441, n114, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n137, n140, n144, n145, n146, n147, n148, n149, n151, n152, n153,
         n154, n156, n157, n158, n159, n161, n162, n163, n164, n166, n167,
         n168, n169, n171, n172, n173, n174, n176, n177, n178, n179, n181,
         n182, n183, n184, n186, n187, n188, n189, n191, n192, n193, n194,
         n196, n197, n198, n199, n201, n202, n203, n204, n207, n208, n209,
         n210, n212, n213, n214, n215, n216, n217, n218, n219, n221, n223,
         n224, n227, n229, n230, n231, n232, n233, n234, n235, n239, n247,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269,
         \add_1308_S2/carry[3] , \add_1308_S2/carry[2] ,
         \add_1300_S2/carry[3] , \add_1300_S2/carry[2] ,
         \add_1292_S2/carry[3] , \add_1292_S2/carry[2] ,
         \add_1284_S2/carry[3] , \add_1284_S2/carry[2] ,
         \add_1276_S2/carry[3] , \add_1276_S2/carry[2] ,
         \add_1268_S2/carry[3] , \add_1268_S2/carry[2] ,
         \add_1260_S2/carry[3] , \add_1260_S2/carry[2] ,
         \add_1252_S2/carry[3] , \add_1252_S2/carry[2] ,
         \add_1244_S2/carry[3] , \add_1244_S2/carry[2] ,
         \add_1236_S2/carry[3] , \add_1236_S2/carry[2] ,
         \add_1228_S2/carry[3] , \add_1228_S2/carry[2] ,
         \add_1220_S2/carry[3] , \add_1220_S2/carry[2] , n1, n2, n3, n5, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107;

  DFF_X1 m_valid_reg ( .D(n268), .CK(clk), .Q(m_valid), .QN(n133) );
  DFF_X1 wr_en_y_reg ( .D(n5), .CK(clk), .Q(wr_en_y) );
  DFF_X1 clear_acc_reg ( .D(N439), .CK(clk), .Q(clear_acc) );
  NAND3_X1 U205 ( .A1(addr_x[1]), .A2(n117), .A3(n214), .ZN(n213) );
  NAND3_X1 U207 ( .A1(n234), .A2(n53), .A3(wr_en_y), .ZN(n235) );
  NAND3_X1 U208 ( .A1(n232), .A2(n53), .A3(n47), .ZN(n233) );
  NAND3_X1 U210 ( .A1(addr_x[2]), .A2(addr_x[0]), .A3(addr_x[1]), .ZN(n247) );
  HA_X1 \add_1308_S2/U1_1_1  ( .A(addr_w_11[1]), .B(addr_w_11[0]), .CO(
        \add_1308_S2/carry[2] ), .S(N422) );
  HA_X1 \add_1308_S2/U1_1_2  ( .A(addr_w_11[2]), .B(\add_1308_S2/carry[2] ), 
        .CO(\add_1308_S2/carry[3] ), .S(N423) );
  HA_X1 \add_1300_S2/U1_1_1  ( .A(addr_w_10[1]), .B(addr_w_10[0]), .CO(
        \add_1300_S2/carry[2] ), .S(N400) );
  HA_X1 \add_1300_S2/U1_1_2  ( .A(addr_w_10[2]), .B(\add_1300_S2/carry[2] ), 
        .CO(\add_1300_S2/carry[3] ), .S(N401) );
  HA_X1 \add_1292_S2/U1_1_1  ( .A(addr_w_9[1]), .B(addr_w_9[0]), .CO(
        \add_1292_S2/carry[2] ), .S(N378) );
  HA_X1 \add_1292_S2/U1_1_2  ( .A(addr_w_9[2]), .B(\add_1292_S2/carry[2] ), 
        .CO(\add_1292_S2/carry[3] ), .S(N379) );
  HA_X1 \add_1284_S2/U1_1_1  ( .A(addr_w_8[1]), .B(addr_w_8[0]), .CO(
        \add_1284_S2/carry[2] ), .S(N356) );
  HA_X1 \add_1284_S2/U1_1_2  ( .A(addr_w_8[2]), .B(\add_1284_S2/carry[2] ), 
        .CO(\add_1284_S2/carry[3] ), .S(N357) );
  HA_X1 \add_1276_S2/U1_1_1  ( .A(addr_w_7[1]), .B(addr_w_7[0]), .CO(
        \add_1276_S2/carry[2] ), .S(N334) );
  HA_X1 \add_1276_S2/U1_1_2  ( .A(addr_w_7[2]), .B(\add_1276_S2/carry[2] ), 
        .CO(\add_1276_S2/carry[3] ), .S(N335) );
  HA_X1 \add_1268_S2/U1_1_1  ( .A(addr_w_6[1]), .B(addr_w_6[0]), .CO(
        \add_1268_S2/carry[2] ), .S(N312) );
  HA_X1 \add_1268_S2/U1_1_2  ( .A(addr_w_6[2]), .B(\add_1268_S2/carry[2] ), 
        .CO(\add_1268_S2/carry[3] ), .S(N313) );
  HA_X1 \add_1260_S2/U1_1_1  ( .A(addr_w_5[1]), .B(addr_w_5[0]), .CO(
        \add_1260_S2/carry[2] ), .S(N290) );
  HA_X1 \add_1260_S2/U1_1_2  ( .A(addr_w_5[2]), .B(\add_1260_S2/carry[2] ), 
        .CO(\add_1260_S2/carry[3] ), .S(N291) );
  HA_X1 \add_1252_S2/U1_1_1  ( .A(addr_w_4[1]), .B(addr_w_4[0]), .CO(
        \add_1252_S2/carry[2] ), .S(N268) );
  HA_X1 \add_1252_S2/U1_1_2  ( .A(addr_w_4[2]), .B(\add_1252_S2/carry[2] ), 
        .CO(\add_1252_S2/carry[3] ), .S(N269) );
  HA_X1 \add_1244_S2/U1_1_1  ( .A(addr_w_3[1]), .B(addr_w_3[0]), .CO(
        \add_1244_S2/carry[2] ), .S(N246) );
  HA_X1 \add_1244_S2/U1_1_2  ( .A(addr_w_3[2]), .B(\add_1244_S2/carry[2] ), 
        .CO(\add_1244_S2/carry[3] ), .S(N247) );
  HA_X1 \add_1236_S2/U1_1_1  ( .A(addr_w_2[1]), .B(addr_w_2[0]), .CO(
        \add_1236_S2/carry[2] ), .S(N224) );
  HA_X1 \add_1236_S2/U1_1_2  ( .A(addr_w_2[2]), .B(\add_1236_S2/carry[2] ), 
        .CO(\add_1236_S2/carry[3] ), .S(N225) );
  HA_X1 \add_1228_S2/U1_1_1  ( .A(addr_w_1[1]), .B(addr_w_1[0]), .CO(
        \add_1228_S2/carry[2] ), .S(N202) );
  HA_X1 \add_1228_S2/U1_1_2  ( .A(addr_w_1[2]), .B(\add_1228_S2/carry[2] ), 
        .CO(\add_1228_S2/carry[3] ), .S(N203) );
  HA_X1 \add_1220_S2/U1_1_1  ( .A(addr_w_0[1]), .B(addr_w_0[0]), .CO(
        \add_1220_S2/carry[2] ), .S(N180) );
  HA_X1 \add_1220_S2/U1_1_2  ( .A(addr_w_0[2]), .B(\add_1220_S2/carry[2] ), 
        .CO(\add_1220_S2/carry[3] ), .S(N181) );
  DFF_X1 \state_reg[2]  ( .D(n2), .CK(clk), .Q(n24), .QN(n36) );
  DFF_X1 clear_acc_delay_reg ( .D(N441), .CK(clk), .Q(clear_acc_delay), .QN(
        n132) );
  DFF_X1 \addr_b_11_reg[0]  ( .D(n258), .CK(clk), .Q(addr_b_11[0]), .QN(n131)
         );
  DFF_X1 \addr_b_10_reg[0]  ( .D(n257), .CK(clk), .Q(addr_b_10[0]), .QN(n130)
         );
  DFF_X1 \addr_b_9_reg[0]  ( .D(n256), .CK(clk), .Q(addr_b_9[0]), .QN(n129) );
  DFF_X1 \addr_b_8_reg[0]  ( .D(n255), .CK(clk), .Q(addr_b_8[0]), .QN(n128) );
  DFF_X1 \addr_b_7_reg[0]  ( .D(n254), .CK(clk), .Q(addr_b_7[0]), .QN(n127) );
  DFF_X1 \addr_b_6_reg[0]  ( .D(n253), .CK(clk), .Q(addr_b_6[0]), .QN(n126) );
  DFF_X1 \addr_b_5_reg[0]  ( .D(n252), .CK(clk), .Q(addr_b_5[0]), .QN(n125) );
  DFF_X1 \addr_b_4_reg[0]  ( .D(n251), .CK(clk), .Q(addr_b_4[0]), .QN(n124) );
  DFF_X1 \addr_b_3_reg[0]  ( .D(n262), .CK(clk), .Q(addr_b_3[0]), .QN(n123) );
  DFF_X1 \addr_b_2_reg[0]  ( .D(n261), .CK(clk), .Q(addr_b_2[0]), .QN(n122) );
  DFF_X1 \addr_b_1_reg[0]  ( .D(n260), .CK(clk), .Q(addr_b_1[0]), .QN(n121) );
  DFF_X1 \addr_b_0_reg[0]  ( .D(n259), .CK(clk), .Q(addr_b_0[0]), .QN(n120) );
  DFF_X1 \sel_count_reg[0]  ( .D(n269), .CK(clk), .Q(sel[0]), .QN(n137) );
  DFF_X1 \state_reg[1]  ( .D(n48), .CK(clk), .Q(\state[1] ), .QN(n114) );
  DFF_X1 \state_reg[0]  ( .D(N11), .CK(clk), .Q(n32), .QN(n35) );
  DFF_X1 \sel_count_reg[1]  ( .D(n57), .CK(clk), .Q(sel[1]), .QN(n17) );
  DFF_X1 \sel_count_reg[3]  ( .D(n267), .CK(clk), .Q(sel[3]), .QN(n134) );
  DFF_X1 \sel_count_reg[2]  ( .D(n266), .CK(clk), .Q(sel[2]), .QN(n135) );
  DFF_X1 \addr_x_reg[0]  ( .D(n264), .CK(clk), .Q(addr_x[0]), .QN(n119) );
  DFF_X1 \addr_w2_11_reg[2]  ( .D(n100), .CK(clk), .Q(addr_w_11[2]) );
  DFF_X1 \addr_w2_11_reg[1]  ( .D(n99), .CK(clk), .Q(addr_w_11[1]) );
  DFF_X1 \addr_w2_10_reg[3]  ( .D(n97), .CK(clk), .Q(addr_w_10[3]) );
  DFF_X1 \addr_w2_10_reg[2]  ( .D(n96), .CK(clk), .Q(addr_w_10[2]) );
  DFF_X1 \addr_w2_10_reg[1]  ( .D(n95), .CK(clk), .Q(addr_w_10[1]) );
  DFF_X1 \addr_w2_10_reg[0]  ( .D(n94), .CK(clk), .Q(addr_w_10[0]), .QN(N399)
         );
  DFF_X1 \addr_w2_9_reg[3]  ( .D(n105), .CK(clk), .Q(addr_w_9[3]) );
  DFF_X1 \addr_w2_8_reg[2]  ( .D(n92), .CK(clk), .Q(addr_w_8[2]) );
  DFF_X1 \addr_w2_8_reg[1]  ( .D(n91), .CK(clk), .Q(addr_w_8[1]) );
  DFF_X1 \addr_w2_7_reg[0]  ( .D(n86), .CK(clk), .Q(addr_w_7[0]), .QN(N333) );
  DFF_X1 \addr_w2_6_reg[2]  ( .D(n84), .CK(clk), .Q(addr_w_6[2]) );
  DFF_X1 \addr_w2_6_reg[1]  ( .D(n83), .CK(clk), .Q(addr_w_6[1]) );
  DFF_X1 \addr_w2_5_reg[2]  ( .D(n80), .CK(clk), .Q(addr_w_5[2]) );
  DFF_X1 \addr_w2_5_reg[1]  ( .D(n79), .CK(clk), .Q(addr_w_5[1]) );
  DFF_X1 \addr_w2_5_reg[0]  ( .D(n78), .CK(clk), .Q(addr_w_5[0]), .QN(N289) );
  DFF_X1 \addr_w2_4_reg[3]  ( .D(n77), .CK(clk), .Q(addr_w_4[3]) );
  DFF_X1 \addr_w2_4_reg[2]  ( .D(n76), .CK(clk), .Q(addr_w_4[2]) );
  DFF_X1 \addr_w2_3_reg[3]  ( .D(n73), .CK(clk), .Q(addr_w_3[3]) );
  DFF_X1 \addr_w2_3_reg[2]  ( .D(n72), .CK(clk), .Q(addr_w_3[2]) );
  DFF_X1 \addr_w2_3_reg[1]  ( .D(n71), .CK(clk), .Q(addr_w_3[1]) );
  DFF_X1 \addr_w2_2_reg[1]  ( .D(n67), .CK(clk), .Q(addr_w_2[1]) );
  DFF_X1 \addr_w2_2_reg[0]  ( .D(n66), .CK(clk), .Q(addr_w_2[0]), .QN(N223) );
  DFF_X1 \addr_w2_1_reg[3]  ( .D(n65), .CK(clk), .Q(addr_w_1[3]) );
  DFF_X1 \addr_w2_1_reg[2]  ( .D(n64), .CK(clk), .Q(addr_w_1[2]) );
  DFF_X1 \addr_w2_1_reg[0]  ( .D(n62), .CK(clk), .Q(addr_w_1[0]), .QN(N201) );
  DFF_X1 \addr_w2_0_reg[3]  ( .D(n61), .CK(clk), .Q(addr_w_0[3]) );
  DFF_X1 \addr_w2_0_reg[1]  ( .D(n59), .CK(clk), .Q(addr_w_0[1]) );
  DFF_X1 \addr_w2_8_reg[3]  ( .D(n93), .CK(clk), .Q(addr_w_8[3]) );
  DFF_X1 \addr_w2_5_reg[3]  ( .D(n81), .CK(clk), .Q(addr_w_5[3]) );
  DFF_X1 \addr_w2_7_reg[2]  ( .D(n88), .CK(clk), .Q(addr_w_7[2]) );
  DFF_X1 \addr_w2_11_reg[3]  ( .D(n101), .CK(clk), .Q(addr_w_11[3]) );
  DFF_X1 \addr_w2_1_reg[1]  ( .D(n63), .CK(clk), .Q(addr_w_1[1]) );
  DFF_X1 \addr_w2_2_reg[2]  ( .D(n68), .CK(clk), .Q(addr_w_2[2]) );
  DFF_X1 \addr_w2_9_reg[0]  ( .D(n102), .CK(clk), .Q(addr_w_9[0]), .QN(N377)
         );
  DFF_X1 \addr_w2_9_reg[1]  ( .D(n103), .CK(clk), .Q(addr_w_9[1]) );
  DFF_X1 \addr_w2_4_reg[1]  ( .D(n75), .CK(clk), .Q(addr_w_4[1]) );
  DFF_X1 \addr_w2_9_reg[2]  ( .D(n104), .CK(clk), .Q(addr_w_9[2]) );
  DFF_X1 \addr_w2_0_reg[2]  ( .D(n60), .CK(clk), .Q(addr_w_0[2]) );
  DFF_X1 \addr_w2_7_reg[1]  ( .D(n87), .CK(clk), .Q(addr_w_7[1]) );
  DFF_X1 \addr_w2_11_reg[0]  ( .D(n98), .CK(clk), .Q(addr_w_11[0]), .QN(N421)
         );
  DFF_X1 \addr_w2_8_reg[0]  ( .D(n90), .CK(clk), .Q(addr_w_8[0]), .QN(N355) );
  DFF_X1 \addr_w2_6_reg[0]  ( .D(n82), .CK(clk), .Q(addr_w_6[0]), .QN(N311) );
  DFF_X1 \addr_w2_3_reg[0]  ( .D(n70), .CK(clk), .Q(addr_w_3[0]), .QN(N245) );
  DFF_X1 \addr_w2_7_reg[3]  ( .D(n89), .CK(clk), .Q(addr_w_7[3]) );
  DFF_X1 \addr_w2_6_reg[3]  ( .D(n85), .CK(clk), .Q(addr_w_6[3]) );
  DFF_X1 \addr_w2_4_reg[0]  ( .D(n74), .CK(clk), .Q(addr_w_4[0]), .QN(N267) );
  DFF_X1 \addr_w2_2_reg[3]  ( .D(n69), .CK(clk), .Q(addr_w_2[3]) );
  DFF_X1 \addr_w2_0_reg[0]  ( .D(n58), .CK(clk), .Q(addr_w_0[0]), .QN(N179) );
  DFF_X1 \addr_x_reg[1]  ( .D(n56), .CK(clk), .Q(addr_x[1]), .QN(n118) );
  DFF_X1 \addr_x_reg[2]  ( .D(n263), .CK(clk), .Q(addr_x[2]), .QN(n117) );
  DFF_X1 \addr_x_reg[3]  ( .D(n265), .CK(clk), .Q(addr_x[3]), .QN(n116) );
  BUF_X1 U3 ( .A(n145), .Z(n15) );
  BUF_X1 U4 ( .A(n145), .Z(n14) );
  NOR2_X1 U5 ( .A1(reset), .A2(n1), .ZN(n2) );
  INV_X1 U6 ( .A(n140), .ZN(n1) );
  CLKBUF_X1 U7 ( .A(n41), .Z(n3) );
  CLKBUF_X3 U8 ( .A(n108), .Z(s_ready) );
  OAI22_X1 U9 ( .A1(reset), .A2(n42), .B1(n41), .B2(n140), .ZN(n108) );
  BUF_X1 U10 ( .A(n9), .Z(n10) );
  BUF_X1 U11 ( .A(n9), .Z(n11) );
  BUF_X1 U12 ( .A(n9), .Z(n13) );
  BUF_X1 U13 ( .A(n9), .Z(n12) );
  OAI21_X1 U14 ( .B1(n208), .B2(wr_en_x), .A(n53), .ZN(n218) );
  NOR3_X1 U15 ( .A1(n223), .A2(n224), .A3(n107), .ZN(n208) );
  NAND4_X1 U16 ( .A1(n221), .A2(n106), .A3(n218), .A4(n53), .ZN(n217) );
  NOR2_X1 U17 ( .A1(n239), .A2(n207), .ZN(n221) );
  AND2_X1 U18 ( .A1(n208), .A2(n53), .ZN(n145) );
  AND2_X1 U19 ( .A1(n8), .A2(n32), .ZN(n5) );
  BUF_X1 U20 ( .A(n146), .Z(n9) );
  NAND2_X1 U21 ( .A1(n221), .A2(n53), .ZN(N439) );
  INV_X1 U22 ( .A(n212), .ZN(n54) );
  NAND2_X1 U23 ( .A1(clear_acc_delay), .A2(n53), .ZN(n210) );
  NOR4_X1 U24 ( .A1(n49), .A2(n207), .A3(n145), .A4(reset), .ZN(n146) );
  NAND4_X1 U25 ( .A1(n47), .A2(m_valid), .A3(m_ready), .A4(n53), .ZN(n232) );
  OAI22_X1 U26 ( .A1(n209), .A2(n123), .B1(addr_b_3[0]), .B2(n210), .ZN(n262)
         );
  OAI22_X1 U27 ( .A1(n209), .A2(n122), .B1(addr_b_2[0]), .B2(n210), .ZN(n261)
         );
  OAI22_X1 U28 ( .A1(n209), .A2(n121), .B1(addr_b_1[0]), .B2(n210), .ZN(n260)
         );
  OAI22_X1 U29 ( .A1(n209), .A2(n120), .B1(addr_b_0[0]), .B2(n210), .ZN(n259)
         );
  OAI22_X1 U30 ( .A1(n209), .A2(n131), .B1(addr_b_11[0]), .B2(n210), .ZN(n258)
         );
  OAI22_X1 U31 ( .A1(n209), .A2(n130), .B1(addr_b_10[0]), .B2(n210), .ZN(n257)
         );
  OAI22_X1 U32 ( .A1(n209), .A2(n129), .B1(addr_b_9[0]), .B2(n210), .ZN(n256)
         );
  OAI22_X1 U33 ( .A1(n209), .A2(n128), .B1(addr_b_8[0]), .B2(n210), .ZN(n255)
         );
  OAI22_X1 U34 ( .A1(n209), .A2(n127), .B1(addr_b_7[0]), .B2(n210), .ZN(n254)
         );
  OAI22_X1 U35 ( .A1(n209), .A2(n126), .B1(addr_b_6[0]), .B2(n210), .ZN(n253)
         );
  OAI22_X1 U36 ( .A1(n209), .A2(n125), .B1(addr_b_5[0]), .B2(n210), .ZN(n252)
         );
  OAI22_X1 U37 ( .A1(n209), .A2(n124), .B1(addr_b_4[0]), .B2(n210), .ZN(n251)
         );
  AOI21_X1 U38 ( .B1(sel[3]), .B2(sel[2]), .A(n7), .ZN(n224) );
  AOI21_X1 U39 ( .B1(n118), .B2(n55), .A(n216), .ZN(n212) );
  NOR2_X1 U40 ( .A1(n232), .A2(n137), .ZN(n227) );
  OAI21_X1 U41 ( .B1(addr_x[0]), .B2(n218), .A(n217), .ZN(n216) );
  NOR2_X1 U42 ( .A1(n218), .A2(n119), .ZN(n214) );
  NOR2_X1 U43 ( .A1(n133), .A2(m_ready), .ZN(n223) );
  INV_X1 U44 ( .A(n204), .ZN(n58) );
  AOI22_X1 U45 ( .A1(N179), .A2(n14), .B1(addr_w_0[0]), .B2(n10), .ZN(n204) );
  OAI22_X1 U46 ( .A1(n119), .A2(n217), .B1(addr_x[0]), .B2(n218), .ZN(n264) );
  INV_X1 U47 ( .A(n189), .ZN(n70) );
  AOI22_X1 U48 ( .A1(N245), .A2(n14), .B1(addr_w_3[0]), .B2(n11), .ZN(n189) );
  INV_X1 U49 ( .A(n171), .ZN(n85) );
  AOI22_X1 U50 ( .A1(N314), .A2(n15), .B1(addr_w_6[3]), .B2(n12), .ZN(n171) );
  XOR2_X1 U51 ( .A(addr_w_6[3]), .B(\add_1268_S2/carry[3] ), .Z(N314) );
  INV_X1 U52 ( .A(n166), .ZN(n89) );
  AOI22_X1 U53 ( .A1(N336), .A2(n15), .B1(addr_w_7[3]), .B2(n12), .ZN(n166) );
  XOR2_X1 U54 ( .A(addr_w_7[3]), .B(\add_1276_S2/carry[3] ), .Z(N336) );
  INV_X1 U55 ( .A(n174), .ZN(n82) );
  AOI22_X1 U56 ( .A1(N311), .A2(n15), .B1(addr_w_6[0]), .B2(n12), .ZN(n174) );
  INV_X1 U57 ( .A(n149), .ZN(n102) );
  AOI22_X1 U58 ( .A1(N377), .A2(n15), .B1(addr_w_9[0]), .B2(n13), .ZN(n149) );
  INV_X1 U59 ( .A(n192), .ZN(n68) );
  AOI22_X1 U60 ( .A1(N225), .A2(n14), .B1(addr_w_2[2]), .B2(n10), .ZN(n192) );
  INV_X1 U61 ( .A(n147), .ZN(n104) );
  AOI22_X1 U62 ( .A1(N379), .A2(n15), .B1(addr_w_9[2]), .B2(n13), .ZN(n147) );
  INV_X1 U63 ( .A(n203), .ZN(n59) );
  AOI22_X1 U64 ( .A1(N180), .A2(n14), .B1(addr_w_0[1]), .B2(n10), .ZN(n203) );
  INV_X1 U65 ( .A(n153), .ZN(n99) );
  AOI22_X1 U66 ( .A1(N422), .A2(n14), .B1(addr_w_11[1]), .B2(n13), .ZN(n153)
         );
  INV_X1 U67 ( .A(n177), .ZN(n80) );
  AOI22_X1 U68 ( .A1(N291), .A2(n14), .B1(addr_w_5[2]), .B2(n11), .ZN(n177) );
  INV_X1 U69 ( .A(n201), .ZN(n61) );
  AOI22_X1 U70 ( .A1(N182), .A2(n14), .B1(addr_w_0[3]), .B2(n10), .ZN(n201) );
  XOR2_X1 U71 ( .A(addr_w_0[3]), .B(\add_1220_S2/carry[3] ), .Z(N182) );
  INV_X1 U72 ( .A(n186), .ZN(n73) );
  AOI22_X1 U73 ( .A1(N248), .A2(n14), .B1(addr_w_3[3]), .B2(n11), .ZN(n186) );
  XOR2_X1 U74 ( .A(addr_w_3[3]), .B(\add_1244_S2/carry[3] ), .Z(N248) );
  INV_X1 U75 ( .A(n181), .ZN(n77) );
  AOI22_X1 U76 ( .A1(N270), .A2(n14), .B1(addr_w_4[3]), .B2(n11), .ZN(n181) );
  XOR2_X1 U77 ( .A(addr_w_4[3]), .B(\add_1252_S2/carry[3] ), .Z(N270) );
  INV_X1 U78 ( .A(n196), .ZN(n65) );
  AOI22_X1 U79 ( .A1(N204), .A2(n14), .B1(addr_w_1[3]), .B2(n10), .ZN(n196) );
  XOR2_X1 U80 ( .A(addr_w_1[3]), .B(\add_1228_S2/carry[3] ), .Z(N204) );
  INV_X1 U81 ( .A(n197), .ZN(n64) );
  AOI22_X1 U82 ( .A1(N203), .A2(n14), .B1(addr_w_1[2]), .B2(n10), .ZN(n197) );
  INV_X1 U83 ( .A(n215), .ZN(n56) );
  AOI22_X1 U84 ( .A1(n216), .A2(addr_x[1]), .B1(n118), .B2(n214), .ZN(n215) );
  NAND4_X1 U85 ( .A1(n227), .A2(sel[2]), .A3(sel[1]), .A4(n134), .ZN(n231) );
  AOI21_X1 U86 ( .B1(n52), .B2(n135), .A(n19), .ZN(n230) );
  AND3_X1 U87 ( .A1(s_valid), .A2(n1), .A3(n40), .ZN(wr_en_x) );
  OAI21_X1 U88 ( .B1(n224), .B2(n223), .A(n53), .ZN(n234) );
  AOI21_X1 U89 ( .B1(n55), .B2(n117), .A(n54), .ZN(n219) );
  AND3_X1 U90 ( .A1(sel[0]), .A2(sel[3]), .A3(sel[1]), .ZN(n7) );
  OAI21_X1 U91 ( .B1(n212), .B2(n117), .A(n213), .ZN(n263) );
  OAI21_X1 U92 ( .B1(sel[0]), .B2(n232), .A(n233), .ZN(n229) );
  AND2_X1 U93 ( .A1(n114), .A2(n24), .ZN(n8) );
  INV_X1 U94 ( .A(n202), .ZN(n60) );
  AOI22_X1 U95 ( .A1(N181), .A2(n14), .B1(addr_w_0[2]), .B2(n10), .ZN(n202) );
  INV_X1 U96 ( .A(n191), .ZN(n69) );
  AOI22_X1 U97 ( .A1(N226), .A2(n14), .B1(addr_w_2[3]), .B2(n10), .ZN(n191) );
  XOR2_X1 U98 ( .A(addr_w_2[3]), .B(\add_1236_S2/carry[3] ), .Z(N226) );
  INV_X1 U99 ( .A(n184), .ZN(n74) );
  AOI22_X1 U100 ( .A1(N267), .A2(n14), .B1(addr_w_4[0]), .B2(n11), .ZN(n184)
         );
  INV_X1 U101 ( .A(n154), .ZN(n98) );
  AOI22_X1 U102 ( .A1(N421), .A2(n15), .B1(addr_w_11[0]), .B2(n13), .ZN(n154)
         );
  INV_X1 U103 ( .A(n168), .ZN(n87) );
  AOI22_X1 U104 ( .A1(N334), .A2(n15), .B1(addr_w_7[1]), .B2(n12), .ZN(n168)
         );
  INV_X1 U105 ( .A(n164), .ZN(n90) );
  AOI22_X1 U106 ( .A1(N355), .A2(n15), .B1(addr_w_8[0]), .B2(n12), .ZN(n164)
         );
  INV_X1 U107 ( .A(n183), .ZN(n75) );
  AOI22_X1 U108 ( .A1(N268), .A2(n14), .B1(addr_w_4[1]), .B2(n11), .ZN(n183)
         );
  INV_X1 U109 ( .A(n151), .ZN(n101) );
  AOI22_X1 U110 ( .A1(N424), .A2(n15), .B1(addr_w_11[3]), .B2(n13), .ZN(n151)
         );
  XOR2_X1 U111 ( .A(addr_w_11[3]), .B(\add_1308_S2/carry[3] ), .Z(N424) );
  INV_X1 U112 ( .A(n148), .ZN(n103) );
  AOI22_X1 U113 ( .A1(N378), .A2(n15), .B1(addr_w_9[1]), .B2(n13), .ZN(n148)
         );
  INV_X1 U114 ( .A(n176), .ZN(n81) );
  AOI22_X1 U115 ( .A1(N292), .A2(n15), .B1(addr_w_5[3]), .B2(n11), .ZN(n176)
         );
  XOR2_X1 U116 ( .A(addr_w_5[3]), .B(\add_1260_S2/carry[3] ), .Z(N292) );
  INV_X1 U117 ( .A(n161), .ZN(n93) );
  AOI22_X1 U118 ( .A1(N358), .A2(n15), .B1(addr_w_8[3]), .B2(n12), .ZN(n161)
         );
  XOR2_X1 U119 ( .A(addr_w_8[3]), .B(\add_1284_S2/carry[3] ), .Z(N358) );
  INV_X1 U120 ( .A(n167), .ZN(n88) );
  AOI22_X1 U121 ( .A1(N335), .A2(n15), .B1(addr_w_7[2]), .B2(n12), .ZN(n167)
         );
  INV_X1 U122 ( .A(n193), .ZN(n67) );
  AOI22_X1 U123 ( .A1(N224), .A2(n14), .B1(addr_w_2[1]), .B2(n10), .ZN(n193)
         );
  INV_X1 U124 ( .A(n194), .ZN(n66) );
  AOI22_X1 U125 ( .A1(N223), .A2(n14), .B1(addr_w_2[0]), .B2(n10), .ZN(n194)
         );
  INV_X1 U126 ( .A(n144), .ZN(n105) );
  AOI22_X1 U127 ( .A1(N380), .A2(n14), .B1(addr_w_9[3]), .B2(n13), .ZN(n144)
         );
  XOR2_X1 U128 ( .A(addr_w_9[3]), .B(\add_1292_S2/carry[3] ), .Z(N380) );
  INV_X1 U129 ( .A(n198), .ZN(n63) );
  AOI22_X1 U130 ( .A1(N202), .A2(n14), .B1(addr_w_1[1]), .B2(n10), .ZN(n198)
         );
  INV_X1 U131 ( .A(n169), .ZN(n86) );
  AOI22_X1 U132 ( .A1(N333), .A2(n15), .B1(addr_w_7[0]), .B2(n12), .ZN(n169)
         );
  INV_X1 U133 ( .A(n156), .ZN(n97) );
  AOI22_X1 U134 ( .A1(N402), .A2(n15), .B1(addr_w_10[3]), .B2(n13), .ZN(n156)
         );
  XOR2_X1 U135 ( .A(addr_w_10[3]), .B(\add_1300_S2/carry[3] ), .Z(N402) );
  INV_X1 U136 ( .A(n158), .ZN(n95) );
  AOI22_X1 U137 ( .A1(N400), .A2(n15), .B1(addr_w_10[1]), .B2(n13), .ZN(n158)
         );
  INV_X1 U138 ( .A(n163), .ZN(n91) );
  AOI22_X1 U139 ( .A1(N356), .A2(n15), .B1(addr_w_8[1]), .B2(n12), .ZN(n163)
         );
  INV_X1 U140 ( .A(n199), .ZN(n62) );
  AOI22_X1 U141 ( .A1(N201), .A2(n14), .B1(addr_w_1[0]), .B2(n10), .ZN(n199)
         );
  INV_X1 U142 ( .A(n179), .ZN(n78) );
  AOI22_X1 U143 ( .A1(N289), .A2(n14), .B1(addr_w_5[0]), .B2(n11), .ZN(n179)
         );
  INV_X1 U144 ( .A(n157), .ZN(n96) );
  AOI22_X1 U145 ( .A1(N401), .A2(n15), .B1(addr_w_10[2]), .B2(n13), .ZN(n157)
         );
  INV_X1 U146 ( .A(n173), .ZN(n83) );
  AOI22_X1 U147 ( .A1(N312), .A2(n15), .B1(addr_w_6[1]), .B2(n12), .ZN(n173)
         );
  INV_X1 U148 ( .A(n178), .ZN(n79) );
  AOI22_X1 U149 ( .A1(N290), .A2(n14), .B1(addr_w_5[1]), .B2(n11), .ZN(n178)
         );
  INV_X1 U150 ( .A(n162), .ZN(n92) );
  AOI22_X1 U151 ( .A1(N357), .A2(n15), .B1(addr_w_8[2]), .B2(n12), .ZN(n162)
         );
  INV_X1 U152 ( .A(n159), .ZN(n94) );
  AOI22_X1 U153 ( .A1(N399), .A2(n15), .B1(addr_w_10[0]), .B2(n13), .ZN(n159)
         );
  INV_X1 U154 ( .A(n152), .ZN(n100) );
  AOI22_X1 U155 ( .A1(N423), .A2(n15), .B1(addr_w_11[2]), .B2(n13), .ZN(n152)
         );
  INV_X1 U156 ( .A(n187), .ZN(n72) );
  AOI22_X1 U157 ( .A1(N247), .A2(n14), .B1(addr_w_3[2]), .B2(n11), .ZN(n187)
         );
  INV_X1 U158 ( .A(n188), .ZN(n71) );
  AOI22_X1 U159 ( .A1(N246), .A2(n14), .B1(addr_w_3[1]), .B2(n11), .ZN(n188)
         );
  INV_X1 U160 ( .A(n182), .ZN(n76) );
  AOI22_X1 U161 ( .A1(N269), .A2(n14), .B1(addr_w_4[2]), .B2(n11), .ZN(n182)
         );
  INV_X1 U162 ( .A(n172), .ZN(n84) );
  AOI22_X1 U163 ( .A1(N313), .A2(n15), .B1(addr_w_6[2]), .B2(n12), .ZN(n172)
         );
  AND2_X1 U164 ( .A1(clear_acc), .A2(n50), .ZN(N441) );
  INV_X1 U165 ( .A(reset), .ZN(n53) );
  INV_X1 U166 ( .A(n229), .ZN(n18) );
  INV_X1 U167 ( .A(n227), .ZN(n16) );
  OAI22_X1 U168 ( .A1(n17), .A2(n18), .B1(sel[1]), .B2(n16), .ZN(n57) );
  OAI21_X1 U169 ( .B1(n232), .B2(sel[1]), .A(n18), .ZN(n19) );
  INV_X1 U170 ( .A(n19), .ZN(n51) );
  NAND3_X1 U171 ( .A1(addr_x[2]), .A2(addr_x[1]), .A3(n214), .ZN(n20) );
  MUX2_X1 U172 ( .A(n219), .B(n20), .S(n116), .Z(n21) );
  INV_X1 U173 ( .A(n21), .ZN(n265) );
  OAI22_X1 U174 ( .A1(n137), .A2(n233), .B1(sel[0]), .B2(n232), .ZN(n269) );
  NAND2_X1 U175 ( .A1(n227), .A2(sel[1]), .ZN(n22) );
  MUX2_X1 U176 ( .A(n51), .B(n22), .S(n135), .Z(n23) );
  NAND2_X1 U177 ( .A1(n53), .A2(n23), .ZN(n266) );
  OAI211_X1 U178 ( .C1(n230), .C2(n134), .A(n231), .B(n53), .ZN(n267) );
  NAND2_X1 U179 ( .A1(n8), .A2(n35), .ZN(n107) );
  AND2_X1 U180 ( .A1(n247), .A2(n116), .ZN(n30) );
  NAND3_X1 U181 ( .A1(\state[1] ), .A2(n35), .A3(n24), .ZN(n37) );
  NAND4_X1 U182 ( .A1(m_valid), .A2(n135), .A3(m_ready), .A4(n7), .ZN(n25) );
  NAND2_X1 U183 ( .A1(\state[1] ), .A2(n32), .ZN(n46) );
  INV_X1 U184 ( .A(n46), .ZN(n34) );
  NAND2_X1 U185 ( .A1(n34), .A2(n24), .ZN(n106) );
  INV_X1 U186 ( .A(n106), .ZN(n49) );
  NAND2_X1 U187 ( .A1(n25), .A2(n49), .ZN(n39) );
  NOR2_X1 U188 ( .A1(addr_x[3]), .A2(n46), .ZN(n27) );
  NAND3_X1 U189 ( .A1(n36), .A2(n114), .A3(n35), .ZN(n42) );
  INV_X1 U190 ( .A(n42), .ZN(n26) );
  AOI22_X1 U191 ( .A1(n27), .A2(n36), .B1(s_valid), .B2(n26), .ZN(n28) );
  NAND3_X1 U192 ( .A1(n37), .A2(n39), .A3(n28), .ZN(n33) );
  INV_X1 U193 ( .A(n33), .ZN(n29) );
  OAI21_X1 U194 ( .B1(n107), .B2(n30), .A(n29), .ZN(n40) );
  INV_X1 U195 ( .A(n40), .ZN(n31) );
  NOR2_X1 U196 ( .A1(reset), .A2(n31), .ZN(N11) );
  OAI21_X1 U197 ( .B1(n133), .B2(n234), .A(n235), .ZN(n268) );
  OAI21_X1 U198 ( .B1(n5), .B2(n33), .A(n53), .ZN(n41) );
  INV_X1 U199 ( .A(n3), .ZN(n48) );
  NAND3_X1 U200 ( .A1(n34), .A2(n36), .A3(addr_x[3]), .ZN(n45) );
  INV_X1 U201 ( .A(n107), .ZN(n50) );
  NAND3_X1 U202 ( .A1(\state[1] ), .A2(n36), .A3(n35), .ZN(n44) );
  NAND2_X1 U203 ( .A1(n44), .A2(n37), .ZN(n43) );
  NOR3_X1 U204 ( .A1(n5), .A2(n50), .A3(n43), .ZN(n38) );
  NAND3_X1 U206 ( .A1(n39), .A2(n45), .A3(n38), .ZN(n140) );
  INV_X1 U209 ( .A(n43), .ZN(n47) );
  INV_X1 U211 ( .A(n44), .ZN(n239) );
  INV_X1 U212 ( .A(n45), .ZN(n207) );
  INV_X1 U213 ( .A(n232), .ZN(n52) );
  INV_X1 U214 ( .A(n218), .ZN(n55) );
  NAND3_X1 U215 ( .A1(n132), .A2(n53), .A3(n46), .ZN(n209) );
endmodule


module layer2_12_8_12_16 ( clk, reset, s_valid, m_ready, data_in, m_valid, 
        s_ready, data_out );
  input [15:0] data_in;
  output [15:0] data_out;
  input clk, reset, s_valid, m_ready;
  output m_valid, s_ready;
  wire   wr_en_x, \addr_b_0[0] , \addr_b_1[0] , \addr_b_2[0] , \addr_b_3[0] ,
         \addr_b_4[0] , \addr_b_5[0] , \addr_b_6[0] , \addr_b_7[0] ,
         \addr_b_8[0] , \addr_b_9[0] , \addr_b_10[0] , \addr_b_11[0] ,
         clear_acc, wr_en_y, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n1, n2, n3, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124;
  wire   [15:0] data_out_x;
  wire   [3:0] addr_x;
  wire   [3:0] addr_w_0;
  wire   [15:0] data_out_w_0;
  wire   [15:0] data_out_b_0;
  wire   [3:0] addr_w_1;
  wire   [15:0] data_out_w_1;
  wire   [15:0] data_out_b_1;
  wire   [3:0] addr_w_2;
  wire   [15:0] data_out_w_2;
  wire   [15:0] data_out_b_2;
  wire   [3:0] addr_w_3;
  wire   [15:0] data_out_w_3;
  wire   [15:0] data_out_b_3;
  wire   [3:0] addr_w_4;
  wire   [15:0] data_out_w_4;
  wire   [15:0] data_out_b_4;
  wire   [3:0] addr_w_5;
  wire   [15:0] data_out_w_5;
  wire   [15:0] data_out_b_5;
  wire   [3:0] addr_w_6;
  wire   [15:0] data_out_w_6;
  wire   [15:0] data_out_b_6;
  wire   [3:0] addr_w_7;
  wire   [15:0] data_out_w_7;
  wire   [15:0] data_out_b_7;
  wire   [3:0] addr_w_8;
  wire   [15:0] data_out_w_8;
  wire   [15:0] data_out_b_8;
  wire   [3:0] addr_w_9;
  wire   [15:0] data_out_w_9;
  wire   [15:0] data_out_b_9;
  wire   [3:0] addr_w_10;
  wire   [15:0] data_out_w_10;
  wire   [15:0] data_out_b_10;
  wire   [3:0] addr_w_11;
  wire   [15:0] data_out_w_11;
  wire   [15:0] data_out_b_11;
  wire   [15:0] data_out_0;
  wire   [3:0] sel;
  wire   [15:0] data_out_1;
  wire   [15:0] data_out_2;
  wire   [15:0] data_out_3;
  wire   [15:0] data_out_4;
  wire   [15:0] data_out_5;
  wire   [15:0] data_out_6;
  wire   [15:0] data_out_7;
  wire   [15:0] data_out_8;
  wire   [15:0] data_out_9;
  wire   [15:0] data_out_10;
  wire   [15:0] data_out_11;
  wire   SYNOPSYS_UNCONNECTED__0;

  AND3_X2 U83 ( .A1(n83), .A2(sel[1]), .A3(sel[2]), .ZN(n13) );
  AND3_X2 U85 ( .A1(sel[2]), .A2(sel[1]), .A3(n84), .ZN(n11) );
  AND3_X2 U87 ( .A1(sel[2]), .A2(n123), .A3(n84), .ZN(n16) );
  memory_WIDTH16_SIZE8_LOGSIZE4 mem_x ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_x), .addr(addr_x), .wr_en(wr_en_x) );
  layer2_12_8_12_16_W_rom_0 mem_w_0 ( .clk(clk), .addr(addr_w_0), .z(
        data_out_w_0) );
  layer2_12_8_12_16_B_rom_0 mem_b_0 ( .clk(clk), .addr(\addr_b_0[0] ) );
  layer2_12_8_12_16_W_rom_1 mem_w_1 ( .clk(clk), .addr(addr_w_1), .z(
        data_out_w_1) );
  layer2_12_8_12_16_B_rom_1 mem_b_1 ( .clk(clk), .addr(\addr_b_1[0] ) );
  layer2_12_8_12_16_W_rom_2 mem_w_2 ( .clk(clk), .addr(addr_w_2), .z(
        data_out_w_2) );
  layer2_12_8_12_16_B_rom_2 mem_b_2 ( .clk(clk), .addr(\addr_b_2[0] ) );
  layer2_12_8_12_16_W_rom_3 mem_w_3 ( .clk(clk), .addr(addr_w_3), .z(
        data_out_w_3) );
  layer2_12_8_12_16_B_rom_3 mem_b_3 ( .clk(clk), .addr(\addr_b_3[0] ) );
  layer2_12_8_12_16_W_rom_4 mem_w_4 ( .clk(clk), .addr(addr_w_4), .z(
        data_out_w_4) );
  layer2_12_8_12_16_B_rom_4 mem_b_4 ( .clk(clk), .addr(\addr_b_4[0] ) );
  layer2_12_8_12_16_W_rom_5 mem_w_5 ( .clk(clk), .addr(addr_w_5), .z(
        data_out_w_5) );
  layer2_12_8_12_16_B_rom_5 mem_b_5 ( .clk(clk), .addr(\addr_b_5[0] ) );
  layer2_12_8_12_16_W_rom_6 mem_w_6 ( .clk(clk), .addr(addr_w_6), .z(
        data_out_w_6) );
  layer2_12_8_12_16_B_rom_6 mem_b_6 ( .clk(clk), .addr(\addr_b_6[0] ) );
  layer2_12_8_12_16_W_rom_7 mem_w_7 ( .clk(clk), .addr(addr_w_7), .z(
        data_out_w_7) );
  layer2_12_8_12_16_B_rom_7 mem_b_7 ( .clk(clk), .addr(\addr_b_7[0] ) );
  layer2_12_8_12_16_W_rom_8 mem_w_8 ( .clk(clk), .addr(addr_w_8), .z(
        data_out_w_8) );
  layer2_12_8_12_16_B_rom_8 mem_b_8 ( .clk(clk), .addr(\addr_b_8[0] ) );
  layer2_12_8_12_16_W_rom_9 mem_w_9 ( .clk(clk), .addr(addr_w_9), .z(
        data_out_w_9) );
  layer2_12_8_12_16_B_rom_9 mem_b_9 ( .clk(clk), .addr(\addr_b_9[0] ) );
  layer2_12_8_12_16_W_rom_10 mem_w_10 ( .clk(clk), .addr(addr_w_10), .z(
        data_out_w_10) );
  layer2_12_8_12_16_B_rom_10 mem_b_10 ( .clk(clk), .addr(\addr_b_10[0] ) );
  layer2_12_8_12_16_W_rom_11 mem_w_11 ( .clk(clk), .addr(addr_w_11), .z({
        data_out_w_11[15:4], SYNOPSYS_UNCONNECTED__0, data_out_w_11[2:0]}) );
  layer2_12_8_12_16_B_rom_11 mem_b_11 ( .clk(clk), .addr(\addr_b_11[0] ) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_0 d_0 ( .clk(clk), .clear_acc(
        clear_acc), .data_out_x({n87, n120, data_out_x[13], n119, 
        data_out_x[11], n91, n88, n96, n116, n1, n104, n113, n101, n92, n108, 
        n90}), .data_out(data_out_0), .data_out_w(data_out_w_0), .data_out_b({
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 
        1'b0, 1'b0, 1'b1, 1'b1}), .wr_en_y(wr_en_y), .m_valid(m_valid), 
        .m_ready(n105), .sel(sel) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_11 d_1 ( .clk(clk), .clear_acc(
        clear_acc), .data_out_x({data_out_x[15], n120, data_out_x[13], n119, 
        data_out_x[11], n118, data_out_x[9], n96, n95, n97, n104, n94, n101, 
        n98, n108, n86}), .data_out(data_out_1), .data_out_w(data_out_w_1), 
        .data_out_b({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1}), .wr_en_y(wr_en_y), 
        .m_valid(m_valid), .m_ready(n106), .sel(sel) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_10 d_2 ( .clk(clk), .clear_acc(
        clear_acc), .data_out_x({n87, n3, data_out_x[13], n119, data_out_x[11], 
        n91, data_out_x[9], n117, n116, n1, n104, n94, n101, n92, n107, n86}), 
        .data_out(data_out_2), .data_out_w(data_out_w_2), .data_out_b({1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b1, 1'b0}), .wr_en_y(wr_en_y), .m_valid(m_valid), .m_ready(
        n106), .sel(sel) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_9 d_3 ( .clk(clk), .clear_acc(
        clear_acc), .data_out_x({n87, n120, data_out_x[13], n119, 
        data_out_x[11], n91, data_out_x[9], n117, n99, n115, n103, n113, n112, 
        n111, n110, n89}), .data_out(data_out_3), .data_out_w(data_out_w_3), 
        .data_out_b({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0}), .wr_en_y(wr_en_y), 
        .m_valid(m_valid), .m_ready(n105), .sel(sel) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_8 d_4 ( .clk(clk), .clear_acc(
        clear_acc), .data_out_x({n87, n3, data_out_x[13], n119, data_out_x[11], 
        n118, data_out_x[9], n117, n99, n2, n103, n94, n102, n111, n108, n109}), .data_out(data_out_4), .data_out_w(data_out_w_4), .data_out_b({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 
        1'b0, 1'b1}), .wr_en_y(wr_en_y), .m_valid(m_valid), .m_ready(n106), 
        .sel(sel) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_7 d_5 ( .clk(clk), .clear_acc(
        clear_acc), .data_out_x({n121, n3, data_out_x[13], n119, 
        data_out_x[11], n91, n85, n96, n95, n1, n103, n94, n101, n98, n107, 
        n89}), .data_out(data_out_5), .data_out_w(data_out_w_5), .data_out_b({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 
        1'b0, 1'b1, 1'b0, 1'b1}), .wr_en_y(wr_en_y), .m_valid(m_valid), 
        .m_ready(n106), .sel(sel) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_6 d_6 ( .clk(clk), .clear_acc(
        clear_acc), .data_out_x({n87, n3, data_out_x[13], n119, data_out_x[11], 
        n100, data_out_x[9], n117, n116, n115, n104, n113, n102, n98, n107, 
        n89}), .data_out(data_out_6), .data_out_w(data_out_w_6), .data_out_b({
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 
        1'b1, 1'b0, 1'b1, 1'b1}), .wr_en_y(wr_en_y), .m_valid(m_valid), 
        .m_ready(n105), .sel(sel) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_5 d_7 ( .clk(clk), .clear_acc(
        clear_acc), .data_out_x({n121, n120, data_out_x[13], n119, 
        data_out_x[11], n118, data_out_x[9], n96, n95, n115, n114, n94, n101, 
        n98, n110, n86}), .data_out(data_out_7), .data_out_w(data_out_w_7), 
        .data_out_b({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1}), .wr_en_y(wr_en_y), 
        .m_valid(m_valid), .m_ready(n105), .sel(sel) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_4 d_8 ( .clk(clk), .clear_acc(
        clear_acc), .data_out_x({data_out_x[15], n120, data_out_x[13], n119, 
        data_out_x[11], n100, n93, n96, n116, n97, n114, n94, n102, n92, n108, 
        n86}), .data_out(data_out_8), .data_out_w(data_out_w_8), .data_out_b({
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 
        1'b1, 1'b1, 1'b1, 1'b1}), .wr_en_y(wr_en_y), .m_valid(m_valid), 
        .m_ready(n105), .sel(sel) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_3 d_9 ( .clk(clk), .clear_acc(
        clear_acc), .data_out_x({n121, n3, data_out_x[13], n119, 
        data_out_x[11], n91, data_out_x[9], n117, n99, n2, n103, n113, n112, 
        n111, n110, n90}), .data_out(data_out_9), .data_out_w(data_out_w_9), 
        .data_out_b({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1}), .wr_en_y(wr_en_y), 
        .m_valid(m_valid), .m_ready(n105), .sel(sel) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_2 d_10 ( .clk(clk), .clear_acc(
        clear_acc), .data_out_x({data_out_x[15], n3, data_out_x[13], n119, 
        data_out_x[11], n118, data_out_x[9], n96, n95, n115, n104, n113, n102, 
        n111, n107, n109}), .data_out(data_out_10), .data_out_w(data_out_w_10), 
        .data_out_b({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1}), .wr_en_y(wr_en_y), 
        .m_valid(m_valid), .m_ready(n106), .sel(sel) );
  layer2_12_8_12_16_datapath_M12_N8_T16_P12_1 d_11 ( .clk(clk), .clear_acc(
        clear_acc), .data_out_x({data_out_x[15], n120, data_out_x[13], n119, 
        data_out_x[11], n118, data_out_x[9], n117, n99, n2, n103, n113, n112, 
        n92, n107, n90}), .data_out(data_out_11), .data_out_w({
        data_out_w_11[15:4], 1'b0, data_out_w_11[2:0]}), .data_out_b({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 
        1'b0, 1'b0, 1'b1}), .wr_en_y(wr_en_y), .m_valid(m_valid), .m_ready(
        n106), .sel(sel) );
  layer2_12_8_12_16_ctrlpath_M12_N8_T16_P12 c ( .clk(clk), .reset(reset), 
        .s_valid(s_valid), .s_ready(s_ready), .m_valid(m_valid), .m_ready(
        m_ready), .clear_acc(clear_acc), .wr_en_x(wr_en_x), .wr_en_y(wr_en_y), 
        .sel(sel), .addr_x(addr_x), .addr_w_0(addr_w_0), .addr_b_0(
        \addr_b_0[0] ), .addr_w_1(addr_w_1), .addr_b_1(\addr_b_1[0] ), 
        .addr_w_2(addr_w_2), .addr_b_2(\addr_b_2[0] ), .addr_w_3(addr_w_3), 
        .addr_b_3(\addr_b_3[0] ), .addr_w_4(addr_w_4), .addr_b_4(\addr_b_4[0] ), .addr_w_5(addr_w_5), .addr_b_5(\addr_b_5[0] ), .addr_w_6(addr_w_6), 
        .addr_b_6(\addr_b_6[0] ), .addr_w_7(addr_w_7), .addr_b_7(\addr_b_7[0] ), .addr_w_8(addr_w_8), .addr_b_8(\addr_b_8[0] ), .addr_w_9(addr_w_9), 
        .addr_b_9(\addr_b_9[0] ), .addr_w_10(addr_w_10), .addr_b_10(
        \addr_b_10[0] ), .addr_w_11(addr_w_11), .addr_b_11(\addr_b_11[0] ) );
  BUF_X1 U1 ( .A(data_out_x[10]), .Z(n100) );
  CLKBUF_X3 U2 ( .A(data_out_x[6]), .Z(n1) );
  CLKBUF_X3 U3 ( .A(data_out_x[6]), .Z(n2) );
  BUF_X1 U4 ( .A(data_out_x[6]), .Z(n97) );
  CLKBUF_X3 U5 ( .A(data_out_x[7]), .Z(n116) );
  CLKBUF_X3 U6 ( .A(data_out_x[5]), .Z(n104) );
  CLKBUF_X3 U7 ( .A(data_out_x[4]), .Z(n94) );
  BUF_X2 U8 ( .A(data_out_x[0]), .Z(n109) );
  CLKBUF_X3 U9 ( .A(data_out_x[4]), .Z(n113) );
  BUF_X1 U10 ( .A(data_out_x[9]), .Z(n85) );
  BUF_X1 U11 ( .A(data_out_x[5]), .Z(n114) );
  BUF_X1 U12 ( .A(data_out_x[9]), .Z(n93) );
  BUF_X1 U13 ( .A(data_out_x[9]), .Z(n88) );
  CLKBUF_X3 U14 ( .A(data_out_x[10]), .Z(n118) );
  BUF_X2 U15 ( .A(data_out_x[14]), .Z(n3) );
  CLKBUF_X3 U16 ( .A(data_out_x[0]), .Z(n86) );
  BUF_X1 U17 ( .A(data_out_x[3]), .Z(n112) );
  CLKBUF_X3 U18 ( .A(data_out_x[2]), .Z(n111) );
  CLKBUF_X3 U19 ( .A(data_out_x[0]), .Z(n90) );
  BUF_X2 U20 ( .A(data_out_x[3]), .Z(n102) );
  BUF_X1 U21 ( .A(data_out_x[15]), .Z(n87) );
  CLKBUF_X3 U22 ( .A(data_out_x[2]), .Z(n92) );
  CLKBUF_X3 U23 ( .A(data_out_x[0]), .Z(n89) );
  CLKBUF_X3 U24 ( .A(data_out_x[10]), .Z(n91) );
  CLKBUF_X3 U25 ( .A(data_out_x[2]), .Z(n98) );
  CLKBUF_X3 U26 ( .A(data_out_x[7]), .Z(n95) );
  BUF_X4 U27 ( .A(data_out_x[12]), .Z(n119) );
  BUF_X4 U28 ( .A(data_out_x[6]), .Z(n115) );
  BUF_X2 U29 ( .A(data_out_x[7]), .Z(n99) );
  BUF_X2 U30 ( .A(data_out_x[1]), .Z(n107) );
  BUF_X1 U31 ( .A(data_out_x[1]), .Z(n110) );
  BUF_X2 U32 ( .A(data_out_x[5]), .Z(n103) );
  BUF_X4 U33 ( .A(data_out_x[8]), .Z(n96) );
  CLKBUF_X3 U34 ( .A(data_out_x[1]), .Z(n108) );
  BUF_X2 U35 ( .A(data_out_x[3]), .Z(n101) );
  CLKBUF_X1 U36 ( .A(m_ready), .Z(n105) );
  CLKBUF_X1 U37 ( .A(m_ready), .Z(n106) );
  BUF_X2 U38 ( .A(data_out_x[14]), .Z(n120) );
  BUF_X1 U39 ( .A(data_out_x[15]), .Z(n121) );
  AND2_X1 U40 ( .A1(n84), .A2(n80), .ZN(n18) );
  AND2_X1 U41 ( .A1(n83), .A2(n82), .ZN(n19) );
  AND2_X1 U42 ( .A1(n84), .A2(n82), .ZN(n17) );
  AND2_X1 U43 ( .A1(n83), .A2(n80), .ZN(n14) );
  NOR2_X2 U44 ( .A1(n124), .A2(n81), .ZN(n9) );
  INV_X1 U45 ( .A(sel[3]), .ZN(n124) );
  AOI21_X1 U46 ( .B1(n80), .B2(sel[0]), .A(sel[2]), .ZN(n81) );
  AND3_X1 U47 ( .A1(sel[3]), .A2(n122), .A3(n82), .ZN(n12) );
  AND3_X1 U48 ( .A1(n83), .A2(n123), .A3(sel[2]), .ZN(n15) );
  NAND4_X1 U49 ( .A1(n76), .A2(n77), .A3(n78), .A4(n79), .ZN(data_out[0]) );
  AOI222_X1 U50 ( .A1(data_out_0[0]), .A2(n17), .B1(data_out_2[0]), .B2(n18), 
        .C1(data_out_1[0]), .C2(n19), .ZN(n76) );
  AOI222_X1 U51 ( .A1(data_out_3[0]), .A2(n14), .B1(data_out_5[0]), .B2(n15), 
        .C1(data_out_4[0]), .C2(n16), .ZN(n77) );
  AOI222_X1 U52 ( .A1(data_out_6[0]), .A2(n11), .B1(data_out_8[0]), .B2(n12), 
        .C1(data_out_7[0]), .C2(n13), .ZN(n78) );
  NAND4_X1 U53 ( .A1(n48), .A2(n49), .A3(n50), .A4(n51), .ZN(data_out[1]) );
  AOI222_X1 U54 ( .A1(data_out_0[1]), .A2(n17), .B1(data_out_2[1]), .B2(n18), 
        .C1(data_out_1[1]), .C2(n19), .ZN(n48) );
  AOI222_X1 U55 ( .A1(data_out_3[1]), .A2(n14), .B1(data_out_5[1]), .B2(n15), 
        .C1(data_out_4[1]), .C2(n16), .ZN(n49) );
  AOI222_X1 U56 ( .A1(data_out_6[1]), .A2(n11), .B1(data_out_8[1]), .B2(n12), 
        .C1(data_out_7[1]), .C2(n13), .ZN(n50) );
  NAND4_X1 U57 ( .A1(n44), .A2(n45), .A3(n46), .A4(n47), .ZN(data_out[2]) );
  AOI222_X1 U58 ( .A1(data_out_0[2]), .A2(n17), .B1(data_out_2[2]), .B2(n18), 
        .C1(data_out_1[2]), .C2(n19), .ZN(n44) );
  AOI222_X1 U59 ( .A1(data_out_3[2]), .A2(n14), .B1(data_out_5[2]), .B2(n15), 
        .C1(data_out_4[2]), .C2(n16), .ZN(n45) );
  AOI222_X1 U60 ( .A1(data_out_6[2]), .A2(n11), .B1(data_out_8[2]), .B2(n12), 
        .C1(data_out_7[2]), .C2(n13), .ZN(n46) );
  NAND4_X1 U61 ( .A1(n40), .A2(n41), .A3(n42), .A4(n43), .ZN(data_out[3]) );
  AOI222_X1 U62 ( .A1(data_out_0[3]), .A2(n17), .B1(data_out_2[3]), .B2(n18), 
        .C1(data_out_1[3]), .C2(n19), .ZN(n40) );
  AOI222_X1 U63 ( .A1(data_out_3[3]), .A2(n14), .B1(data_out_5[3]), .B2(n15), 
        .C1(data_out_4[3]), .C2(n16), .ZN(n41) );
  AOI222_X1 U64 ( .A1(data_out_6[3]), .A2(n11), .B1(data_out_8[3]), .B2(n12), 
        .C1(data_out_7[3]), .C2(n13), .ZN(n42) );
  NAND4_X1 U65 ( .A1(n36), .A2(n37), .A3(n38), .A4(n39), .ZN(data_out[4]) );
  AOI222_X1 U66 ( .A1(data_out_0[4]), .A2(n17), .B1(data_out_2[4]), .B2(n18), 
        .C1(data_out_1[4]), .C2(n19), .ZN(n36) );
  AOI222_X1 U67 ( .A1(data_out_3[4]), .A2(n14), .B1(data_out_5[4]), .B2(n15), 
        .C1(data_out_4[4]), .C2(n16), .ZN(n37) );
  AOI222_X1 U68 ( .A1(data_out_6[4]), .A2(n11), .B1(data_out_8[4]), .B2(n12), 
        .C1(data_out_7[4]), .C2(n13), .ZN(n38) );
  NAND4_X1 U69 ( .A1(n32), .A2(n33), .A3(n34), .A4(n35), .ZN(data_out[5]) );
  AOI222_X1 U70 ( .A1(data_out_0[5]), .A2(n17), .B1(data_out_2[5]), .B2(n18), 
        .C1(data_out_1[5]), .C2(n19), .ZN(n32) );
  AOI222_X1 U71 ( .A1(data_out_3[5]), .A2(n14), .B1(data_out_5[5]), .B2(n15), 
        .C1(data_out_4[5]), .C2(n16), .ZN(n33) );
  AOI222_X1 U72 ( .A1(data_out_6[5]), .A2(n11), .B1(data_out_8[5]), .B2(n12), 
        .C1(data_out_7[5]), .C2(n13), .ZN(n34) );
  NAND4_X1 U73 ( .A1(n28), .A2(n29), .A3(n30), .A4(n31), .ZN(data_out[6]) );
  AOI222_X1 U74 ( .A1(data_out_0[6]), .A2(n17), .B1(data_out_2[6]), .B2(n18), 
        .C1(data_out_1[6]), .C2(n19), .ZN(n28) );
  AOI222_X1 U75 ( .A1(data_out_3[6]), .A2(n14), .B1(data_out_5[6]), .B2(n15), 
        .C1(data_out_4[6]), .C2(n16), .ZN(n29) );
  AOI222_X1 U76 ( .A1(data_out_6[6]), .A2(n11), .B1(data_out_8[6]), .B2(n12), 
        .C1(data_out_7[6]), .C2(n13), .ZN(n30) );
  NAND4_X1 U77 ( .A1(n24), .A2(n25), .A3(n26), .A4(n27), .ZN(data_out[7]) );
  AOI222_X1 U78 ( .A1(data_out_0[7]), .A2(n17), .B1(data_out_2[7]), .B2(n18), 
        .C1(data_out_1[7]), .C2(n19), .ZN(n24) );
  AOI222_X1 U79 ( .A1(data_out_3[7]), .A2(n14), .B1(data_out_5[7]), .B2(n15), 
        .C1(data_out_4[7]), .C2(n16), .ZN(n25) );
  AOI222_X1 U80 ( .A1(data_out_6[7]), .A2(n11), .B1(data_out_8[7]), .B2(n12), 
        .C1(data_out_7[7]), .C2(n13), .ZN(n26) );
  NAND4_X1 U81 ( .A1(n20), .A2(n21), .A3(n22), .A4(n23), .ZN(data_out[8]) );
  AOI222_X1 U82 ( .A1(data_out_0[8]), .A2(n17), .B1(data_out_2[8]), .B2(n18), 
        .C1(data_out_1[8]), .C2(n19), .ZN(n20) );
  AOI222_X1 U84 ( .A1(data_out_3[8]), .A2(n14), .B1(data_out_5[8]), .B2(n15), 
        .C1(data_out_4[8]), .C2(n16), .ZN(n21) );
  AOI222_X1 U86 ( .A1(data_out_6[8]), .A2(n11), .B1(data_out_8[8]), .B2(n12), 
        .C1(data_out_7[8]), .C2(n13), .ZN(n22) );
  NAND4_X1 U88 ( .A1(n4), .A2(n5), .A3(n6), .A4(n7), .ZN(data_out[9]) );
  AOI222_X1 U89 ( .A1(data_out_0[9]), .A2(n17), .B1(data_out_2[9]), .B2(n18), 
        .C1(data_out_1[9]), .C2(n19), .ZN(n4) );
  AOI222_X1 U90 ( .A1(data_out_3[9]), .A2(n14), .B1(data_out_5[9]), .B2(n15), 
        .C1(data_out_4[9]), .C2(n16), .ZN(n5) );
  AOI222_X1 U91 ( .A1(data_out_6[9]), .A2(n11), .B1(data_out_8[9]), .B2(n12), 
        .C1(data_out_7[9]), .C2(n13), .ZN(n6) );
  NAND4_X1 U92 ( .A1(n72), .A2(n73), .A3(n74), .A4(n75), .ZN(data_out[10]) );
  AOI222_X1 U93 ( .A1(data_out_0[10]), .A2(n17), .B1(data_out_2[10]), .B2(n18), 
        .C1(data_out_1[10]), .C2(n19), .ZN(n72) );
  AOI222_X1 U94 ( .A1(data_out_3[10]), .A2(n14), .B1(data_out_5[10]), .B2(n15), 
        .C1(data_out_4[10]), .C2(n16), .ZN(n73) );
  AOI222_X1 U95 ( .A1(data_out_6[10]), .A2(n11), .B1(data_out_8[10]), .B2(n12), 
        .C1(data_out_7[10]), .C2(n13), .ZN(n74) );
  NAND4_X1 U96 ( .A1(n68), .A2(n69), .A3(n70), .A4(n71), .ZN(data_out[11]) );
  AOI222_X1 U97 ( .A1(data_out_0[11]), .A2(n17), .B1(data_out_2[11]), .B2(n18), 
        .C1(data_out_1[11]), .C2(n19), .ZN(n68) );
  AOI222_X1 U98 ( .A1(data_out_3[11]), .A2(n14), .B1(data_out_5[11]), .B2(n15), 
        .C1(data_out_4[11]), .C2(n16), .ZN(n69) );
  AOI222_X1 U99 ( .A1(data_out_6[11]), .A2(n11), .B1(data_out_8[11]), .B2(n12), 
        .C1(data_out_7[11]), .C2(n13), .ZN(n70) );
  NAND4_X1 U100 ( .A1(n64), .A2(n65), .A3(n66), .A4(n67), .ZN(data_out[12]) );
  AOI222_X1 U101 ( .A1(data_out_0[12]), .A2(n17), .B1(data_out_2[12]), .B2(n18), .C1(data_out_1[12]), .C2(n19), .ZN(n64) );
  AOI222_X1 U102 ( .A1(data_out_3[12]), .A2(n14), .B1(data_out_5[12]), .B2(n15), .C1(data_out_4[12]), .C2(n16), .ZN(n65) );
  AOI222_X1 U103 ( .A1(data_out_6[12]), .A2(n11), .B1(data_out_8[12]), .B2(n12), .C1(data_out_7[12]), .C2(n13), .ZN(n66) );
  NAND4_X1 U104 ( .A1(n60), .A2(n61), .A3(n62), .A4(n63), .ZN(data_out[13]) );
  AOI222_X1 U105 ( .A1(data_out_0[13]), .A2(n17), .B1(data_out_2[13]), .B2(n18), .C1(data_out_1[13]), .C2(n19), .ZN(n60) );
  AOI222_X1 U106 ( .A1(data_out_3[13]), .A2(n14), .B1(data_out_5[13]), .B2(n15), .C1(data_out_4[13]), .C2(n16), .ZN(n61) );
  AOI222_X1 U107 ( .A1(data_out_6[13]), .A2(n11), .B1(data_out_8[13]), .B2(n12), .C1(data_out_7[13]), .C2(n13), .ZN(n62) );
  NAND4_X1 U108 ( .A1(n56), .A2(n57), .A3(n58), .A4(n59), .ZN(data_out[14]) );
  AOI222_X1 U109 ( .A1(data_out_0[14]), .A2(n17), .B1(data_out_2[14]), .B2(n18), .C1(data_out_1[14]), .C2(n19), .ZN(n56) );
  AOI222_X1 U110 ( .A1(data_out_3[14]), .A2(n14), .B1(data_out_5[14]), .B2(n15), .C1(data_out_4[14]), .C2(n16), .ZN(n57) );
  AOI222_X1 U111 ( .A1(data_out_6[14]), .A2(n11), .B1(data_out_8[14]), .B2(n12), .C1(data_out_7[14]), .C2(n13), .ZN(n58) );
  NAND4_X1 U112 ( .A1(n52), .A2(n53), .A3(n54), .A4(n55), .ZN(data_out[15]) );
  AOI222_X1 U113 ( .A1(data_out_0[15]), .A2(n17), .B1(data_out_2[15]), .B2(n18), .C1(data_out_1[15]), .C2(n19), .ZN(n52) );
  AOI222_X1 U114 ( .A1(data_out_3[15]), .A2(n14), .B1(data_out_5[15]), .B2(n15), .C1(data_out_4[15]), .C2(n16), .ZN(n53) );
  AOI222_X1 U115 ( .A1(data_out_6[15]), .A2(n11), .B1(data_out_8[15]), .B2(n12), .C1(data_out_7[15]), .C2(n13), .ZN(n54) );
  AND3_X1 U116 ( .A1(n80), .A2(n122), .A3(sel[3]), .ZN(n10) );
  AND3_X1 U117 ( .A1(sel[3]), .A2(sel[0]), .A3(n82), .ZN(n8) );
  AOI222_X1 U118 ( .A1(data_out_9[0]), .A2(n8), .B1(data_out_11[0]), .B2(n9), 
        .C1(data_out_10[0]), .C2(n10), .ZN(n79) );
  AOI222_X1 U119 ( .A1(data_out_9[1]), .A2(n8), .B1(data_out_11[1]), .B2(n9), 
        .C1(data_out_10[1]), .C2(n10), .ZN(n51) );
  AOI222_X1 U120 ( .A1(data_out_9[2]), .A2(n8), .B1(data_out_11[2]), .B2(n9), 
        .C1(data_out_10[2]), .C2(n10), .ZN(n47) );
  AOI222_X1 U121 ( .A1(data_out_9[3]), .A2(n8), .B1(data_out_11[3]), .B2(n9), 
        .C1(data_out_10[3]), .C2(n10), .ZN(n43) );
  AOI222_X1 U122 ( .A1(data_out_9[4]), .A2(n8), .B1(data_out_11[4]), .B2(n9), 
        .C1(data_out_10[4]), .C2(n10), .ZN(n39) );
  AOI222_X1 U123 ( .A1(data_out_9[5]), .A2(n8), .B1(data_out_11[5]), .B2(n9), 
        .C1(data_out_10[5]), .C2(n10), .ZN(n35) );
  AOI222_X1 U124 ( .A1(data_out_9[6]), .A2(n8), .B1(data_out_11[6]), .B2(n9), 
        .C1(data_out_10[6]), .C2(n10), .ZN(n31) );
  AOI222_X1 U125 ( .A1(data_out_9[7]), .A2(n8), .B1(data_out_11[7]), .B2(n9), 
        .C1(data_out_10[7]), .C2(n10), .ZN(n27) );
  AOI222_X1 U126 ( .A1(data_out_9[8]), .A2(n8), .B1(data_out_11[8]), .B2(n9), 
        .C1(data_out_10[8]), .C2(n10), .ZN(n23) );
  AOI222_X1 U127 ( .A1(data_out_9[9]), .A2(n8), .B1(data_out_11[9]), .B2(n9), 
        .C1(data_out_10[9]), .C2(n10), .ZN(n7) );
  AOI222_X1 U128 ( .A1(data_out_9[10]), .A2(n8), .B1(data_out_11[10]), .B2(n9), 
        .C1(data_out_10[10]), .C2(n10), .ZN(n75) );
  AOI222_X1 U129 ( .A1(data_out_9[11]), .A2(n8), .B1(data_out_11[11]), .B2(n9), 
        .C1(data_out_10[11]), .C2(n10), .ZN(n71) );
  AOI222_X1 U130 ( .A1(data_out_9[12]), .A2(n8), .B1(data_out_11[12]), .B2(n9), 
        .C1(data_out_10[12]), .C2(n10), .ZN(n67) );
  AOI222_X1 U131 ( .A1(data_out_9[13]), .A2(n8), .B1(data_out_11[13]), .B2(n9), 
        .C1(data_out_10[13]), .C2(n10), .ZN(n63) );
  AOI222_X1 U132 ( .A1(data_out_9[14]), .A2(n8), .B1(data_out_11[14]), .B2(n9), 
        .C1(data_out_10[14]), .C2(n10), .ZN(n59) );
  AOI222_X1 U133 ( .A1(data_out_9[15]), .A2(n8), .B1(data_out_11[15]), .B2(n9), 
        .C1(data_out_10[15]), .C2(n10), .ZN(n55) );
  NOR2_X1 U134 ( .A1(n123), .A2(sel[2]), .ZN(n80) );
  NOR2_X1 U135 ( .A1(sel[2]), .A2(sel[1]), .ZN(n82) );
  BUF_X4 U136 ( .A(data_out_x[8]), .Z(n117) );
  NOR2_X1 U137 ( .A1(sel[3]), .A2(sel[0]), .ZN(n84) );
  NOR2_X1 U138 ( .A1(n122), .A2(sel[3]), .ZN(n83) );
  INV_X1 U139 ( .A(sel[1]), .ZN(n123) );
  INV_X1 U140 ( .A(sel[0]), .ZN(n122) );
endmodule


module memory_WIDTH16_SIZE12_LOGSIZE4 ( clk, data_in, data_out, addr, wr_en );
  input [15:0] data_in;
  output [15:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   \mem[11][15] , \mem[11][14] , \mem[11][13] , \mem[11][12] ,
         \mem[11][11] , \mem[11][10] , \mem[11][9] , \mem[11][8] ,
         \mem[11][7] , \mem[11][6] , \mem[11][5] , \mem[11][4] , \mem[11][3] ,
         \mem[11][2] , \mem[11][1] , \mem[11][0] , \mem[10][15] ,
         \mem[10][14] , \mem[10][13] , \mem[10][12] , \mem[10][11] ,
         \mem[10][10] , \mem[10][9] , \mem[10][8] , \mem[10][7] , \mem[10][6] ,
         \mem[10][5] , \mem[10][4] , \mem[10][3] , \mem[10][2] , \mem[10][1] ,
         \mem[10][0] , \mem[9][15] , \mem[9][14] , \mem[9][13] , \mem[9][12] ,
         \mem[9][11] , \mem[9][10] , \mem[9][9] , \mem[9][8] , \mem[9][7] ,
         \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] ,
         \mem[9][1] , \mem[9][0] , \mem[8][15] , \mem[8][14] , \mem[8][13] ,
         \mem[8][12] , \mem[8][11] , \mem[8][10] , \mem[8][9] , \mem[8][8] ,
         \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] , \mem[8][3] ,
         \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][15] , \mem[7][14] ,
         \mem[7][13] , \mem[7][12] , \mem[7][11] , \mem[7][10] , \mem[7][9] ,
         \mem[7][8] , \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] ,
         \mem[7][3] , \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][15] ,
         \mem[6][14] , \mem[6][13] , \mem[6][12] , \mem[6][11] , \mem[6][10] ,
         \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][15] , \mem[5][14] , \mem[5][13] , \mem[5][12] , \mem[5][11] ,
         \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[4][15] , \mem[4][14] , \mem[4][13] , \mem[4][12] ,
         \mem[4][11] , \mem[4][10] , \mem[4][9] , \mem[4][8] , \mem[4][7] ,
         \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] ,
         \mem[4][1] , \mem[4][0] , \mem[3][15] , \mem[3][14] , \mem[3][13] ,
         \mem[3][12] , \mem[3][11] , \mem[3][10] , \mem[3][9] , \mem[3][8] ,
         \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] , \mem[3][3] ,
         \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][15] , \mem[2][14] ,
         \mem[2][13] , \mem[2][12] , \mem[2][11] , \mem[2][10] , \mem[2][9] ,
         \mem[2][8] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][15] ,
         \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] , \mem[1][10] ,
         \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64,
         N65, N66, N67, N68, N69, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476;

  DFF_X1 \mem_reg[11][15]  ( .D(n53), .CK(clk), .Q(\mem[11][15] ) );
  DFF_X1 \mem_reg[11][14]  ( .D(n65), .CK(clk), .Q(\mem[11][14] ) );
  DFF_X1 \mem_reg[11][13]  ( .D(n77), .CK(clk), .Q(\mem[11][13] ) );
  DFF_X1 \mem_reg[11][12]  ( .D(n89), .CK(clk), .Q(\mem[11][12] ) );
  DFF_X1 \mem_reg[11][11]  ( .D(n101), .CK(clk), .Q(\mem[11][11] ) );
  DFF_X1 \mem_reg[11][10]  ( .D(n113), .CK(clk), .Q(\mem[11][10] ) );
  DFF_X1 \mem_reg[11][9]  ( .D(n125), .CK(clk), .Q(\mem[11][9] ) );
  DFF_X1 \mem_reg[11][8]  ( .D(n137), .CK(clk), .Q(\mem[11][8] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n149), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n161), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n173), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n185), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n197), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n427), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n439), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n451), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][15]  ( .D(n54), .CK(clk), .Q(\mem[10][15] ) );
  DFF_X1 \mem_reg[10][14]  ( .D(n66), .CK(clk), .Q(\mem[10][14] ) );
  DFF_X1 \mem_reg[10][13]  ( .D(n78), .CK(clk), .Q(\mem[10][13] ) );
  DFF_X1 \mem_reg[10][12]  ( .D(n90), .CK(clk), .Q(\mem[10][12] ) );
  DFF_X1 \mem_reg[10][11]  ( .D(n102), .CK(clk), .Q(\mem[10][11] ) );
  DFF_X1 \mem_reg[10][10]  ( .D(n114), .CK(clk), .Q(\mem[10][10] ) );
  DFF_X1 \mem_reg[10][9]  ( .D(n126), .CK(clk), .Q(\mem[10][9] ) );
  DFF_X1 \mem_reg[10][8]  ( .D(n138), .CK(clk), .Q(\mem[10][8] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n150), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n162), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n174), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n186), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n198), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n428), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n440), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n452), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][15]  ( .D(n55), .CK(clk), .Q(\mem[9][15] ) );
  DFF_X1 \mem_reg[9][14]  ( .D(n67), .CK(clk), .Q(\mem[9][14] ) );
  DFF_X1 \mem_reg[9][13]  ( .D(n79), .CK(clk), .Q(\mem[9][13] ) );
  DFF_X1 \mem_reg[9][12]  ( .D(n91), .CK(clk), .Q(\mem[9][12] ) );
  DFF_X1 \mem_reg[9][11]  ( .D(n103), .CK(clk), .Q(\mem[9][11] ) );
  DFF_X1 \mem_reg[9][10]  ( .D(n115), .CK(clk), .Q(\mem[9][10] ) );
  DFF_X1 \mem_reg[9][9]  ( .D(n127), .CK(clk), .Q(\mem[9][9] ) );
  DFF_X1 \mem_reg[9][8]  ( .D(n139), .CK(clk), .Q(\mem[9][8] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n151), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n163), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n175), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n187), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n199), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n429), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n441), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n453), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][15]  ( .D(n56), .CK(clk), .Q(\mem[8][15] ) );
  DFF_X1 \mem_reg[8][14]  ( .D(n68), .CK(clk), .Q(\mem[8][14] ) );
  DFF_X1 \mem_reg[8][13]  ( .D(n80), .CK(clk), .Q(\mem[8][13] ) );
  DFF_X1 \mem_reg[8][12]  ( .D(n92), .CK(clk), .Q(\mem[8][12] ) );
  DFF_X1 \mem_reg[8][11]  ( .D(n104), .CK(clk), .Q(\mem[8][11] ) );
  DFF_X1 \mem_reg[8][10]  ( .D(n116), .CK(clk), .Q(\mem[8][10] ) );
  DFF_X1 \mem_reg[8][9]  ( .D(n128), .CK(clk), .Q(\mem[8][9] ) );
  DFF_X1 \mem_reg[8][8]  ( .D(n140), .CK(clk), .Q(\mem[8][8] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n152), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n164), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n176), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n188), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n200), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n430), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n442), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n454), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][15]  ( .D(n57), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n69), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n81), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n93), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n105), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n117), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n129), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n141), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n153), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n165), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n177), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n189), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n201), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n431), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n443), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n455), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n58), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n70), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n82), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n94), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n106), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n118), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n130), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n142), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n154), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n166), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n178), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n190), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n202), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n432), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n444), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n456), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n59), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n71), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n83), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n95), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n107), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n119), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n131), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n143), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n155), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n167), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n179), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n191), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n203), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n433), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n445), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n457), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n60), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n72), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n84), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n96), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n108), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n120), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n132), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n144), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n156), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n168), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n180), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n192), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n204), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n434), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n446), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n458), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n61), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n73), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n85), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n97), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n109), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n121), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n133), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n145), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n157), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n169), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n181), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n193), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n205), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n435), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n447), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n459), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n62), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n74), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n86), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n98), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n110), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n122), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n134), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n146), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n158), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n170), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n182), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n194), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n206), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n436), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n448), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n460), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n63), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n75), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n87), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n99), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n111), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n123), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n135), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n147), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n159), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n171), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n183), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n195), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n425), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n437), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n449), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n461), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n64), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(N54), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n76), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(N55), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n88), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(N56), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n100), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(N57), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n112), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(N58), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n124), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(N59), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n136), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(N60), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n148), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(N61), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n160), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(N62), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n172), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(N63), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n184), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(N64), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n196), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(N65), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n426), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(N66), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n438), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(N67), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n450), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(N68), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n462), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(N69), .CK(clk), .Q(data_out[0]) );
  INV_X1 U3 ( .A(n353), .ZN(n470) );
  INV_X1 U4 ( .A(n299), .ZN(n465) );
  INV_X1 U5 ( .A(n226), .ZN(n474) );
  INV_X1 U6 ( .A(n244), .ZN(n473) );
  INV_X1 U7 ( .A(n262), .ZN(n472) );
  INV_X1 U8 ( .A(n372), .ZN(n469) );
  INV_X1 U9 ( .A(n390), .ZN(n468) );
  INV_X1 U10 ( .A(n408), .ZN(n467) );
  INV_X1 U11 ( .A(n280), .ZN(n466) );
  INV_X1 U12 ( .A(n317), .ZN(n464) );
  INV_X1 U13 ( .A(n335), .ZN(n463) );
  INV_X1 U14 ( .A(n208), .ZN(n475) );
  NAND2_X1 U15 ( .A1(wr_en), .A2(n224), .ZN(n208) );
  NAND2_X1 U16 ( .A1(n369), .A2(n370), .ZN(n353) );
  NAND2_X1 U17 ( .A1(n388), .A2(n370), .ZN(n372) );
  NAND2_X1 U18 ( .A1(n406), .A2(n370), .ZN(n390) );
  NAND2_X1 U19 ( .A1(n424), .A2(n370), .ZN(n408) );
  NAND2_X1 U20 ( .A1(n296), .A2(n297), .ZN(n280) );
  NAND2_X1 U21 ( .A1(n315), .A2(n297), .ZN(n299) );
  NAND2_X1 U22 ( .A1(n333), .A2(n297), .ZN(n317) );
  NAND2_X1 U23 ( .A1(n351), .A2(n297), .ZN(n335) );
  NAND2_X1 U24 ( .A1(n242), .A2(wr_en), .ZN(n226) );
  NAND2_X1 U25 ( .A1(n260), .A2(wr_en), .ZN(n244) );
  NAND2_X1 U26 ( .A1(n278), .A2(wr_en), .ZN(n262) );
  AND2_X1 U27 ( .A1(n491), .A2(n493), .ZN(n242) );
  AND2_X1 U28 ( .A1(n493), .A2(n492), .ZN(n224) );
  AND2_X1 U29 ( .A1(n489), .A2(n493), .ZN(n260) );
  AND2_X1 U30 ( .A1(n490), .A2(n493), .ZN(n278) );
  INV_X1 U31 ( .A(wr_en), .ZN(n471) );
  AND2_X1 U32 ( .A1(addr[2]), .A2(n491), .ZN(n315) );
  AND2_X1 U33 ( .A1(addr[3]), .A2(n492), .ZN(n369) );
  AOI222_X1 U34 ( .A1(\mem[9][13] ), .A2(n388), .B1(\mem[11][13] ), .B2(n424), 
        .C1(\mem[10][13] ), .C2(n406), .ZN(n480) );
  AOI222_X1 U35 ( .A1(\mem[9][14] ), .A2(n388), .B1(\mem[11][14] ), .B2(n424), 
        .C1(\mem[10][14] ), .C2(n406), .ZN(n484) );
  AOI222_X1 U36 ( .A1(\mem[9][15] ), .A2(n388), .B1(\mem[11][15] ), .B2(n424), 
        .C1(\mem[10][15] ), .C2(n406), .ZN(n488) );
  NOR2_X1 U37 ( .A1(addr[2]), .A2(addr[3]), .ZN(n493) );
  NOR2_X1 U38 ( .A1(n471), .A2(addr[2]), .ZN(n370) );
  NOR2_X1 U39 ( .A1(n471), .A2(addr[3]), .ZN(n297) );
  NOR2_X1 U40 ( .A1(addr[0]), .A2(addr[1]), .ZN(n492) );
  NOR2_X1 U41 ( .A1(n476), .A2(addr[1]), .ZN(n491) );
  AND2_X1 U42 ( .A1(addr[2]), .A2(n492), .ZN(n296) );
  AND2_X1 U43 ( .A1(addr[2]), .A2(n490), .ZN(n351) );
  AND2_X1 U44 ( .A1(addr[3]), .A2(n489), .ZN(n406) );
  AND2_X1 U45 ( .A1(addr[2]), .A2(n489), .ZN(n333) );
  AND2_X1 U46 ( .A1(addr[3]), .A2(n490), .ZN(n424) );
  AND2_X1 U47 ( .A1(addr[3]), .A2(n491), .ZN(n388) );
  NAND4_X1 U48 ( .A1(n477), .A2(n478), .A3(n479), .A4(n480), .ZN(N56) );
  AOI222_X1 U49 ( .A1(\mem[6][13] ), .A2(n333), .B1(\mem[8][13] ), .B2(n369), 
        .C1(\mem[7][13] ), .C2(n351), .ZN(n479) );
  AOI222_X1 U50 ( .A1(\mem[3][13] ), .A2(n278), .B1(\mem[5][13] ), .B2(n315), 
        .C1(\mem[4][13] ), .C2(n296), .ZN(n478) );
  AOI222_X1 U51 ( .A1(\mem[0][13] ), .A2(n224), .B1(\mem[2][13] ), .B2(n260), 
        .C1(\mem[1][13] ), .C2(n242), .ZN(n477) );
  NAND4_X1 U52 ( .A1(n481), .A2(n482), .A3(n483), .A4(n484), .ZN(N55) );
  AOI222_X1 U53 ( .A1(\mem[6][14] ), .A2(n333), .B1(\mem[8][14] ), .B2(n369), 
        .C1(\mem[7][14] ), .C2(n351), .ZN(n483) );
  AOI222_X1 U54 ( .A1(\mem[3][14] ), .A2(n278), .B1(\mem[5][14] ), .B2(n315), 
        .C1(\mem[4][14] ), .C2(n296), .ZN(n482) );
  AOI222_X1 U55 ( .A1(\mem[0][14] ), .A2(n224), .B1(\mem[2][14] ), .B2(n260), 
        .C1(\mem[1][14] ), .C2(n242), .ZN(n481) );
  NAND4_X1 U56 ( .A1(n485), .A2(n486), .A3(n487), .A4(n488), .ZN(N54) );
  AOI222_X1 U57 ( .A1(\mem[6][15] ), .A2(n333), .B1(\mem[8][15] ), .B2(n369), 
        .C1(\mem[7][15] ), .C2(n351), .ZN(n487) );
  AOI222_X1 U58 ( .A1(\mem[3][15] ), .A2(n278), .B1(\mem[5][15] ), .B2(n315), 
        .C1(\mem[4][15] ), .C2(n296), .ZN(n486) );
  AOI222_X1 U59 ( .A1(\mem[0][15] ), .A2(n224), .B1(\mem[2][15] ), .B2(n260), 
        .C1(\mem[1][15] ), .C2(n242), .ZN(n485) );
  AND2_X1 U60 ( .A1(addr[1]), .A2(addr[0]), .ZN(n490) );
  AND2_X1 U61 ( .A1(addr[1]), .A2(n476), .ZN(n489) );
  INV_X1 U62 ( .A(addr[0]), .ZN(n476) );
  INV_X1 U63 ( .A(n352), .ZN(n454) );
  AOI22_X1 U64 ( .A1(data_in[0]), .A2(n470), .B1(n353), .B2(\mem[8][0] ), .ZN(
        n352) );
  INV_X1 U65 ( .A(n354), .ZN(n442) );
  AOI22_X1 U66 ( .A1(data_in[1]), .A2(n470), .B1(n353), .B2(\mem[8][1] ), .ZN(
        n354) );
  INV_X1 U67 ( .A(n355), .ZN(n430) );
  AOI22_X1 U68 ( .A1(data_in[2]), .A2(n470), .B1(n353), .B2(\mem[8][2] ), .ZN(
        n355) );
  INV_X1 U69 ( .A(n356), .ZN(n200) );
  AOI22_X1 U70 ( .A1(data_in[3]), .A2(n470), .B1(n353), .B2(\mem[8][3] ), .ZN(
        n356) );
  INV_X1 U71 ( .A(n357), .ZN(n188) );
  AOI22_X1 U72 ( .A1(data_in[4]), .A2(n470), .B1(n353), .B2(\mem[8][4] ), .ZN(
        n357) );
  INV_X1 U73 ( .A(n358), .ZN(n176) );
  AOI22_X1 U74 ( .A1(data_in[5]), .A2(n470), .B1(n353), .B2(\mem[8][5] ), .ZN(
        n358) );
  INV_X1 U75 ( .A(n359), .ZN(n164) );
  AOI22_X1 U76 ( .A1(data_in[6]), .A2(n470), .B1(n353), .B2(\mem[8][6] ), .ZN(
        n359) );
  INV_X1 U77 ( .A(n360), .ZN(n152) );
  AOI22_X1 U78 ( .A1(data_in[7]), .A2(n470), .B1(n353), .B2(\mem[8][7] ), .ZN(
        n360) );
  INV_X1 U79 ( .A(n361), .ZN(n140) );
  AOI22_X1 U80 ( .A1(data_in[8]), .A2(n470), .B1(n353), .B2(\mem[8][8] ), .ZN(
        n361) );
  INV_X1 U81 ( .A(n362), .ZN(n128) );
  AOI22_X1 U82 ( .A1(data_in[9]), .A2(n470), .B1(n353), .B2(\mem[8][9] ), .ZN(
        n362) );
  INV_X1 U83 ( .A(n363), .ZN(n116) );
  AOI22_X1 U84 ( .A1(data_in[10]), .A2(n470), .B1(n353), .B2(\mem[8][10] ), 
        .ZN(n363) );
  INV_X1 U85 ( .A(n364), .ZN(n104) );
  AOI22_X1 U86 ( .A1(data_in[11]), .A2(n470), .B1(n353), .B2(\mem[8][11] ), 
        .ZN(n364) );
  INV_X1 U87 ( .A(n365), .ZN(n92) );
  AOI22_X1 U88 ( .A1(data_in[12]), .A2(n470), .B1(n353), .B2(\mem[8][12] ), 
        .ZN(n365) );
  INV_X1 U89 ( .A(n366), .ZN(n80) );
  AOI22_X1 U90 ( .A1(data_in[13]), .A2(n470), .B1(n353), .B2(\mem[8][13] ), 
        .ZN(n366) );
  INV_X1 U91 ( .A(n367), .ZN(n68) );
  AOI22_X1 U92 ( .A1(data_in[14]), .A2(n470), .B1(n353), .B2(\mem[8][14] ), 
        .ZN(n367) );
  INV_X1 U93 ( .A(n368), .ZN(n56) );
  AOI22_X1 U94 ( .A1(data_in[15]), .A2(n470), .B1(n353), .B2(\mem[8][15] ), 
        .ZN(n368) );
  INV_X1 U95 ( .A(n371), .ZN(n453) );
  AOI22_X1 U96 ( .A1(data_in[0]), .A2(n469), .B1(n372), .B2(\mem[9][0] ), .ZN(
        n371) );
  INV_X1 U97 ( .A(n373), .ZN(n441) );
  AOI22_X1 U98 ( .A1(data_in[1]), .A2(n469), .B1(n372), .B2(\mem[9][1] ), .ZN(
        n373) );
  INV_X1 U99 ( .A(n374), .ZN(n429) );
  AOI22_X1 U100 ( .A1(data_in[2]), .A2(n469), .B1(n372), .B2(\mem[9][2] ), 
        .ZN(n374) );
  INV_X1 U101 ( .A(n375), .ZN(n199) );
  AOI22_X1 U102 ( .A1(data_in[3]), .A2(n469), .B1(n372), .B2(\mem[9][3] ), 
        .ZN(n375) );
  INV_X1 U103 ( .A(n376), .ZN(n187) );
  AOI22_X1 U104 ( .A1(data_in[4]), .A2(n469), .B1(n372), .B2(\mem[9][4] ), 
        .ZN(n376) );
  INV_X1 U105 ( .A(n377), .ZN(n175) );
  AOI22_X1 U106 ( .A1(data_in[5]), .A2(n469), .B1(n372), .B2(\mem[9][5] ), 
        .ZN(n377) );
  INV_X1 U107 ( .A(n378), .ZN(n163) );
  AOI22_X1 U108 ( .A1(data_in[6]), .A2(n469), .B1(n372), .B2(\mem[9][6] ), 
        .ZN(n378) );
  INV_X1 U109 ( .A(n379), .ZN(n151) );
  AOI22_X1 U110 ( .A1(data_in[7]), .A2(n469), .B1(n372), .B2(\mem[9][7] ), 
        .ZN(n379) );
  INV_X1 U111 ( .A(n380), .ZN(n139) );
  AOI22_X1 U112 ( .A1(data_in[8]), .A2(n469), .B1(n372), .B2(\mem[9][8] ), 
        .ZN(n380) );
  INV_X1 U113 ( .A(n381), .ZN(n127) );
  AOI22_X1 U114 ( .A1(data_in[9]), .A2(n469), .B1(n372), .B2(\mem[9][9] ), 
        .ZN(n381) );
  INV_X1 U115 ( .A(n382), .ZN(n115) );
  AOI22_X1 U116 ( .A1(data_in[10]), .A2(n469), .B1(n372), .B2(\mem[9][10] ), 
        .ZN(n382) );
  INV_X1 U117 ( .A(n383), .ZN(n103) );
  AOI22_X1 U118 ( .A1(data_in[11]), .A2(n469), .B1(n372), .B2(\mem[9][11] ), 
        .ZN(n383) );
  INV_X1 U119 ( .A(n384), .ZN(n91) );
  AOI22_X1 U120 ( .A1(data_in[12]), .A2(n469), .B1(n372), .B2(\mem[9][12] ), 
        .ZN(n384) );
  INV_X1 U121 ( .A(n385), .ZN(n79) );
  AOI22_X1 U122 ( .A1(data_in[13]), .A2(n469), .B1(n372), .B2(\mem[9][13] ), 
        .ZN(n385) );
  INV_X1 U123 ( .A(n386), .ZN(n67) );
  AOI22_X1 U124 ( .A1(data_in[14]), .A2(n469), .B1(n372), .B2(\mem[9][14] ), 
        .ZN(n386) );
  INV_X1 U125 ( .A(n387), .ZN(n55) );
  AOI22_X1 U126 ( .A1(data_in[15]), .A2(n469), .B1(n372), .B2(\mem[9][15] ), 
        .ZN(n387) );
  INV_X1 U127 ( .A(n389), .ZN(n452) );
  AOI22_X1 U128 ( .A1(data_in[0]), .A2(n468), .B1(n390), .B2(\mem[10][0] ), 
        .ZN(n389) );
  INV_X1 U129 ( .A(n391), .ZN(n440) );
  AOI22_X1 U130 ( .A1(data_in[1]), .A2(n468), .B1(n390), .B2(\mem[10][1] ), 
        .ZN(n391) );
  INV_X1 U131 ( .A(n392), .ZN(n428) );
  AOI22_X1 U132 ( .A1(data_in[2]), .A2(n468), .B1(n390), .B2(\mem[10][2] ), 
        .ZN(n392) );
  INV_X1 U133 ( .A(n393), .ZN(n198) );
  AOI22_X1 U134 ( .A1(data_in[3]), .A2(n468), .B1(n390), .B2(\mem[10][3] ), 
        .ZN(n393) );
  INV_X1 U135 ( .A(n394), .ZN(n186) );
  AOI22_X1 U136 ( .A1(data_in[4]), .A2(n468), .B1(n390), .B2(\mem[10][4] ), 
        .ZN(n394) );
  INV_X1 U137 ( .A(n395), .ZN(n174) );
  AOI22_X1 U138 ( .A1(data_in[5]), .A2(n468), .B1(n390), .B2(\mem[10][5] ), 
        .ZN(n395) );
  INV_X1 U139 ( .A(n396), .ZN(n162) );
  AOI22_X1 U140 ( .A1(data_in[6]), .A2(n468), .B1(n390), .B2(\mem[10][6] ), 
        .ZN(n396) );
  INV_X1 U141 ( .A(n397), .ZN(n150) );
  AOI22_X1 U142 ( .A1(data_in[7]), .A2(n468), .B1(n390), .B2(\mem[10][7] ), 
        .ZN(n397) );
  INV_X1 U143 ( .A(n398), .ZN(n138) );
  AOI22_X1 U144 ( .A1(data_in[8]), .A2(n468), .B1(n390), .B2(\mem[10][8] ), 
        .ZN(n398) );
  INV_X1 U145 ( .A(n399), .ZN(n126) );
  AOI22_X1 U146 ( .A1(data_in[9]), .A2(n468), .B1(n390), .B2(\mem[10][9] ), 
        .ZN(n399) );
  INV_X1 U147 ( .A(n400), .ZN(n114) );
  AOI22_X1 U148 ( .A1(data_in[10]), .A2(n468), .B1(n390), .B2(\mem[10][10] ), 
        .ZN(n400) );
  INV_X1 U149 ( .A(n401), .ZN(n102) );
  AOI22_X1 U150 ( .A1(data_in[11]), .A2(n468), .B1(n390), .B2(\mem[10][11] ), 
        .ZN(n401) );
  INV_X1 U151 ( .A(n402), .ZN(n90) );
  AOI22_X1 U152 ( .A1(data_in[12]), .A2(n468), .B1(n390), .B2(\mem[10][12] ), 
        .ZN(n402) );
  INV_X1 U153 ( .A(n403), .ZN(n78) );
  AOI22_X1 U154 ( .A1(data_in[13]), .A2(n468), .B1(n390), .B2(\mem[10][13] ), 
        .ZN(n403) );
  INV_X1 U155 ( .A(n404), .ZN(n66) );
  AOI22_X1 U156 ( .A1(data_in[14]), .A2(n468), .B1(n390), .B2(\mem[10][14] ), 
        .ZN(n404) );
  INV_X1 U157 ( .A(n405), .ZN(n54) );
  AOI22_X1 U158 ( .A1(data_in[15]), .A2(n468), .B1(n390), .B2(\mem[10][15] ), 
        .ZN(n405) );
  INV_X1 U159 ( .A(n407), .ZN(n451) );
  AOI22_X1 U160 ( .A1(data_in[0]), .A2(n467), .B1(n408), .B2(\mem[11][0] ), 
        .ZN(n407) );
  INV_X1 U161 ( .A(n409), .ZN(n439) );
  AOI22_X1 U162 ( .A1(data_in[1]), .A2(n467), .B1(n408), .B2(\mem[11][1] ), 
        .ZN(n409) );
  INV_X1 U163 ( .A(n410), .ZN(n427) );
  AOI22_X1 U164 ( .A1(data_in[2]), .A2(n467), .B1(n408), .B2(\mem[11][2] ), 
        .ZN(n410) );
  INV_X1 U165 ( .A(n411), .ZN(n197) );
  AOI22_X1 U166 ( .A1(data_in[3]), .A2(n467), .B1(n408), .B2(\mem[11][3] ), 
        .ZN(n411) );
  INV_X1 U167 ( .A(n412), .ZN(n185) );
  AOI22_X1 U168 ( .A1(data_in[4]), .A2(n467), .B1(n408), .B2(\mem[11][4] ), 
        .ZN(n412) );
  INV_X1 U169 ( .A(n413), .ZN(n173) );
  AOI22_X1 U170 ( .A1(data_in[5]), .A2(n467), .B1(n408), .B2(\mem[11][5] ), 
        .ZN(n413) );
  INV_X1 U171 ( .A(n414), .ZN(n161) );
  AOI22_X1 U172 ( .A1(data_in[6]), .A2(n467), .B1(n408), .B2(\mem[11][6] ), 
        .ZN(n414) );
  INV_X1 U173 ( .A(n415), .ZN(n149) );
  AOI22_X1 U174 ( .A1(data_in[7]), .A2(n467), .B1(n408), .B2(\mem[11][7] ), 
        .ZN(n415) );
  INV_X1 U175 ( .A(n416), .ZN(n137) );
  AOI22_X1 U176 ( .A1(data_in[8]), .A2(n467), .B1(n408), .B2(\mem[11][8] ), 
        .ZN(n416) );
  INV_X1 U177 ( .A(n417), .ZN(n125) );
  AOI22_X1 U178 ( .A1(data_in[9]), .A2(n467), .B1(n408), .B2(\mem[11][9] ), 
        .ZN(n417) );
  INV_X1 U179 ( .A(n418), .ZN(n113) );
  AOI22_X1 U180 ( .A1(data_in[10]), .A2(n467), .B1(n408), .B2(\mem[11][10] ), 
        .ZN(n418) );
  INV_X1 U181 ( .A(n419), .ZN(n101) );
  AOI22_X1 U182 ( .A1(data_in[11]), .A2(n467), .B1(n408), .B2(\mem[11][11] ), 
        .ZN(n419) );
  INV_X1 U183 ( .A(n420), .ZN(n89) );
  AOI22_X1 U184 ( .A1(data_in[12]), .A2(n467), .B1(n408), .B2(\mem[11][12] ), 
        .ZN(n420) );
  INV_X1 U185 ( .A(n421), .ZN(n77) );
  AOI22_X1 U186 ( .A1(data_in[13]), .A2(n467), .B1(n408), .B2(\mem[11][13] ), 
        .ZN(n421) );
  INV_X1 U187 ( .A(n422), .ZN(n65) );
  AOI22_X1 U188 ( .A1(data_in[14]), .A2(n467), .B1(n408), .B2(\mem[11][14] ), 
        .ZN(n422) );
  INV_X1 U189 ( .A(n423), .ZN(n53) );
  AOI22_X1 U190 ( .A1(data_in[15]), .A2(n467), .B1(n408), .B2(\mem[11][15] ), 
        .ZN(n423) );
  INV_X1 U191 ( .A(n279), .ZN(n458) );
  AOI22_X1 U192 ( .A1(data_in[0]), .A2(n466), .B1(n280), .B2(\mem[4][0] ), 
        .ZN(n279) );
  INV_X1 U193 ( .A(n281), .ZN(n446) );
  AOI22_X1 U194 ( .A1(data_in[1]), .A2(n466), .B1(n280), .B2(\mem[4][1] ), 
        .ZN(n281) );
  INV_X1 U195 ( .A(n282), .ZN(n434) );
  AOI22_X1 U196 ( .A1(data_in[2]), .A2(n466), .B1(n280), .B2(\mem[4][2] ), 
        .ZN(n282) );
  INV_X1 U197 ( .A(n283), .ZN(n204) );
  AOI22_X1 U198 ( .A1(data_in[3]), .A2(n466), .B1(n280), .B2(\mem[4][3] ), 
        .ZN(n283) );
  INV_X1 U199 ( .A(n284), .ZN(n192) );
  AOI22_X1 U200 ( .A1(data_in[4]), .A2(n466), .B1(n280), .B2(\mem[4][4] ), 
        .ZN(n284) );
  INV_X1 U201 ( .A(n285), .ZN(n180) );
  AOI22_X1 U202 ( .A1(data_in[5]), .A2(n466), .B1(n280), .B2(\mem[4][5] ), 
        .ZN(n285) );
  INV_X1 U203 ( .A(n286), .ZN(n168) );
  AOI22_X1 U204 ( .A1(data_in[6]), .A2(n466), .B1(n280), .B2(\mem[4][6] ), 
        .ZN(n286) );
  INV_X1 U205 ( .A(n287), .ZN(n156) );
  AOI22_X1 U206 ( .A1(data_in[7]), .A2(n466), .B1(n280), .B2(\mem[4][7] ), 
        .ZN(n287) );
  INV_X1 U207 ( .A(n288), .ZN(n144) );
  AOI22_X1 U208 ( .A1(data_in[8]), .A2(n466), .B1(n280), .B2(\mem[4][8] ), 
        .ZN(n288) );
  INV_X1 U209 ( .A(n289), .ZN(n132) );
  AOI22_X1 U210 ( .A1(data_in[9]), .A2(n466), .B1(n280), .B2(\mem[4][9] ), 
        .ZN(n289) );
  INV_X1 U211 ( .A(n290), .ZN(n120) );
  AOI22_X1 U212 ( .A1(data_in[10]), .A2(n466), .B1(n280), .B2(\mem[4][10] ), 
        .ZN(n290) );
  INV_X1 U213 ( .A(n291), .ZN(n108) );
  AOI22_X1 U214 ( .A1(data_in[11]), .A2(n466), .B1(n280), .B2(\mem[4][11] ), 
        .ZN(n291) );
  INV_X1 U215 ( .A(n292), .ZN(n96) );
  AOI22_X1 U216 ( .A1(data_in[12]), .A2(n466), .B1(n280), .B2(\mem[4][12] ), 
        .ZN(n292) );
  INV_X1 U217 ( .A(n293), .ZN(n84) );
  AOI22_X1 U218 ( .A1(data_in[13]), .A2(n466), .B1(n280), .B2(\mem[4][13] ), 
        .ZN(n293) );
  INV_X1 U219 ( .A(n294), .ZN(n72) );
  AOI22_X1 U220 ( .A1(data_in[14]), .A2(n466), .B1(n280), .B2(\mem[4][14] ), 
        .ZN(n294) );
  INV_X1 U221 ( .A(n295), .ZN(n60) );
  AOI22_X1 U222 ( .A1(data_in[15]), .A2(n466), .B1(n280), .B2(\mem[4][15] ), 
        .ZN(n295) );
  INV_X1 U223 ( .A(n298), .ZN(n457) );
  AOI22_X1 U224 ( .A1(data_in[0]), .A2(n465), .B1(n299), .B2(\mem[5][0] ), 
        .ZN(n298) );
  INV_X1 U225 ( .A(n300), .ZN(n445) );
  AOI22_X1 U226 ( .A1(data_in[1]), .A2(n465), .B1(n299), .B2(\mem[5][1] ), 
        .ZN(n300) );
  INV_X1 U227 ( .A(n301), .ZN(n433) );
  AOI22_X1 U228 ( .A1(data_in[2]), .A2(n465), .B1(n299), .B2(\mem[5][2] ), 
        .ZN(n301) );
  INV_X1 U229 ( .A(n302), .ZN(n203) );
  AOI22_X1 U230 ( .A1(data_in[3]), .A2(n465), .B1(n299), .B2(\mem[5][3] ), 
        .ZN(n302) );
  INV_X1 U231 ( .A(n303), .ZN(n191) );
  AOI22_X1 U232 ( .A1(data_in[4]), .A2(n465), .B1(n299), .B2(\mem[5][4] ), 
        .ZN(n303) );
  INV_X1 U233 ( .A(n304), .ZN(n179) );
  AOI22_X1 U234 ( .A1(data_in[5]), .A2(n465), .B1(n299), .B2(\mem[5][5] ), 
        .ZN(n304) );
  INV_X1 U235 ( .A(n305), .ZN(n167) );
  AOI22_X1 U236 ( .A1(data_in[6]), .A2(n465), .B1(n299), .B2(\mem[5][6] ), 
        .ZN(n305) );
  INV_X1 U237 ( .A(n306), .ZN(n155) );
  AOI22_X1 U238 ( .A1(data_in[7]), .A2(n465), .B1(n299), .B2(\mem[5][7] ), 
        .ZN(n306) );
  INV_X1 U239 ( .A(n307), .ZN(n143) );
  AOI22_X1 U240 ( .A1(data_in[8]), .A2(n465), .B1(n299), .B2(\mem[5][8] ), 
        .ZN(n307) );
  INV_X1 U241 ( .A(n308), .ZN(n131) );
  AOI22_X1 U242 ( .A1(data_in[9]), .A2(n465), .B1(n299), .B2(\mem[5][9] ), 
        .ZN(n308) );
  INV_X1 U243 ( .A(n309), .ZN(n119) );
  AOI22_X1 U244 ( .A1(data_in[10]), .A2(n465), .B1(n299), .B2(\mem[5][10] ), 
        .ZN(n309) );
  INV_X1 U245 ( .A(n310), .ZN(n107) );
  AOI22_X1 U246 ( .A1(data_in[11]), .A2(n465), .B1(n299), .B2(\mem[5][11] ), 
        .ZN(n310) );
  INV_X1 U247 ( .A(n311), .ZN(n95) );
  AOI22_X1 U248 ( .A1(data_in[12]), .A2(n465), .B1(n299), .B2(\mem[5][12] ), 
        .ZN(n311) );
  INV_X1 U249 ( .A(n312), .ZN(n83) );
  AOI22_X1 U250 ( .A1(data_in[13]), .A2(n465), .B1(n299), .B2(\mem[5][13] ), 
        .ZN(n312) );
  INV_X1 U251 ( .A(n313), .ZN(n71) );
  AOI22_X1 U252 ( .A1(data_in[14]), .A2(n465), .B1(n299), .B2(\mem[5][14] ), 
        .ZN(n313) );
  INV_X1 U253 ( .A(n314), .ZN(n59) );
  AOI22_X1 U254 ( .A1(data_in[15]), .A2(n465), .B1(n299), .B2(\mem[5][15] ), 
        .ZN(n314) );
  INV_X1 U255 ( .A(n316), .ZN(n456) );
  AOI22_X1 U256 ( .A1(data_in[0]), .A2(n464), .B1(n317), .B2(\mem[6][0] ), 
        .ZN(n316) );
  INV_X1 U257 ( .A(n318), .ZN(n444) );
  AOI22_X1 U258 ( .A1(data_in[1]), .A2(n464), .B1(n317), .B2(\mem[6][1] ), 
        .ZN(n318) );
  INV_X1 U259 ( .A(n319), .ZN(n432) );
  AOI22_X1 U260 ( .A1(data_in[2]), .A2(n464), .B1(n317), .B2(\mem[6][2] ), 
        .ZN(n319) );
  INV_X1 U261 ( .A(n320), .ZN(n202) );
  AOI22_X1 U262 ( .A1(data_in[3]), .A2(n464), .B1(n317), .B2(\mem[6][3] ), 
        .ZN(n320) );
  INV_X1 U263 ( .A(n321), .ZN(n190) );
  AOI22_X1 U264 ( .A1(data_in[4]), .A2(n464), .B1(n317), .B2(\mem[6][4] ), 
        .ZN(n321) );
  INV_X1 U265 ( .A(n322), .ZN(n178) );
  AOI22_X1 U266 ( .A1(data_in[5]), .A2(n464), .B1(n317), .B2(\mem[6][5] ), 
        .ZN(n322) );
  INV_X1 U267 ( .A(n323), .ZN(n166) );
  AOI22_X1 U268 ( .A1(data_in[6]), .A2(n464), .B1(n317), .B2(\mem[6][6] ), 
        .ZN(n323) );
  INV_X1 U269 ( .A(n324), .ZN(n154) );
  AOI22_X1 U270 ( .A1(data_in[7]), .A2(n464), .B1(n317), .B2(\mem[6][7] ), 
        .ZN(n324) );
  INV_X1 U271 ( .A(n325), .ZN(n142) );
  AOI22_X1 U272 ( .A1(data_in[8]), .A2(n464), .B1(n317), .B2(\mem[6][8] ), 
        .ZN(n325) );
  INV_X1 U273 ( .A(n326), .ZN(n130) );
  AOI22_X1 U274 ( .A1(data_in[9]), .A2(n464), .B1(n317), .B2(\mem[6][9] ), 
        .ZN(n326) );
  INV_X1 U275 ( .A(n327), .ZN(n118) );
  AOI22_X1 U276 ( .A1(data_in[10]), .A2(n464), .B1(n317), .B2(\mem[6][10] ), 
        .ZN(n327) );
  INV_X1 U277 ( .A(n328), .ZN(n106) );
  AOI22_X1 U278 ( .A1(data_in[11]), .A2(n464), .B1(n317), .B2(\mem[6][11] ), 
        .ZN(n328) );
  INV_X1 U279 ( .A(n329), .ZN(n94) );
  AOI22_X1 U280 ( .A1(data_in[12]), .A2(n464), .B1(n317), .B2(\mem[6][12] ), 
        .ZN(n329) );
  INV_X1 U281 ( .A(n330), .ZN(n82) );
  AOI22_X1 U282 ( .A1(data_in[13]), .A2(n464), .B1(n317), .B2(\mem[6][13] ), 
        .ZN(n330) );
  INV_X1 U283 ( .A(n331), .ZN(n70) );
  AOI22_X1 U284 ( .A1(data_in[14]), .A2(n464), .B1(n317), .B2(\mem[6][14] ), 
        .ZN(n331) );
  INV_X1 U285 ( .A(n332), .ZN(n58) );
  AOI22_X1 U286 ( .A1(data_in[15]), .A2(n464), .B1(n317), .B2(\mem[6][15] ), 
        .ZN(n332) );
  INV_X1 U287 ( .A(n334), .ZN(n455) );
  AOI22_X1 U288 ( .A1(data_in[0]), .A2(n463), .B1(n335), .B2(\mem[7][0] ), 
        .ZN(n334) );
  INV_X1 U289 ( .A(n336), .ZN(n443) );
  AOI22_X1 U290 ( .A1(data_in[1]), .A2(n463), .B1(n335), .B2(\mem[7][1] ), 
        .ZN(n336) );
  INV_X1 U291 ( .A(n337), .ZN(n431) );
  AOI22_X1 U292 ( .A1(data_in[2]), .A2(n463), .B1(n335), .B2(\mem[7][2] ), 
        .ZN(n337) );
  INV_X1 U293 ( .A(n338), .ZN(n201) );
  AOI22_X1 U294 ( .A1(data_in[3]), .A2(n463), .B1(n335), .B2(\mem[7][3] ), 
        .ZN(n338) );
  INV_X1 U295 ( .A(n339), .ZN(n189) );
  AOI22_X1 U296 ( .A1(data_in[4]), .A2(n463), .B1(n335), .B2(\mem[7][4] ), 
        .ZN(n339) );
  INV_X1 U297 ( .A(n340), .ZN(n177) );
  AOI22_X1 U298 ( .A1(data_in[5]), .A2(n463), .B1(n335), .B2(\mem[7][5] ), 
        .ZN(n340) );
  INV_X1 U299 ( .A(n341), .ZN(n165) );
  AOI22_X1 U300 ( .A1(data_in[6]), .A2(n463), .B1(n335), .B2(\mem[7][6] ), 
        .ZN(n341) );
  INV_X1 U301 ( .A(n342), .ZN(n153) );
  AOI22_X1 U302 ( .A1(data_in[7]), .A2(n463), .B1(n335), .B2(\mem[7][7] ), 
        .ZN(n342) );
  INV_X1 U303 ( .A(n343), .ZN(n141) );
  AOI22_X1 U304 ( .A1(data_in[8]), .A2(n463), .B1(n335), .B2(\mem[7][8] ), 
        .ZN(n343) );
  INV_X1 U305 ( .A(n344), .ZN(n129) );
  AOI22_X1 U306 ( .A1(data_in[9]), .A2(n463), .B1(n335), .B2(\mem[7][9] ), 
        .ZN(n344) );
  INV_X1 U307 ( .A(n345), .ZN(n117) );
  AOI22_X1 U308 ( .A1(data_in[10]), .A2(n463), .B1(n335), .B2(\mem[7][10] ), 
        .ZN(n345) );
  INV_X1 U309 ( .A(n346), .ZN(n105) );
  AOI22_X1 U310 ( .A1(data_in[11]), .A2(n463), .B1(n335), .B2(\mem[7][11] ), 
        .ZN(n346) );
  INV_X1 U311 ( .A(n347), .ZN(n93) );
  AOI22_X1 U312 ( .A1(data_in[12]), .A2(n463), .B1(n335), .B2(\mem[7][12] ), 
        .ZN(n347) );
  INV_X1 U313 ( .A(n348), .ZN(n81) );
  AOI22_X1 U314 ( .A1(data_in[13]), .A2(n463), .B1(n335), .B2(\mem[7][13] ), 
        .ZN(n348) );
  INV_X1 U315 ( .A(n349), .ZN(n69) );
  AOI22_X1 U316 ( .A1(data_in[14]), .A2(n463), .B1(n335), .B2(\mem[7][14] ), 
        .ZN(n349) );
  INV_X1 U317 ( .A(n350), .ZN(n57) );
  AOI22_X1 U318 ( .A1(data_in[15]), .A2(n463), .B1(n335), .B2(\mem[7][15] ), 
        .ZN(n350) );
  INV_X1 U319 ( .A(n225), .ZN(n461) );
  AOI22_X1 U320 ( .A1(data_in[0]), .A2(n474), .B1(n226), .B2(\mem[1][0] ), 
        .ZN(n225) );
  INV_X1 U321 ( .A(n227), .ZN(n449) );
  AOI22_X1 U322 ( .A1(data_in[1]), .A2(n474), .B1(n226), .B2(\mem[1][1] ), 
        .ZN(n227) );
  INV_X1 U323 ( .A(n228), .ZN(n437) );
  AOI22_X1 U324 ( .A1(data_in[2]), .A2(n474), .B1(n226), .B2(\mem[1][2] ), 
        .ZN(n228) );
  INV_X1 U325 ( .A(n229), .ZN(n425) );
  AOI22_X1 U326 ( .A1(data_in[3]), .A2(n474), .B1(n226), .B2(\mem[1][3] ), 
        .ZN(n229) );
  INV_X1 U327 ( .A(n230), .ZN(n195) );
  AOI22_X1 U328 ( .A1(data_in[4]), .A2(n474), .B1(n226), .B2(\mem[1][4] ), 
        .ZN(n230) );
  INV_X1 U329 ( .A(n231), .ZN(n183) );
  AOI22_X1 U330 ( .A1(data_in[5]), .A2(n474), .B1(n226), .B2(\mem[1][5] ), 
        .ZN(n231) );
  INV_X1 U331 ( .A(n232), .ZN(n171) );
  AOI22_X1 U332 ( .A1(data_in[6]), .A2(n474), .B1(n226), .B2(\mem[1][6] ), 
        .ZN(n232) );
  INV_X1 U333 ( .A(n233), .ZN(n159) );
  AOI22_X1 U334 ( .A1(data_in[7]), .A2(n474), .B1(n226), .B2(\mem[1][7] ), 
        .ZN(n233) );
  INV_X1 U335 ( .A(n234), .ZN(n147) );
  AOI22_X1 U336 ( .A1(data_in[8]), .A2(n474), .B1(n226), .B2(\mem[1][8] ), 
        .ZN(n234) );
  INV_X1 U337 ( .A(n235), .ZN(n135) );
  AOI22_X1 U338 ( .A1(data_in[9]), .A2(n474), .B1(n226), .B2(\mem[1][9] ), 
        .ZN(n235) );
  INV_X1 U339 ( .A(n236), .ZN(n123) );
  AOI22_X1 U340 ( .A1(data_in[10]), .A2(n474), .B1(n226), .B2(\mem[1][10] ), 
        .ZN(n236) );
  INV_X1 U341 ( .A(n237), .ZN(n111) );
  AOI22_X1 U342 ( .A1(data_in[11]), .A2(n474), .B1(n226), .B2(\mem[1][11] ), 
        .ZN(n237) );
  INV_X1 U343 ( .A(n238), .ZN(n99) );
  AOI22_X1 U344 ( .A1(data_in[12]), .A2(n474), .B1(n226), .B2(\mem[1][12] ), 
        .ZN(n238) );
  INV_X1 U345 ( .A(n239), .ZN(n87) );
  AOI22_X1 U346 ( .A1(data_in[13]), .A2(n474), .B1(n226), .B2(\mem[1][13] ), 
        .ZN(n239) );
  INV_X1 U347 ( .A(n240), .ZN(n75) );
  AOI22_X1 U348 ( .A1(data_in[14]), .A2(n474), .B1(n226), .B2(\mem[1][14] ), 
        .ZN(n240) );
  INV_X1 U349 ( .A(n241), .ZN(n63) );
  AOI22_X1 U350 ( .A1(data_in[15]), .A2(n474), .B1(n226), .B2(\mem[1][15] ), 
        .ZN(n241) );
  INV_X1 U351 ( .A(n243), .ZN(n460) );
  AOI22_X1 U352 ( .A1(data_in[0]), .A2(n473), .B1(n244), .B2(\mem[2][0] ), 
        .ZN(n243) );
  INV_X1 U353 ( .A(n245), .ZN(n448) );
  AOI22_X1 U354 ( .A1(data_in[1]), .A2(n473), .B1(n244), .B2(\mem[2][1] ), 
        .ZN(n245) );
  INV_X1 U355 ( .A(n246), .ZN(n436) );
  AOI22_X1 U356 ( .A1(data_in[2]), .A2(n473), .B1(n244), .B2(\mem[2][2] ), 
        .ZN(n246) );
  INV_X1 U357 ( .A(n247), .ZN(n206) );
  AOI22_X1 U358 ( .A1(data_in[3]), .A2(n473), .B1(n244), .B2(\mem[2][3] ), 
        .ZN(n247) );
  INV_X1 U359 ( .A(n248), .ZN(n194) );
  AOI22_X1 U360 ( .A1(data_in[4]), .A2(n473), .B1(n244), .B2(\mem[2][4] ), 
        .ZN(n248) );
  INV_X1 U361 ( .A(n249), .ZN(n182) );
  AOI22_X1 U362 ( .A1(data_in[5]), .A2(n473), .B1(n244), .B2(\mem[2][5] ), 
        .ZN(n249) );
  INV_X1 U363 ( .A(n250), .ZN(n170) );
  AOI22_X1 U364 ( .A1(data_in[6]), .A2(n473), .B1(n244), .B2(\mem[2][6] ), 
        .ZN(n250) );
  INV_X1 U365 ( .A(n251), .ZN(n158) );
  AOI22_X1 U366 ( .A1(data_in[7]), .A2(n473), .B1(n244), .B2(\mem[2][7] ), 
        .ZN(n251) );
  INV_X1 U367 ( .A(n252), .ZN(n146) );
  AOI22_X1 U368 ( .A1(data_in[8]), .A2(n473), .B1(n244), .B2(\mem[2][8] ), 
        .ZN(n252) );
  INV_X1 U369 ( .A(n253), .ZN(n134) );
  AOI22_X1 U370 ( .A1(data_in[9]), .A2(n473), .B1(n244), .B2(\mem[2][9] ), 
        .ZN(n253) );
  INV_X1 U371 ( .A(n254), .ZN(n122) );
  AOI22_X1 U372 ( .A1(data_in[10]), .A2(n473), .B1(n244), .B2(\mem[2][10] ), 
        .ZN(n254) );
  INV_X1 U373 ( .A(n255), .ZN(n110) );
  AOI22_X1 U374 ( .A1(data_in[11]), .A2(n473), .B1(n244), .B2(\mem[2][11] ), 
        .ZN(n255) );
  INV_X1 U375 ( .A(n256), .ZN(n98) );
  AOI22_X1 U376 ( .A1(data_in[12]), .A2(n473), .B1(n244), .B2(\mem[2][12] ), 
        .ZN(n256) );
  INV_X1 U377 ( .A(n257), .ZN(n86) );
  AOI22_X1 U378 ( .A1(data_in[13]), .A2(n473), .B1(n244), .B2(\mem[2][13] ), 
        .ZN(n257) );
  INV_X1 U379 ( .A(n258), .ZN(n74) );
  AOI22_X1 U380 ( .A1(data_in[14]), .A2(n473), .B1(n244), .B2(\mem[2][14] ), 
        .ZN(n258) );
  INV_X1 U381 ( .A(n259), .ZN(n62) );
  AOI22_X1 U382 ( .A1(data_in[15]), .A2(n473), .B1(n244), .B2(\mem[2][15] ), 
        .ZN(n259) );
  INV_X1 U383 ( .A(n261), .ZN(n459) );
  AOI22_X1 U384 ( .A1(data_in[0]), .A2(n472), .B1(n262), .B2(\mem[3][0] ), 
        .ZN(n261) );
  INV_X1 U385 ( .A(n263), .ZN(n447) );
  AOI22_X1 U386 ( .A1(data_in[1]), .A2(n472), .B1(n262), .B2(\mem[3][1] ), 
        .ZN(n263) );
  INV_X1 U387 ( .A(n264), .ZN(n435) );
  AOI22_X1 U388 ( .A1(data_in[2]), .A2(n472), .B1(n262), .B2(\mem[3][2] ), 
        .ZN(n264) );
  INV_X1 U389 ( .A(n265), .ZN(n205) );
  AOI22_X1 U390 ( .A1(data_in[3]), .A2(n472), .B1(n262), .B2(\mem[3][3] ), 
        .ZN(n265) );
  INV_X1 U391 ( .A(n266), .ZN(n193) );
  AOI22_X1 U392 ( .A1(data_in[4]), .A2(n472), .B1(n262), .B2(\mem[3][4] ), 
        .ZN(n266) );
  INV_X1 U393 ( .A(n267), .ZN(n181) );
  AOI22_X1 U394 ( .A1(data_in[5]), .A2(n472), .B1(n262), .B2(\mem[3][5] ), 
        .ZN(n267) );
  INV_X1 U395 ( .A(n268), .ZN(n169) );
  AOI22_X1 U396 ( .A1(data_in[6]), .A2(n472), .B1(n262), .B2(\mem[3][6] ), 
        .ZN(n268) );
  INV_X1 U397 ( .A(n269), .ZN(n157) );
  AOI22_X1 U398 ( .A1(data_in[7]), .A2(n472), .B1(n262), .B2(\mem[3][7] ), 
        .ZN(n269) );
  INV_X1 U399 ( .A(n270), .ZN(n145) );
  AOI22_X1 U400 ( .A1(data_in[8]), .A2(n472), .B1(n262), .B2(\mem[3][8] ), 
        .ZN(n270) );
  INV_X1 U401 ( .A(n271), .ZN(n133) );
  AOI22_X1 U402 ( .A1(data_in[9]), .A2(n472), .B1(n262), .B2(\mem[3][9] ), 
        .ZN(n271) );
  INV_X1 U403 ( .A(n272), .ZN(n121) );
  AOI22_X1 U404 ( .A1(data_in[10]), .A2(n472), .B1(n262), .B2(\mem[3][10] ), 
        .ZN(n272) );
  INV_X1 U405 ( .A(n273), .ZN(n109) );
  AOI22_X1 U406 ( .A1(data_in[11]), .A2(n472), .B1(n262), .B2(\mem[3][11] ), 
        .ZN(n273) );
  INV_X1 U407 ( .A(n274), .ZN(n97) );
  AOI22_X1 U408 ( .A1(data_in[12]), .A2(n472), .B1(n262), .B2(\mem[3][12] ), 
        .ZN(n274) );
  INV_X1 U409 ( .A(n275), .ZN(n85) );
  AOI22_X1 U410 ( .A1(data_in[13]), .A2(n472), .B1(n262), .B2(\mem[3][13] ), 
        .ZN(n275) );
  INV_X1 U411 ( .A(n276), .ZN(n73) );
  AOI22_X1 U412 ( .A1(data_in[14]), .A2(n472), .B1(n262), .B2(\mem[3][14] ), 
        .ZN(n276) );
  INV_X1 U413 ( .A(n277), .ZN(n61) );
  AOI22_X1 U414 ( .A1(data_in[15]), .A2(n472), .B1(n262), .B2(\mem[3][15] ), 
        .ZN(n277) );
  INV_X1 U415 ( .A(n207), .ZN(n462) );
  AOI22_X1 U416 ( .A1(n475), .A2(data_in[0]), .B1(n208), .B2(\mem[0][0] ), 
        .ZN(n207) );
  INV_X1 U417 ( .A(n209), .ZN(n450) );
  AOI22_X1 U418 ( .A1(n475), .A2(data_in[1]), .B1(n208), .B2(\mem[0][1] ), 
        .ZN(n209) );
  INV_X1 U419 ( .A(n210), .ZN(n438) );
  AOI22_X1 U420 ( .A1(n475), .A2(data_in[2]), .B1(n208), .B2(\mem[0][2] ), 
        .ZN(n210) );
  INV_X1 U421 ( .A(n211), .ZN(n426) );
  AOI22_X1 U422 ( .A1(n475), .A2(data_in[3]), .B1(n208), .B2(\mem[0][3] ), 
        .ZN(n211) );
  INV_X1 U423 ( .A(n212), .ZN(n196) );
  AOI22_X1 U424 ( .A1(n475), .A2(data_in[4]), .B1(n208), .B2(\mem[0][4] ), 
        .ZN(n212) );
  INV_X1 U425 ( .A(n213), .ZN(n184) );
  AOI22_X1 U426 ( .A1(n475), .A2(data_in[5]), .B1(n208), .B2(\mem[0][5] ), 
        .ZN(n213) );
  INV_X1 U427 ( .A(n214), .ZN(n172) );
  AOI22_X1 U428 ( .A1(n475), .A2(data_in[6]), .B1(n208), .B2(\mem[0][6] ), 
        .ZN(n214) );
  INV_X1 U429 ( .A(n215), .ZN(n160) );
  AOI22_X1 U430 ( .A1(n475), .A2(data_in[7]), .B1(n208), .B2(\mem[0][7] ), 
        .ZN(n215) );
  INV_X1 U431 ( .A(n216), .ZN(n148) );
  AOI22_X1 U432 ( .A1(n475), .A2(data_in[8]), .B1(n208), .B2(\mem[0][8] ), 
        .ZN(n216) );
  INV_X1 U433 ( .A(n217), .ZN(n136) );
  AOI22_X1 U434 ( .A1(n475), .A2(data_in[9]), .B1(n208), .B2(\mem[0][9] ), 
        .ZN(n217) );
  INV_X1 U435 ( .A(n218), .ZN(n124) );
  AOI22_X1 U436 ( .A1(n475), .A2(data_in[10]), .B1(n208), .B2(\mem[0][10] ), 
        .ZN(n218) );
  INV_X1 U437 ( .A(n219), .ZN(n112) );
  AOI22_X1 U438 ( .A1(n475), .A2(data_in[11]), .B1(n208), .B2(\mem[0][11] ), 
        .ZN(n219) );
  INV_X1 U439 ( .A(n220), .ZN(n100) );
  AOI22_X1 U440 ( .A1(n475), .A2(data_in[12]), .B1(n208), .B2(\mem[0][12] ), 
        .ZN(n220) );
  INV_X1 U441 ( .A(n221), .ZN(n88) );
  AOI22_X1 U442 ( .A1(n475), .A2(data_in[13]), .B1(n208), .B2(\mem[0][13] ), 
        .ZN(n221) );
  INV_X1 U443 ( .A(n222), .ZN(n76) );
  AOI22_X1 U444 ( .A1(n475), .A2(data_in[14]), .B1(n208), .B2(\mem[0][14] ), 
        .ZN(n222) );
  INV_X1 U445 ( .A(n223), .ZN(n64) );
  AOI22_X1 U446 ( .A1(n475), .A2(data_in[15]), .B1(n208), .B2(\mem[0][15] ), 
        .ZN(n223) );
  AOI222_X1 U447 ( .A1(\mem[1][0] ), .A2(n242), .B1(\mem[0][0] ), .B2(n224), 
        .C1(\mem[2][0] ), .C2(n260), .ZN(n4) );
  AOI222_X1 U448 ( .A1(\mem[4][0] ), .A2(n296), .B1(\mem[3][0] ), .B2(n278), 
        .C1(\mem[5][0] ), .C2(n315), .ZN(n3) );
  AOI222_X1 U449 ( .A1(\mem[7][0] ), .A2(n351), .B1(\mem[6][0] ), .B2(n333), 
        .C1(\mem[8][0] ), .C2(n369), .ZN(n2) );
  AOI222_X1 U450 ( .A1(\mem[10][0] ), .A2(n406), .B1(\mem[9][0] ), .B2(n388), 
        .C1(\mem[11][0] ), .C2(n424), .ZN(n1) );
  NAND4_X1 U451 ( .A1(n4), .A2(n3), .A3(n2), .A4(n1), .ZN(N69) );
  AOI222_X1 U452 ( .A1(\mem[1][1] ), .A2(n242), .B1(\mem[0][1] ), .B2(n224), 
        .C1(\mem[2][1] ), .C2(n260), .ZN(n8) );
  AOI222_X1 U453 ( .A1(\mem[4][1] ), .A2(n296), .B1(\mem[3][1] ), .B2(n278), 
        .C1(\mem[5][1] ), .C2(n315), .ZN(n7) );
  AOI222_X1 U454 ( .A1(\mem[7][1] ), .A2(n351), .B1(\mem[6][1] ), .B2(n333), 
        .C1(\mem[8][1] ), .C2(n369), .ZN(n6) );
  AOI222_X1 U455 ( .A1(\mem[10][1] ), .A2(n406), .B1(\mem[9][1] ), .B2(n388), 
        .C1(\mem[11][1] ), .C2(n424), .ZN(n5) );
  NAND4_X1 U456 ( .A1(n8), .A2(n7), .A3(n6), .A4(n5), .ZN(N68) );
  AOI222_X1 U457 ( .A1(\mem[1][2] ), .A2(n242), .B1(\mem[0][2] ), .B2(n224), 
        .C1(\mem[2][2] ), .C2(n260), .ZN(n12) );
  AOI222_X1 U458 ( .A1(\mem[4][2] ), .A2(n296), .B1(\mem[3][2] ), .B2(n278), 
        .C1(\mem[5][2] ), .C2(n315), .ZN(n11) );
  AOI222_X1 U459 ( .A1(\mem[7][2] ), .A2(n351), .B1(\mem[6][2] ), .B2(n333), 
        .C1(\mem[8][2] ), .C2(n369), .ZN(n10) );
  AOI222_X1 U460 ( .A1(\mem[10][2] ), .A2(n406), .B1(\mem[9][2] ), .B2(n388), 
        .C1(\mem[11][2] ), .C2(n424), .ZN(n9) );
  NAND4_X1 U461 ( .A1(n12), .A2(n11), .A3(n10), .A4(n9), .ZN(N67) );
  AOI222_X1 U462 ( .A1(\mem[1][3] ), .A2(n242), .B1(\mem[0][3] ), .B2(n224), 
        .C1(\mem[2][3] ), .C2(n260), .ZN(n16) );
  AOI222_X1 U463 ( .A1(\mem[4][3] ), .A2(n296), .B1(\mem[3][3] ), .B2(n278), 
        .C1(\mem[5][3] ), .C2(n315), .ZN(n15) );
  AOI222_X1 U464 ( .A1(\mem[7][3] ), .A2(n351), .B1(\mem[6][3] ), .B2(n333), 
        .C1(\mem[8][3] ), .C2(n369), .ZN(n14) );
  AOI222_X1 U465 ( .A1(\mem[10][3] ), .A2(n406), .B1(\mem[9][3] ), .B2(n388), 
        .C1(\mem[11][3] ), .C2(n424), .ZN(n13) );
  NAND4_X1 U466 ( .A1(n16), .A2(n15), .A3(n14), .A4(n13), .ZN(N66) );
  AOI222_X1 U467 ( .A1(\mem[1][4] ), .A2(n242), .B1(\mem[0][4] ), .B2(n224), 
        .C1(\mem[2][4] ), .C2(n260), .ZN(n20) );
  AOI222_X1 U468 ( .A1(\mem[4][4] ), .A2(n296), .B1(\mem[3][4] ), .B2(n278), 
        .C1(\mem[5][4] ), .C2(n315), .ZN(n19) );
  AOI222_X1 U469 ( .A1(\mem[7][4] ), .A2(n351), .B1(\mem[6][4] ), .B2(n333), 
        .C1(\mem[8][4] ), .C2(n369), .ZN(n18) );
  AOI222_X1 U470 ( .A1(\mem[10][4] ), .A2(n406), .B1(\mem[9][4] ), .B2(n388), 
        .C1(\mem[11][4] ), .C2(n424), .ZN(n17) );
  NAND4_X1 U471 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .ZN(N65) );
  AOI222_X1 U472 ( .A1(\mem[1][5] ), .A2(n242), .B1(\mem[0][5] ), .B2(n224), 
        .C1(\mem[2][5] ), .C2(n260), .ZN(n24) );
  AOI222_X1 U473 ( .A1(\mem[4][5] ), .A2(n296), .B1(\mem[3][5] ), .B2(n278), 
        .C1(\mem[5][5] ), .C2(n315), .ZN(n23) );
  AOI222_X1 U474 ( .A1(\mem[7][5] ), .A2(n351), .B1(\mem[6][5] ), .B2(n333), 
        .C1(\mem[8][5] ), .C2(n369), .ZN(n22) );
  AOI222_X1 U475 ( .A1(\mem[10][5] ), .A2(n406), .B1(\mem[9][5] ), .B2(n388), 
        .C1(\mem[11][5] ), .C2(n424), .ZN(n21) );
  NAND4_X1 U476 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(N64) );
  AOI222_X1 U477 ( .A1(\mem[1][6] ), .A2(n242), .B1(\mem[0][6] ), .B2(n224), 
        .C1(\mem[2][6] ), .C2(n260), .ZN(n28) );
  AOI222_X1 U478 ( .A1(\mem[4][6] ), .A2(n296), .B1(\mem[3][6] ), .B2(n278), 
        .C1(\mem[5][6] ), .C2(n315), .ZN(n27) );
  AOI222_X1 U479 ( .A1(\mem[7][6] ), .A2(n351), .B1(\mem[6][6] ), .B2(n333), 
        .C1(\mem[8][6] ), .C2(n369), .ZN(n26) );
  AOI222_X1 U480 ( .A1(\mem[10][6] ), .A2(n406), .B1(\mem[9][6] ), .B2(n388), 
        .C1(\mem[11][6] ), .C2(n424), .ZN(n25) );
  NAND4_X1 U481 ( .A1(n28), .A2(n27), .A3(n26), .A4(n25), .ZN(N63) );
  AOI222_X1 U482 ( .A1(\mem[1][7] ), .A2(n242), .B1(\mem[0][7] ), .B2(n224), 
        .C1(\mem[2][7] ), .C2(n260), .ZN(n32) );
  AOI222_X1 U483 ( .A1(\mem[4][7] ), .A2(n296), .B1(\mem[3][7] ), .B2(n278), 
        .C1(\mem[5][7] ), .C2(n315), .ZN(n31) );
  AOI222_X1 U484 ( .A1(\mem[7][7] ), .A2(n351), .B1(\mem[6][7] ), .B2(n333), 
        .C1(\mem[8][7] ), .C2(n369), .ZN(n30) );
  AOI222_X1 U485 ( .A1(\mem[10][7] ), .A2(n406), .B1(\mem[9][7] ), .B2(n388), 
        .C1(\mem[11][7] ), .C2(n424), .ZN(n29) );
  NAND4_X1 U486 ( .A1(n32), .A2(n31), .A3(n30), .A4(n29), .ZN(N62) );
  AOI222_X1 U487 ( .A1(\mem[1][8] ), .A2(n242), .B1(\mem[0][8] ), .B2(n224), 
        .C1(\mem[2][8] ), .C2(n260), .ZN(n36) );
  AOI222_X1 U488 ( .A1(\mem[4][8] ), .A2(n296), .B1(\mem[3][8] ), .B2(n278), 
        .C1(\mem[5][8] ), .C2(n315), .ZN(n35) );
  AOI222_X1 U489 ( .A1(\mem[7][8] ), .A2(n351), .B1(\mem[6][8] ), .B2(n333), 
        .C1(\mem[8][8] ), .C2(n369), .ZN(n34) );
  AOI222_X1 U490 ( .A1(\mem[10][8] ), .A2(n406), .B1(\mem[9][8] ), .B2(n388), 
        .C1(\mem[11][8] ), .C2(n424), .ZN(n33) );
  NAND4_X1 U491 ( .A1(n36), .A2(n35), .A3(n34), .A4(n33), .ZN(N61) );
  AOI222_X1 U492 ( .A1(\mem[1][9] ), .A2(n242), .B1(\mem[0][9] ), .B2(n224), 
        .C1(\mem[2][9] ), .C2(n260), .ZN(n40) );
  AOI222_X1 U493 ( .A1(\mem[4][9] ), .A2(n296), .B1(\mem[3][9] ), .B2(n278), 
        .C1(\mem[5][9] ), .C2(n315), .ZN(n39) );
  AOI222_X1 U494 ( .A1(\mem[7][9] ), .A2(n351), .B1(\mem[6][9] ), .B2(n333), 
        .C1(\mem[8][9] ), .C2(n369), .ZN(n38) );
  AOI222_X1 U495 ( .A1(\mem[10][9] ), .A2(n406), .B1(\mem[9][9] ), .B2(n388), 
        .C1(\mem[11][9] ), .C2(n424), .ZN(n37) );
  NAND4_X1 U496 ( .A1(n40), .A2(n39), .A3(n38), .A4(n37), .ZN(N60) );
  AOI222_X1 U497 ( .A1(\mem[1][10] ), .A2(n242), .B1(\mem[0][10] ), .B2(n224), 
        .C1(\mem[2][10] ), .C2(n260), .ZN(n44) );
  AOI222_X1 U498 ( .A1(\mem[4][10] ), .A2(n296), .B1(\mem[3][10] ), .B2(n278), 
        .C1(\mem[5][10] ), .C2(n315), .ZN(n43) );
  AOI222_X1 U499 ( .A1(\mem[7][10] ), .A2(n351), .B1(\mem[6][10] ), .B2(n333), 
        .C1(\mem[8][10] ), .C2(n369), .ZN(n42) );
  AOI222_X1 U500 ( .A1(\mem[10][10] ), .A2(n406), .B1(\mem[9][10] ), .B2(n388), 
        .C1(\mem[11][10] ), .C2(n424), .ZN(n41) );
  NAND4_X1 U501 ( .A1(n44), .A2(n43), .A3(n42), .A4(n41), .ZN(N59) );
  AOI222_X1 U502 ( .A1(\mem[1][11] ), .A2(n242), .B1(\mem[0][11] ), .B2(n224), 
        .C1(\mem[2][11] ), .C2(n260), .ZN(n48) );
  AOI222_X1 U503 ( .A1(\mem[4][11] ), .A2(n296), .B1(\mem[3][11] ), .B2(n278), 
        .C1(\mem[5][11] ), .C2(n315), .ZN(n47) );
  AOI222_X1 U504 ( .A1(\mem[7][11] ), .A2(n351), .B1(\mem[6][11] ), .B2(n333), 
        .C1(\mem[8][11] ), .C2(n369), .ZN(n46) );
  AOI222_X1 U505 ( .A1(\mem[10][11] ), .A2(n406), .B1(\mem[9][11] ), .B2(n388), 
        .C1(\mem[11][11] ), .C2(n424), .ZN(n45) );
  NAND4_X1 U506 ( .A1(n48), .A2(n47), .A3(n46), .A4(n45), .ZN(N58) );
  AOI222_X1 U507 ( .A1(\mem[1][12] ), .A2(n242), .B1(\mem[0][12] ), .B2(n224), 
        .C1(\mem[2][12] ), .C2(n260), .ZN(n52) );
  AOI222_X1 U508 ( .A1(\mem[4][12] ), .A2(n296), .B1(\mem[3][12] ), .B2(n278), 
        .C1(\mem[5][12] ), .C2(n315), .ZN(n51) );
  AOI222_X1 U509 ( .A1(\mem[7][12] ), .A2(n351), .B1(\mem[6][12] ), .B2(n333), 
        .C1(\mem[8][12] ), .C2(n369), .ZN(n50) );
  AOI222_X1 U510 ( .A1(\mem[10][12] ), .A2(n406), .B1(\mem[9][12] ), .B2(n388), 
        .C1(\mem[11][12] ), .C2(n424), .ZN(n49) );
  NAND4_X1 U511 ( .A1(n52), .A2(n51), .A3(n50), .A4(n49), .ZN(N57) );
endmodule


module layer3_16_12_16_16_W_rom_0 ( clk, addr, z );
  input [3:0] addr;
  output [15:0] z;
  input clk;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n19, n36, n37, n38,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n13, n14, n15, n16, n17, n18, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n39, n40, n62, n63, n64, n65, n66, n67, n68, n69, n70;

  DFF_X1 \z_reg[15]  ( .D(n61), .CK(clk), .Q(z[15]), .QN(n1) );
  DFF_X1 \z_reg[14]  ( .D(n60), .CK(clk), .Q(z[14]), .QN(n2) );
  DFF_X1 \z_reg[13]  ( .D(n59), .CK(clk), .Q(z[13]), .QN(n3) );
  DFF_X1 \z_reg[12]  ( .D(n58), .CK(clk), .Q(z[12]), .QN(n4) );
  DFF_X1 \z_reg[11]  ( .D(n57), .CK(clk), .Q(z[11]), .QN(n5) );
  DFF_X1 \z_reg[10]  ( .D(n56), .CK(clk), .Q(z[10]), .QN(n6) );
  DFF_X1 \z_reg[9]  ( .D(n55), .CK(clk), .Q(z[9]), .QN(n7) );
  DFF_X1 \z_reg[8]  ( .D(n54), .CK(clk), .Q(z[8]), .QN(n8) );
  DFF_X1 \z_reg[7]  ( .D(n53), .CK(clk), .Q(z[7]), .QN(n9) );
  DFF_X1 \z_reg[6]  ( .D(n52), .CK(clk), .Q(z[6]), .QN(n16) );
  DFF_X1 \z_reg[5]  ( .D(n51), .CK(clk), .Q(z[5]) );
  DFF_X1 \z_reg[4]  ( .D(n50), .CK(clk), .Q(z[4]), .QN(n10) );
  DFF_X1 \z_reg[3]  ( .D(n49), .CK(clk), .Q(z[3]), .QN(n11) );
  DFF_X1 \z_reg[2]  ( .D(n48), .CK(clk), .Q(z[2]) );
  DFF_X1 \z_reg[1]  ( .D(n47), .CK(clk), .Q(z[1]) );
  DFF_X1 \z_reg[0]  ( .D(n46), .CK(clk), .Q(z[0]), .QN(n12) );
  NAND3_X1 U46 ( .A1(n42), .A2(n69), .A3(addr[2]), .ZN(n36) );
  NAND3_X1 U47 ( .A1(n42), .A2(addr[1]), .A3(addr[2]), .ZN(n38) );
  NAND3_X1 U49 ( .A1(n44), .A2(n69), .A3(addr[2]), .ZN(n37) );
  AND2_X1 U3 ( .A1(n28), .A2(n25), .ZN(n13) );
  AND2_X1 U4 ( .A1(addr[3]), .A2(n45), .ZN(n14) );
  AND3_X1 U5 ( .A1(n36), .A2(n41), .A3(n38), .ZN(n15) );
  NAND3_X1 U6 ( .A1(n13), .A2(n29), .A3(n23), .ZN(n19) );
  AND2_X1 U7 ( .A1(n67), .A2(n15), .ZN(n17) );
  NAND2_X1 U8 ( .A1(n43), .A2(n42), .ZN(n41) );
  NOR2_X1 U9 ( .A1(addr[2]), .A2(addr[1]), .ZN(n43) );
  NOR2_X1 U10 ( .A1(addr[3]), .A2(addr[0]), .ZN(n42) );
  NOR2_X1 U11 ( .A1(n68), .A2(addr[3]), .ZN(n44) );
  OAI21_X1 U12 ( .B1(n19), .B2(n4), .A(n17), .ZN(n58) );
  OAI21_X1 U13 ( .B1(n19), .B2(n3), .A(n17), .ZN(n59) );
  OAI21_X1 U14 ( .B1(n19), .B2(n2), .A(n17), .ZN(n60) );
  OAI21_X1 U15 ( .B1(n19), .B2(n1), .A(n17), .ZN(n61) );
  NOR2_X1 U16 ( .A1(n69), .A2(addr[2]), .ZN(n45) );
  INV_X1 U17 ( .A(n43), .ZN(n70) );
  INV_X1 U18 ( .A(addr[1]), .ZN(n69) );
  INV_X1 U19 ( .A(addr[0]), .ZN(n68) );
  NAND2_X1 U20 ( .A1(n14), .A2(n68), .ZN(n28) );
  NAND2_X1 U21 ( .A1(n42), .A2(n45), .ZN(n25) );
  NAND3_X1 U22 ( .A1(addr[3]), .A2(n43), .A3(addr[0]), .ZN(n29) );
  NAND2_X1 U23 ( .A1(n44), .A2(n43), .ZN(n66) );
  NAND2_X1 U24 ( .A1(n14), .A2(addr[0]), .ZN(n33) );
  OAI211_X1 U25 ( .C1(n70), .C2(addr[0]), .A(n66), .B(n33), .ZN(n18) );
  INV_X1 U26 ( .A(n18), .ZN(n67) );
  INV_X1 U27 ( .A(n44), .ZN(n20) );
  OAI21_X1 U28 ( .B1(n20), .B2(n69), .A(n41), .ZN(n21) );
  INV_X1 U29 ( .A(n21), .ZN(n31) );
  NAND3_X1 U30 ( .A1(n37), .A2(n67), .A3(n31), .ZN(n24) );
  INV_X1 U31 ( .A(n36), .ZN(n22) );
  INV_X1 U32 ( .A(n38), .ZN(n63) );
  NOR3_X1 U33 ( .A1(n24), .A2(n22), .A3(n63), .ZN(n23) );
  INV_X1 U34 ( .A(n24), .ZN(n32) );
  OAI211_X1 U35 ( .C1(n12), .C2(n19), .A(n13), .B(n32), .ZN(n46) );
  NAND3_X1 U36 ( .A1(n37), .A2(n36), .A3(n29), .ZN(n62) );
  INV_X1 U37 ( .A(n62), .ZN(n34) );
  INV_X1 U38 ( .A(n19), .ZN(n39) );
  INV_X1 U39 ( .A(n25), .ZN(n26) );
  AOI21_X1 U40 ( .B1(z[1]), .B2(n39), .A(n26), .ZN(n27) );
  NAND3_X1 U41 ( .A1(n34), .A2(n31), .A3(n27), .ZN(n47) );
  INV_X1 U42 ( .A(n28), .ZN(n64) );
  INV_X1 U43 ( .A(n29), .ZN(n35) );
  AOI211_X1 U44 ( .C1(z[2]), .C2(n39), .A(n64), .B(n35), .ZN(n30) );
  NAND4_X1 U45 ( .A1(n38), .A2(n67), .A3(n31), .A4(n30), .ZN(n48) );
  OAI21_X1 U48 ( .B1(n11), .B2(n19), .A(n32), .ZN(n49) );
  OAI211_X1 U50 ( .C1(n10), .C2(n19), .A(n34), .B(n33), .ZN(n50) );
  AOI21_X1 U51 ( .B1(z[5]), .B2(n39), .A(n35), .ZN(n40) );
  NAND3_X1 U52 ( .A1(n13), .A2(n15), .A3(n40), .ZN(n51) );
  NOR3_X1 U53 ( .A1(n64), .A2(n63), .A3(n62), .ZN(n65) );
  OAI211_X1 U54 ( .C1(n19), .C2(n16), .A(n66), .B(n65), .ZN(n52) );
  OAI21_X1 U55 ( .B1(n9), .B2(n19), .A(n17), .ZN(n53) );
  OAI21_X1 U56 ( .B1(n8), .B2(n19), .A(n17), .ZN(n54) );
  OAI21_X1 U57 ( .B1(n7), .B2(n19), .A(n17), .ZN(n55) );
  OAI21_X1 U58 ( .B1(n6), .B2(n19), .A(n17), .ZN(n56) );
  OAI21_X1 U59 ( .B1(n5), .B2(n19), .A(n17), .ZN(n57) );
endmodule


module layer3_16_12_16_16_B_rom_0 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b1;
  assign z[14] = 1'b1;
  assign z[13] = 1'b1;
  assign z[12] = 1'b1;
  assign z[11] = 1'b1;
  assign z[10] = 1'b1;
  assign z[9] = 1'b1;
  assign z[8] = 1'b1;
  assign z[7] = 1'b1;
  assign z[6] = 1'b1;
  assign z[5] = 1'b1;
  assign z[4] = 1'b0;
  assign z[3] = 1'b1;
  assign z[2] = 1'b1;
  assign z[1] = 1'b1;
  assign z[0] = 1'b1;

endmodule


module layer3_16_12_16_16_W_rom_1 ( clk, addr, z );
  input [3:0] addr;
  output [15:0] z;
  input clk;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n26, n27, n31,
         n33, n38, n42, n43, n44, n45, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n28, n29, n30, n32, n34,
         n35, n36, n37, n39, n40, n41, n46, n47, n48, n49, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82;

  DFF_X1 \z_reg[15]  ( .D(n68), .CK(clk), .Q(z[15]), .QN(n1) );
  DFF_X1 \z_reg[14]  ( .D(n67), .CK(clk), .Q(z[14]), .QN(n2) );
  DFF_X1 \z_reg[13]  ( .D(n66), .CK(clk), .Q(z[13]), .QN(n3) );
  DFF_X1 \z_reg[12]  ( .D(n65), .CK(clk), .Q(z[12]), .QN(n4) );
  DFF_X1 \z_reg[11]  ( .D(n64), .CK(clk), .Q(z[11]), .QN(n5) );
  DFF_X1 \z_reg[10]  ( .D(n63), .CK(clk), .Q(z[10]), .QN(n6) );
  DFF_X1 \z_reg[9]  ( .D(n62), .CK(clk), .Q(z[9]), .QN(n7) );
  DFF_X1 \z_reg[8]  ( .D(n61), .CK(clk), .Q(z[8]), .QN(n8) );
  DFF_X1 \z_reg[7]  ( .D(n60), .CK(clk), .Q(z[7]), .QN(n9) );
  DFF_X1 \z_reg[6]  ( .D(n59), .CK(clk), .Q(z[6]) );
  DFF_X1 \z_reg[5]  ( .D(n58), .CK(clk), .Q(z[5]), .QN(n10) );
  DFF_X1 \z_reg[4]  ( .D(n57), .CK(clk), .Q(z[4]), .QN(n11) );
  DFF_X1 \z_reg[3]  ( .D(n56), .CK(clk), .Q(z[3]) );
  DFF_X1 \z_reg[2]  ( .D(n55), .CK(clk), .Q(z[2]), .QN(n12) );
  DFF_X1 \z_reg[1]  ( .D(n54), .CK(clk), .Q(z[1]), .QN(n13) );
  DFF_X1 \z_reg[0]  ( .D(n53), .CK(clk), .Q(z[0]), .QN(n14) );
  NAND3_X1 U57 ( .A1(n82), .A2(n81), .A3(n52), .ZN(n33) );
  AND2_X1 U3 ( .A1(n78), .A2(n23), .ZN(n15) );
  AND4_X1 U4 ( .A1(n38), .A2(n79), .A3(n21), .A4(n25), .ZN(n16) );
  NAND2_X1 U5 ( .A1(n79), .A2(n33), .ZN(n26) );
  NAND2_X1 U6 ( .A1(n51), .A2(n82), .ZN(n38) );
  NAND2_X1 U7 ( .A1(n42), .A2(n52), .ZN(n31) );
  NOR2_X1 U8 ( .A1(addr[3]), .A2(addr[2]), .ZN(n52) );
  NOR2_X1 U9 ( .A1(n81), .A2(addr[0]), .ZN(n42) );
  NOR2_X1 U10 ( .A1(n82), .A2(addr[1]), .ZN(n45) );
  OAI21_X1 U11 ( .B1(n27), .B2(n4), .A(n16), .ZN(n65) );
  OAI21_X1 U12 ( .B1(n27), .B2(n3), .A(n16), .ZN(n66) );
  OAI21_X1 U13 ( .B1(n27), .B2(n2), .A(n16), .ZN(n67) );
  OAI21_X1 U14 ( .B1(n27), .B2(n1), .A(n16), .ZN(n68) );
  NOR2_X1 U15 ( .A1(n80), .A2(addr[2]), .ZN(n50) );
  OR2_X1 U16 ( .A1(n45), .A2(addr[2]), .ZN(n43) );
  AND2_X1 U17 ( .A1(addr[2]), .A2(n80), .ZN(n51) );
  NAND2_X1 U18 ( .A1(addr[1]), .A2(addr[0]), .ZN(n44) );
  INV_X1 U19 ( .A(n45), .ZN(n19) );
  INV_X1 U20 ( .A(n52), .ZN(n30) );
  INV_X1 U21 ( .A(n51), .ZN(n18) );
  INV_X1 U22 ( .A(n42), .ZN(n17) );
  INV_X1 U23 ( .A(addr[0]), .ZN(n82) );
  INV_X1 U24 ( .A(addr[1]), .ZN(n81) );
  NAND3_X1 U25 ( .A1(n50), .A2(n82), .A3(n81), .ZN(n77) );
  OAI221_X1 U26 ( .B1(n19), .B2(n30), .C1(n18), .C2(n17), .A(n77), .ZN(n20) );
  INV_X1 U27 ( .A(n20), .ZN(n79) );
  NAND2_X1 U28 ( .A1(n42), .A2(n50), .ZN(n72) );
  NAND2_X1 U29 ( .A1(n51), .A2(n45), .ZN(n24) );
  NAND2_X1 U30 ( .A1(n72), .A2(n24), .ZN(n41) );
  INV_X1 U31 ( .A(n41), .ZN(n21) );
  NAND2_X1 U32 ( .A1(n45), .A2(n50), .ZN(n25) );
  INV_X1 U33 ( .A(n50), .ZN(n48) );
  OAI21_X1 U34 ( .B1(n44), .B2(n48), .A(n31), .ZN(n22) );
  INV_X1 U35 ( .A(n22), .ZN(n78) );
  INV_X1 U36 ( .A(n44), .ZN(n36) );
  OAI21_X1 U37 ( .B1(n52), .B2(n51), .A(n36), .ZN(n23) );
  NAND3_X1 U38 ( .A1(n33), .A2(n16), .A3(n15), .ZN(n27) );
  INV_X1 U39 ( .A(n24), .ZN(n28) );
  INV_X1 U40 ( .A(n25), .ZN(n73) );
  NOR3_X1 U41 ( .A1(n26), .A2(n28), .A3(n73), .ZN(n29) );
  OAI221_X1 U42 ( .B1(n27), .B2(n14), .C1(n44), .C2(n30), .A(n29), .ZN(n53) );
  INV_X1 U43 ( .A(n26), .ZN(n35) );
  INV_X1 U44 ( .A(n31), .ZN(n32) );
  NOR2_X1 U45 ( .A1(n41), .A2(n32), .ZN(n34) );
  OAI211_X1 U46 ( .C1(n13), .C2(n27), .A(n35), .B(n34), .ZN(n54) );
  AOI21_X1 U47 ( .B1(n51), .B2(n36), .A(n26), .ZN(n37) );
  OAI211_X1 U48 ( .C1(n12), .C2(n27), .A(n31), .B(n37), .ZN(n55) );
  INV_X1 U49 ( .A(n27), .ZN(n75) );
  INV_X1 U50 ( .A(n77), .ZN(n39) );
  AOI21_X1 U51 ( .B1(z[3]), .B2(n75), .A(n39), .ZN(n40) );
  NAND3_X1 U52 ( .A1(n15), .A2(n38), .A3(n40), .ZN(n56) );
  INV_X1 U53 ( .A(n38), .ZN(n46) );
  NOR2_X1 U54 ( .A1(n46), .A2(n41), .ZN(n47) );
  OAI211_X1 U55 ( .C1(n11), .C2(n27), .A(n78), .B(n47), .ZN(n57) );
  INV_X1 U56 ( .A(addr[3]), .ZN(n80) );
  OAI21_X1 U58 ( .B1(n10), .B2(n80), .A(n48), .ZN(n71) );
  INV_X1 U59 ( .A(addr[2]), .ZN(n69) );
  OAI21_X1 U60 ( .B1(n43), .B2(n42), .A(n80), .ZN(n49) );
  OAI21_X1 U61 ( .B1(n10), .B2(n69), .A(n49), .ZN(n70) );
  MUX2_X1 U62 ( .A(n71), .B(n70), .S(n44), .Z(n58) );
  INV_X1 U63 ( .A(n72), .ZN(n74) );
  AOI211_X1 U64 ( .C1(z[6]), .C2(n75), .A(n74), .B(n73), .ZN(n76) );
  NAND4_X1 U65 ( .A1(n78), .A2(n33), .A3(n77), .A4(n76), .ZN(n59) );
  OAI21_X1 U66 ( .B1(n9), .B2(n27), .A(n16), .ZN(n60) );
  OAI21_X1 U67 ( .B1(n8), .B2(n27), .A(n16), .ZN(n61) );
  OAI21_X1 U68 ( .B1(n7), .B2(n27), .A(n16), .ZN(n62) );
  OAI21_X1 U69 ( .B1(n6), .B2(n27), .A(n16), .ZN(n63) );
  OAI21_X1 U70 ( .B1(n5), .B2(n27), .A(n16), .ZN(n64) );
endmodule


module layer3_16_12_16_16_B_rom_1 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b0;
  assign z[14] = 1'b0;
  assign z[13] = 1'b0;
  assign z[12] = 1'b0;
  assign z[11] = 1'b0;
  assign z[10] = 1'b0;
  assign z[9] = 1'b0;
  assign z[8] = 1'b0;
  assign z[7] = 1'b0;
  assign z[6] = 1'b0;
  assign z[5] = 1'b1;
  assign z[4] = 1'b0;
  assign z[3] = 1'b1;
  assign z[2] = 1'b1;
  assign z[1] = 1'b1;
  assign z[0] = 1'b1;

endmodule


module layer3_16_12_16_16_W_rom_2 ( clk, addr, z );
  input [3:0] addr;
  output [15:0] z;
  input clk;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n11, n12, n27, n28, n32, n33, n42,
         n43, n44, n45, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n10, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n29, n30, n31, n34, n35,
         n36, n37, n38, n39, n40, n41, n46, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFF_X1 \z_reg[14]  ( .D(n64), .CK(clk), .Q(z[14]), .QN(n2) );
  DFF_X1 \z_reg[13]  ( .D(n63), .CK(clk), .Q(z[13]), .QN(n3) );
  DFF_X1 \z_reg[12]  ( .D(n62), .CK(clk), .Q(z[12]), .QN(n4) );
  DFF_X1 \z_reg[11]  ( .D(n61), .CK(clk), .Q(z[11]), .QN(n5) );
  DFF_X1 \z_reg[10]  ( .D(n60), .CK(clk), .Q(z[10]), .QN(n6) );
  DFF_X1 \z_reg[9]  ( .D(n59), .CK(clk), .Q(z[9]), .QN(n7) );
  DFF_X1 \z_reg[8]  ( .D(n58), .CK(clk), .Q(z[8]), .QN(n8) );
  DFF_X1 \z_reg[7]  ( .D(n57), .CK(clk), .Q(z[7]), .QN(n9) );
  DFF_X1 \z_reg[6]  ( .D(n80), .CK(clk), .Q(z[6]), .QN(n14) );
  DFF_X1 \z_reg[5]  ( .D(n56), .CK(clk), .Q(z[5]) );
  DFF_X1 \z_reg[4]  ( .D(n55), .CK(clk), .Q(z[4]), .QN(n11) );
  DFF_X1 \z_reg[3]  ( .D(n54), .CK(clk), .Q(z[3]), .QN(n13) );
  DFF_X1 \z_reg[2]  ( .D(n53), .CK(clk), .Q(z[2]), .QN(n12) );
  DFF_X1 \z_reg[1]  ( .D(n52), .CK(clk), .Q(z[1]) );
  DFF_X1 \z_reg[0]  ( .D(n51), .CK(clk), .Q(z[0]) );
  NAND3_X1 U55 ( .A1(n79), .A2(n78), .A3(n47), .ZN(n44) );
  DFF_X1 \z_reg[15]  ( .D(n65), .CK(clk), .Q(z[15]), .QN(n1) );
  AND2_X1 U3 ( .A1(n30), .A2(n73), .ZN(n10) );
  NAND3_X1 U4 ( .A1(n72), .A2(n36), .A3(n29), .ZN(n28) );
  AND4_X1 U5 ( .A1(n42), .A2(n45), .A3(n43), .A4(n77), .ZN(n15) );
  AND3_X1 U6 ( .A1(n44), .A2(n68), .A3(n21), .ZN(n16) );
  AND2_X1 U7 ( .A1(n16), .A2(n26), .ZN(n17) );
  NOR2_X1 U8 ( .A1(n78), .A2(n79), .ZN(n48) );
  NAND2_X1 U9 ( .A1(n33), .A2(n50), .ZN(n43) );
  NAND2_X1 U10 ( .A1(n49), .A2(n33), .ZN(n45) );
  NAND2_X1 U11 ( .A1(n49), .A2(n48), .ZN(n42) );
  NAND2_X1 U12 ( .A1(n32), .A2(n47), .ZN(n27) );
  NOR2_X1 U13 ( .A1(addr[3]), .A2(addr[2]), .ZN(n49) );
  NOR2_X1 U14 ( .A1(n81), .A2(addr[2]), .ZN(n50) );
  NOR2_X1 U15 ( .A1(n78), .A2(addr[0]), .ZN(n32) );
  NOR2_X1 U16 ( .A1(n79), .A2(addr[1]), .ZN(n33) );
  OAI21_X1 U17 ( .B1(n28), .B2(n4), .A(n15), .ZN(n62) );
  OAI21_X1 U18 ( .B1(n28), .B2(n3), .A(n15), .ZN(n63) );
  OAI21_X1 U19 ( .B1(n28), .B2(n2), .A(n15), .ZN(n64) );
  OAI21_X1 U20 ( .B1(n28), .B2(n1), .A(n15), .ZN(n65) );
  AND2_X1 U21 ( .A1(addr[2]), .A2(n81), .ZN(n47) );
  INV_X1 U22 ( .A(n47), .ZN(n23) );
  INV_X1 U23 ( .A(n33), .ZN(n37) );
  OAI21_X1 U24 ( .B1(n23), .B2(n37), .A(n43), .ZN(n18) );
  INV_X1 U25 ( .A(n18), .ZN(n72) );
  INV_X1 U26 ( .A(n48), .ZN(n22) );
  NAND2_X1 U27 ( .A1(n49), .A2(n32), .ZN(n68) );
  INV_X1 U28 ( .A(n42), .ZN(n20) );
  INV_X1 U29 ( .A(n45), .ZN(n46) );
  INV_X1 U30 ( .A(n27), .ZN(n19) );
  NOR3_X1 U31 ( .A1(n20), .A2(n46), .A3(n19), .ZN(n21) );
  INV_X1 U32 ( .A(addr[0]), .ZN(n79) );
  INV_X1 U33 ( .A(addr[1]), .ZN(n78) );
  NAND3_X1 U34 ( .A1(n49), .A2(n79), .A3(n78), .ZN(n26) );
  NAND2_X1 U35 ( .A1(n48), .A2(n50), .ZN(n30) );
  NAND3_X1 U36 ( .A1(n50), .A2(n79), .A3(n78), .ZN(n73) );
  OAI211_X1 U37 ( .C1(n23), .C2(n22), .A(n17), .B(n10), .ZN(n24) );
  INV_X1 U38 ( .A(n24), .ZN(n36) );
  NAND2_X1 U39 ( .A1(n50), .A2(n32), .ZN(n29) );
  INV_X1 U40 ( .A(n28), .ZN(n70) );
  INV_X1 U41 ( .A(n29), .ZN(n76) );
  AOI21_X1 U42 ( .B1(z[0]), .B2(n70), .A(n76), .ZN(n25) );
  NAND3_X1 U43 ( .A1(n10), .A2(n16), .A3(n25), .ZN(n51) );
  NAND3_X1 U44 ( .A1(n43), .A2(n29), .A3(n26), .ZN(n66) );
  INV_X1 U45 ( .A(n66), .ZN(n35) );
  INV_X1 U46 ( .A(n30), .ZN(n31) );
  AOI21_X1 U47 ( .B1(z[1]), .B2(n70), .A(n31), .ZN(n34) );
  NAND3_X1 U48 ( .A1(n35), .A2(n27), .A3(n34), .ZN(n52) );
  OAI21_X1 U49 ( .B1(n12), .B2(n28), .A(n36), .ZN(n53) );
  INV_X1 U50 ( .A(n32), .ZN(n38) );
  NAND2_X1 U51 ( .A1(n38), .A2(n37), .ZN(n41) );
  INV_X1 U52 ( .A(addr[2]), .ZN(n39) );
  NOR2_X1 U53 ( .A1(n13), .A2(n39), .ZN(n40) );
  MUX2_X1 U54 ( .A(n41), .B(n40), .S(addr[3]), .Z(n54) );
  INV_X1 U56 ( .A(n44), .ZN(n74) );
  NOR3_X1 U57 ( .A1(n66), .A2(n46), .A3(n74), .ZN(n67) );
  OAI211_X1 U58 ( .C1(n11), .C2(n28), .A(n73), .B(n67), .ZN(n55) );
  INV_X1 U59 ( .A(n68), .ZN(n69) );
  AOI21_X1 U60 ( .B1(z[5]), .B2(n70), .A(n69), .ZN(n71) );
  NAND3_X1 U61 ( .A1(n72), .A2(n10), .A3(n71), .ZN(n56) );
  OAI211_X1 U62 ( .C1(n28), .C2(n14), .A(n72), .B(n17), .ZN(n80) );
  INV_X1 U63 ( .A(n73), .ZN(n75) );
  NOR3_X1 U64 ( .A1(n76), .A2(n75), .A3(n74), .ZN(n77) );
  OAI21_X1 U65 ( .B1(n9), .B2(n28), .A(n15), .ZN(n57) );
  OAI21_X1 U66 ( .B1(n8), .B2(n28), .A(n15), .ZN(n58) );
  OAI21_X1 U67 ( .B1(n7), .B2(n28), .A(n15), .ZN(n59) );
  OAI21_X1 U68 ( .B1(n6), .B2(n28), .A(n15), .ZN(n60) );
  OAI21_X1 U69 ( .B1(n5), .B2(n28), .A(n15), .ZN(n61) );
  INV_X1 U70 ( .A(addr[3]), .ZN(n81) );
endmodule


module layer3_16_12_16_16_B_rom_2 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b1;
  assign z[14] = 1'b1;
  assign z[13] = 1'b1;
  assign z[12] = 1'b1;
  assign z[11] = 1'b1;
  assign z[10] = 1'b1;
  assign z[9] = 1'b1;
  assign z[8] = 1'b1;
  assign z[7] = 1'b1;
  assign z[6] = 1'b0;
  assign z[5] = 1'b1;
  assign z[4] = 1'b1;
  assign z[3] = 1'b0;
  assign z[2] = 1'b0;
  assign z[1] = 1'b0;
  assign z[0] = 1'b1;

endmodule


module layer3_16_12_16_16_W_rom_3 ( clk, addr, z );
  input [3:0] addr;
  output [15:0] z;
  input clk;
  wire   n11, n24, n42, n43, n44, n48, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n45,
         n46, n47, n49, n50, n51, n52, n65, n66, n67, n68, n69, n70, n71, n72;

  DFF_X1 \z_reg[12]  ( .D(n66), .CK(clk), .Q(z[12]) );
  DFF_X1 \z_reg[11]  ( .D(n67), .CK(clk), .Q(z[11]), .QN(n7) );
  DFF_X1 \z_reg[10]  ( .D(n68), .CK(clk), .Q(z[10]), .QN(n6) );
  DFF_X1 \z_reg[9]  ( .D(n69), .CK(clk), .Q(z[9]), .QN(n5) );
  DFF_X1 \z_reg[8]  ( .D(n70), .CK(clk), .Q(z[8]), .QN(n4) );
  DFF_X1 \z_reg[7]  ( .D(n71), .CK(clk), .Q(z[7]), .QN(n3) );
  DFF_X1 \z_reg[6]  ( .D(n72), .CK(clk), .Q(z[6]), .QN(n2) );
  DFF_X1 \z_reg[5]  ( .D(n64), .CK(clk), .Q(z[5]) );
  DFF_X1 \z_reg[4]  ( .D(n63), .CK(clk), .Q(z[4]), .QN(n11) );
  DFF_X1 \z_reg[3]  ( .D(n62), .CK(clk), .Q(z[3]), .QN(n1) );
  DFF_X1 \z_reg[2]  ( .D(n61), .CK(clk), .Q(z[2]) );
  DFF_X1 \z_reg[1]  ( .D(n60), .CK(clk), .Q(z[1]) );
  DFF_X1 \z_reg[0]  ( .D(n59), .CK(clk), .Q(z[0]) );
  NAND3_X1 U58 ( .A1(n50), .A2(n46), .A3(n57), .ZN(n44) );
  NAND3_X1 U60 ( .A1(addr[1]), .A2(addr[2]), .A3(n58), .ZN(n42) );
  NAND3_X1 U65 ( .A1(n49), .A2(n47), .A3(addr[0]), .ZN(n43) );
  DFF_X1 \z_reg[15]  ( .D(n51), .CK(clk), .Q(z[15]) );
  DFF_X1 \z_reg[14]  ( .D(n52), .CK(clk), .Q(z[14]) );
  DFF_X1 \z_reg[13]  ( .D(n65), .CK(clk), .Q(z[13]) );
  AND2_X1 U3 ( .A1(n22), .A2(n39), .ZN(n8) );
  NOR2_X1 U4 ( .A1(n49), .A2(addr[2]), .ZN(n57) );
  NOR2_X1 U5 ( .A1(n50), .A2(addr[3]), .ZN(n58) );
  AND2_X1 U6 ( .A1(addr[2]), .A2(addr[3]), .ZN(n9) );
  AND2_X1 U7 ( .A1(n57), .A2(addr[3]), .ZN(n10) );
  AND4_X1 U8 ( .A1(n13), .A2(n43), .A3(n23), .A4(n33), .ZN(n12) );
  AND2_X1 U9 ( .A1(n42), .A2(n44), .ZN(n13) );
  OAI21_X1 U10 ( .B1(addr[3]), .B2(addr[2]), .A(n49), .ZN(n24) );
  INV_X1 U11 ( .A(n53), .ZN(n66) );
  AOI21_X1 U12 ( .B1(z[12]), .B2(n45), .A(n48), .ZN(n53) );
  INV_X1 U13 ( .A(n54), .ZN(n65) );
  AOI21_X1 U14 ( .B1(z[13]), .B2(n45), .A(n48), .ZN(n54) );
  INV_X1 U15 ( .A(n55), .ZN(n52) );
  AOI21_X1 U16 ( .B1(z[14]), .B2(n45), .A(n48), .ZN(n55) );
  INV_X1 U17 ( .A(n56), .ZN(n51) );
  AOI21_X1 U18 ( .B1(z[15]), .B2(n45), .A(n48), .ZN(n56) );
  INV_X1 U19 ( .A(addr[0]), .ZN(n50) );
  XOR2_X1 U20 ( .A(n50), .B(n24), .Z(n14) );
  MUX2_X1 U21 ( .A(n14), .B(z[0]), .S(n9), .Z(n59) );
  INV_X1 U22 ( .A(addr[1]), .ZN(n49) );
  NAND2_X1 U23 ( .A1(n50), .A2(n49), .ZN(n18) );
  INV_X1 U24 ( .A(n57), .ZN(n16) );
  INV_X1 U25 ( .A(n58), .ZN(n15) );
  INV_X1 U26 ( .A(addr[3]), .ZN(n46) );
  INV_X1 U27 ( .A(addr[2]), .ZN(n47) );
  INV_X1 U28 ( .A(n18), .ZN(n34) );
  NAND3_X1 U29 ( .A1(n46), .A2(n47), .A3(n34), .ZN(n25) );
  NAND2_X1 U30 ( .A1(n10), .A2(addr[0]), .ZN(n36) );
  OAI211_X1 U31 ( .C1(n16), .C2(n15), .A(n25), .B(n36), .ZN(n29) );
  INV_X1 U32 ( .A(n29), .ZN(n17) );
  OAI211_X1 U33 ( .C1(addr[2]), .C2(n18), .A(n43), .B(n17), .ZN(n19) );
  INV_X1 U34 ( .A(n19), .ZN(n22) );
  NAND3_X1 U35 ( .A1(addr[2]), .A2(n50), .A3(n46), .ZN(n39) );
  NAND3_X1 U36 ( .A1(n58), .A2(addr[2]), .A3(n49), .ZN(n28) );
  NAND3_X1 U37 ( .A1(n8), .A2(n28), .A3(n13), .ZN(n48) );
  NAND2_X1 U38 ( .A1(n10), .A2(n50), .ZN(n33) );
  INV_X1 U39 ( .A(n48), .ZN(n40) );
  NAND2_X1 U40 ( .A1(n33), .A2(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n41), .ZN(n45) );
  INV_X1 U42 ( .A(n33), .ZN(n20) );
  AOI21_X1 U43 ( .B1(z[1]), .B2(n45), .A(n20), .ZN(n21) );
  NAND3_X1 U44 ( .A1(n22), .A2(n44), .A3(n21), .ZN(n60) );
  NAND3_X1 U45 ( .A1(addr[2]), .A2(n46), .A3(n34), .ZN(n23) );
  INV_X1 U46 ( .A(n25), .ZN(n26) );
  AOI21_X1 U47 ( .B1(z[2]), .B2(n45), .A(n26), .ZN(n27) );
  NAND3_X1 U48 ( .A1(n12), .A2(n28), .A3(n27), .ZN(n61) );
  INV_X1 U49 ( .A(n39), .ZN(n31) );
  INV_X1 U50 ( .A(n28), .ZN(n30) );
  NOR3_X1 U51 ( .A1(n31), .A2(n30), .A3(n29), .ZN(n32) );
  OAI211_X1 U52 ( .C1(n41), .C2(n1), .A(n33), .B(n32), .ZN(n62) );
  MUX2_X1 U53 ( .A(n34), .B(n11), .S(n9), .Z(n35) );
  INV_X1 U54 ( .A(n35), .ZN(n63) );
  INV_X1 U55 ( .A(n36), .ZN(n37) );
  AOI21_X1 U56 ( .B1(z[5]), .B2(n45), .A(n37), .ZN(n38) );
  NAND3_X1 U57 ( .A1(n12), .A2(n39), .A3(n38), .ZN(n64) );
  OAI21_X1 U59 ( .B1(n41), .B2(n2), .A(n8), .ZN(n72) );
  OAI21_X1 U61 ( .B1(n41), .B2(n3), .A(n40), .ZN(n71) );
  OAI21_X1 U62 ( .B1(n41), .B2(n4), .A(n40), .ZN(n70) );
  OAI21_X1 U63 ( .B1(n41), .B2(n5), .A(n40), .ZN(n69) );
  OAI21_X1 U64 ( .B1(n41), .B2(n6), .A(n40), .ZN(n68) );
  OAI21_X1 U66 ( .B1(n41), .B2(n7), .A(n40), .ZN(n67) );
endmodule


module layer3_16_12_16_16_B_rom_3 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b1;
  assign z[14] = 1'b1;
  assign z[13] = 1'b1;
  assign z[12] = 1'b1;
  assign z[11] = 1'b1;
  assign z[10] = 1'b1;
  assign z[9] = 1'b1;
  assign z[8] = 1'b1;
  assign z[7] = 1'b1;
  assign z[6] = 1'b1;
  assign z[5] = 1'b0;
  assign z[4] = 1'b0;
  assign z[3] = 1'b0;
  assign z[2] = 1'b1;
  assign z[1] = 1'b1;
  assign z[0] = 1'b1;

endmodule


module layer3_16_12_16_16_W_rom_4 ( clk, addr, z );
  input [3:0] addr;
  output [15:0] z;
  input clk;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n19, n27, n30, n34,
         n36, n37, n38, n43, n45, n46, n47, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n12, n14, n15, n16,
         n17, n18, n20, n21, n22, n23, n24, n25, n26, n28, n29, n31, n32, n33,
         n35, n39, n40, n41, n42, n44, n48, n66, n67, n68, n69, n70, n71, n72;

  DFF_X1 \z_reg[15]  ( .D(n65), .CK(clk), .Q(z[15]), .QN(n1) );
  DFF_X1 \z_reg[14]  ( .D(n64), .CK(clk), .Q(z[14]), .QN(n2) );
  DFF_X1 \z_reg[13]  ( .D(n63), .CK(clk), .Q(z[13]), .QN(n3) );
  DFF_X1 \z_reg[12]  ( .D(n62), .CK(clk), .Q(z[12]), .QN(n4) );
  DFF_X1 \z_reg[11]  ( .D(n61), .CK(clk), .Q(z[11]), .QN(n5) );
  DFF_X1 \z_reg[10]  ( .D(n60), .CK(clk), .Q(z[10]), .QN(n6) );
  DFF_X1 \z_reg[9]  ( .D(n59), .CK(clk), .Q(z[9]), .QN(n7) );
  DFF_X1 \z_reg[8]  ( .D(n58), .CK(clk), .Q(z[8]), .QN(n8) );
  DFF_X1 \z_reg[7]  ( .D(n57), .CK(clk), .Q(z[7]), .QN(n9) );
  DFF_X1 \z_reg[6]  ( .D(n56), .CK(clk), .Q(z[6]) );
  DFF_X1 \z_reg[5]  ( .D(n55), .CK(clk), .Q(z[5]), .QN(n10) );
  DFF_X1 \z_reg[4]  ( .D(n54), .CK(clk), .Q(z[4]), .QN(n11) );
  DFF_X1 \z_reg[3]  ( .D(n53), .CK(clk), .Q(z[3]) );
  DFF_X1 \z_reg[2]  ( .D(n52), .CK(clk), .Q(z[2]) );
  DFF_X1 \z_reg[1]  ( .D(n71), .CK(clk), .Q(z[1]), .QN(n15) );
  DFF_X1 \z_reg[0]  ( .D(n51), .CK(clk), .Q(z[0]), .QN(n13) );
  NAND3_X1 U50 ( .A1(n47), .A2(addr[0]), .A3(addr[3]), .ZN(n38) );
  NAND3_X1 U51 ( .A1(n47), .A2(n72), .A3(addr[3]), .ZN(n34) );
  NAND3_X1 U53 ( .A1(n49), .A2(n70), .A3(addr[2]), .ZN(n36) );
  NAND3_X1 U55 ( .A1(n46), .A2(n72), .A3(addr[3]), .ZN(n27) );
  AND3_X1 U3 ( .A1(n38), .A2(n30), .A3(n18), .ZN(n12) );
  AND4_X1 U4 ( .A1(n50), .A2(n37), .A3(n27), .A4(n28), .ZN(n14) );
  AND2_X1 U5 ( .A1(n36), .A2(n34), .ZN(n16) );
  NAND3_X1 U6 ( .A1(n14), .A2(n12), .A3(n35), .ZN(n19) );
  AND3_X1 U7 ( .A1(n12), .A2(n69), .A3(n16), .ZN(n17) );
  NAND2_X1 U8 ( .A1(n45), .A2(n47), .ZN(n30) );
  NAND2_X1 U9 ( .A1(n46), .A2(n49), .ZN(n37) );
  NOR2_X1 U10 ( .A1(addr[3]), .A2(addr[0]), .ZN(n45) );
  NOR2_X1 U11 ( .A1(n72), .A2(addr[3]), .ZN(n49) );
  NOR2_X1 U12 ( .A1(n70), .A2(addr[2]), .ZN(n47) );
  NOR2_X1 U13 ( .A1(addr[2]), .A2(addr[1]), .ZN(n46) );
  OAI21_X1 U14 ( .B1(n19), .B2(n4), .A(n17), .ZN(n62) );
  OAI21_X1 U15 ( .B1(n19), .B2(n3), .A(n17), .ZN(n63) );
  OAI21_X1 U16 ( .B1(n19), .B2(n2), .A(n17), .ZN(n64) );
  OAI21_X1 U17 ( .B1(n19), .B2(n1), .A(n17), .ZN(n65) );
  OAI21_X1 U18 ( .B1(addr[3]), .B2(addr[2]), .A(addr[1]), .ZN(n43) );
  NAND2_X1 U19 ( .A1(addr[2]), .A2(n45), .ZN(n50) );
  INV_X1 U20 ( .A(addr[0]), .ZN(n72) );
  NAND2_X1 U21 ( .A1(n47), .A2(n49), .ZN(n28) );
  NAND3_X1 U22 ( .A1(n49), .A2(addr[2]), .A3(addr[1]), .ZN(n18) );
  NAND2_X1 U23 ( .A1(n46), .A2(n45), .ZN(n44) );
  NAND3_X1 U24 ( .A1(addr[3]), .A2(n46), .A3(addr[0]), .ZN(n42) );
  NAND3_X1 U25 ( .A1(n44), .A2(n42), .A3(n16), .ZN(n23) );
  INV_X1 U26 ( .A(n23), .ZN(n35) );
  NAND3_X1 U27 ( .A1(n14), .A2(n34), .A3(n18), .ZN(n39) );
  INV_X1 U28 ( .A(n39), .ZN(n20) );
  OAI211_X1 U29 ( .C1(n13), .C2(n19), .A(n20), .B(n30), .ZN(n51) );
  INV_X1 U30 ( .A(addr[1]), .ZN(n70) );
  NAND3_X1 U31 ( .A1(n45), .A2(addr[2]), .A3(n70), .ZN(n69) );
  INV_X1 U32 ( .A(n30), .ZN(n22) );
  INV_X1 U33 ( .A(n27), .ZN(n21) );
  NOR3_X1 U34 ( .A1(n23), .A2(n22), .A3(n21), .ZN(n24) );
  OAI211_X1 U35 ( .C1(n19), .C2(n15), .A(n69), .B(n24), .ZN(n71) );
  INV_X1 U36 ( .A(n19), .ZN(n32) );
  INV_X1 U37 ( .A(n69), .ZN(n31) );
  INV_X1 U38 ( .A(n42), .ZN(n25) );
  AOI211_X1 U39 ( .C1(z[2]), .C2(n32), .A(n31), .B(n25), .ZN(n26) );
  NAND4_X1 U40 ( .A1(n27), .A2(n37), .A3(n12), .A4(n26), .ZN(n52) );
  INV_X1 U41 ( .A(n28), .ZN(n29) );
  AOI211_X1 U42 ( .C1(z[3]), .C2(n32), .A(n31), .B(n29), .ZN(n33) );
  NAND4_X1 U43 ( .A1(n37), .A2(n38), .A3(n35), .A4(n33), .ZN(n53) );
  INV_X1 U44 ( .A(n36), .ZN(n40) );
  NOR2_X1 U45 ( .A1(n40), .A2(n39), .ZN(n41) );
  OAI211_X1 U46 ( .C1(n11), .C2(n19), .A(n42), .B(n41), .ZN(n54) );
  OAI211_X1 U47 ( .C1(n10), .C2(n19), .A(n14), .B(n44), .ZN(n55) );
  XOR2_X1 U48 ( .A(n72), .B(n43), .Z(n68) );
  INV_X1 U49 ( .A(addr[2]), .ZN(n66) );
  INV_X1 U52 ( .A(addr[3]), .ZN(n48) );
  NOR2_X1 U54 ( .A1(n66), .A2(n48), .ZN(n67) );
  MUX2_X1 U56 ( .A(n68), .B(z[6]), .S(n67), .Z(n56) );
  OAI21_X1 U57 ( .B1(n9), .B2(n19), .A(n17), .ZN(n57) );
  OAI21_X1 U58 ( .B1(n8), .B2(n19), .A(n17), .ZN(n58) );
  OAI21_X1 U59 ( .B1(n7), .B2(n19), .A(n17), .ZN(n59) );
  OAI21_X1 U60 ( .B1(n6), .B2(n19), .A(n17), .ZN(n60) );
  OAI21_X1 U61 ( .B1(n5), .B2(n19), .A(n17), .ZN(n61) );
endmodule


module layer3_16_12_16_16_B_rom_4 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b1;
  assign z[14] = 1'b1;
  assign z[13] = 1'b1;
  assign z[12] = 1'b1;
  assign z[11] = 1'b1;
  assign z[10] = 1'b1;
  assign z[9] = 1'b1;
  assign z[8] = 1'b1;
  assign z[7] = 1'b1;
  assign z[6] = 1'b0;
  assign z[5] = 1'b0;
  assign z[4] = 1'b0;
  assign z[3] = 1'b0;
  assign z[2] = 1'b0;
  assign z[1] = 1'b0;
  assign z[0] = 1'b0;

endmodule


module layer3_16_12_16_16_W_rom_5 ( clk, addr, z );
  input [3:0] addr;
  output [15:0] z;
  input clk;
  wire   n10, n33, n41, n42, n43, n47, n49, n54, n55, n56, n57, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n1, n2, n3, n4, n5, n6, n7, n8, n9, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n34, n35, n36, n37, n38, n39, n40,
         n44, n45, n46, n48, n50, n51, n52, n53, n58, n59, n69, n70, n71, n72,
         n73, n74, n75, n76, n77;

  DFF_X1 \z_reg[14]  ( .D(n76), .CK(clk), .Q(z[14]) );
  DFF_X1 \z_reg[13]  ( .D(n75), .CK(clk), .Q(z[13]) );
  DFF_X1 \z_reg[12]  ( .D(n74), .CK(clk), .Q(z[12]) );
  DFF_X1 \z_reg[11]  ( .D(n73), .CK(clk), .Q(z[11]), .QN(n9) );
  DFF_X1 \z_reg[10]  ( .D(n72), .CK(clk), .Q(z[10]), .QN(n8) );
  DFF_X1 \z_reg[9]  ( .D(n71), .CK(clk), .Q(z[9]), .QN(n7) );
  DFF_X1 \z_reg[8]  ( .D(n70), .CK(clk), .Q(z[8]), .QN(n6) );
  DFF_X1 \z_reg[7]  ( .D(n69), .CK(clk), .Q(z[7]), .QN(n5) );
  DFF_X1 \z_reg[6]  ( .D(n68), .CK(clk), .Q(z[6]) );
  DFF_X1 \z_reg[5]  ( .D(n67), .CK(clk), .Q(z[5]), .QN(n4) );
  DFF_X1 \z_reg[4]  ( .D(n66), .CK(clk), .Q(z[4]), .QN(n10) );
  DFF_X1 \z_reg[3]  ( .D(n65), .CK(clk), .Q(z[3]) );
  DFF_X1 \z_reg[2]  ( .D(n64), .CK(clk), .Q(z[2]), .QN(n3) );
  DFF_X1 \z_reg[1]  ( .D(n63), .CK(clk), .Q(z[1]), .QN(n2) );
  DFF_X1 \z_reg[0]  ( .D(n62), .CK(clk), .Q(z[0]) );
  NAND3_X1 U66 ( .A1(n53), .A2(n52), .A3(n47), .ZN(n43) );
  DFF_X1 \z_reg[15]  ( .D(n77), .CK(clk), .Q(z[15]) );
  AND2_X1 U3 ( .A1(n61), .A2(n58), .ZN(n1) );
  NAND3_X1 U4 ( .A1(n35), .A2(n15), .A3(n14), .ZN(n50) );
  NOR2_X1 U5 ( .A1(n59), .A2(n58), .ZN(n41) );
  AND3_X1 U6 ( .A1(n59), .A2(n58), .A3(n42), .ZN(n33) );
  NOR2_X1 U7 ( .A1(n59), .A2(addr[1]), .ZN(n47) );
  NOR3_X1 U8 ( .A1(addr[2]), .A2(addr[3]), .A3(addr[0]), .ZN(n61) );
  NOR2_X1 U9 ( .A1(n53), .A2(addr[3]), .ZN(n42) );
  AND2_X1 U10 ( .A1(n61), .A2(addr[1]), .ZN(n60) );
  INV_X1 U11 ( .A(n54), .ZN(n74) );
  AOI21_X1 U12 ( .B1(n51), .B2(z[12]), .A(n49), .ZN(n54) );
  INV_X1 U13 ( .A(n55), .ZN(n75) );
  AOI21_X1 U14 ( .B1(n51), .B2(z[13]), .A(n49), .ZN(n55) );
  INV_X1 U15 ( .A(n56), .ZN(n76) );
  AOI21_X1 U16 ( .B1(n51), .B2(z[14]), .A(n49), .ZN(n56) );
  INV_X1 U17 ( .A(n57), .ZN(n77) );
  AOI21_X1 U18 ( .B1(n51), .B2(z[15]), .A(n49), .ZN(n57) );
  INV_X1 U19 ( .A(addr[2]), .ZN(n53) );
  NAND2_X1 U20 ( .A1(addr[3]), .A2(n53), .ZN(n46) );
  INV_X1 U21 ( .A(n46), .ZN(n12) );
  INV_X1 U22 ( .A(addr[0]), .ZN(n59) );
  NAND2_X1 U23 ( .A1(addr[1]), .A2(n59), .ZN(n37) );
  INV_X1 U24 ( .A(n37), .ZN(n11) );
  NAND2_X1 U25 ( .A1(n12), .A2(n11), .ZN(n44) );
  INV_X1 U26 ( .A(addr[1]), .ZN(n58) );
  NAND3_X1 U27 ( .A1(n58), .A2(n59), .A3(n12), .ZN(n32) );
  NAND3_X1 U28 ( .A1(n43), .A2(n44), .A3(n32), .ZN(n49) );
  NAND2_X1 U29 ( .A1(n41), .A2(n12), .ZN(n15) );
  NAND2_X1 U30 ( .A1(n15), .A2(n32), .ZN(n28) );
  INV_X1 U31 ( .A(n28), .ZN(n18) );
  OAI21_X1 U32 ( .B1(n47), .B2(addr[1]), .A(n42), .ZN(n35) );
  INV_X1 U33 ( .A(addr[3]), .ZN(n52) );
  NAND3_X1 U34 ( .A1(n41), .A2(n53), .A3(n52), .ZN(n19) );
  INV_X1 U35 ( .A(n19), .ZN(n16) );
  INV_X1 U36 ( .A(n33), .ZN(n13) );
  OAI21_X1 U37 ( .B1(n45), .B2(n46), .A(n13), .ZN(n27) );
  OR3_X1 U38 ( .A1(n16), .A2(n27), .A3(n60), .ZN(n31) );
  NOR3_X1 U39 ( .A1(n1), .A2(n49), .A3(n31), .ZN(n14) );
  INV_X1 U40 ( .A(n50), .ZN(n51) );
  AOI21_X1 U41 ( .B1(z[0]), .B2(n51), .A(n16), .ZN(n17) );
  NAND3_X1 U42 ( .A1(n18), .A2(n44), .A3(n17), .ZN(n62) );
  INV_X1 U43 ( .A(n42), .ZN(n25) );
  INV_X1 U44 ( .A(n32), .ZN(n21) );
  INV_X1 U45 ( .A(n41), .ZN(n20) );
  OAI211_X1 U46 ( .C1(n20), .C2(n25), .A(n43), .B(n19), .ZN(n26) );
  NOR3_X1 U47 ( .A1(n1), .A2(n21), .A3(n26), .ZN(n22) );
  OAI221_X1 U48 ( .B1(n50), .B2(n2), .C1(n58), .C2(n25), .A(n22), .ZN(n63) );
  INV_X1 U49 ( .A(n47), .ZN(n45) );
  INV_X1 U50 ( .A(n44), .ZN(n23) );
  NOR3_X1 U51 ( .A1(n33), .A2(n23), .A3(n1), .ZN(n24) );
  OAI221_X1 U52 ( .B1(n50), .B2(n3), .C1(n25), .C2(n45), .A(n24), .ZN(n64) );
  INV_X1 U53 ( .A(n26), .ZN(n36) );
  INV_X1 U54 ( .A(n27), .ZN(n30) );
  AOI21_X1 U55 ( .B1(z[3]), .B2(n51), .A(n28), .ZN(n29) );
  NAND3_X1 U56 ( .A1(n36), .A2(n30), .A3(n29), .ZN(n65) );
  INV_X1 U57 ( .A(n31), .ZN(n34) );
  OAI211_X1 U58 ( .C1(n10), .C2(n50), .A(n34), .B(n32), .ZN(n66) );
  OAI211_X1 U59 ( .C1(n50), .C2(n4), .A(n36), .B(n35), .ZN(n67) );
  OAI211_X1 U60 ( .C1(n41), .C2(n53), .A(n37), .B(n45), .ZN(n39) );
  NAND2_X1 U61 ( .A1(z[6]), .A2(addr[2]), .ZN(n38) );
  MUX2_X1 U62 ( .A(n39), .B(n38), .S(addr[3]), .Z(n40) );
  OAI211_X1 U63 ( .C1(n46), .C2(n45), .A(n44), .B(n40), .ZN(n68) );
  INV_X1 U64 ( .A(n49), .ZN(n48) );
  OAI21_X1 U65 ( .B1(n50), .B2(n5), .A(n48), .ZN(n69) );
  OAI21_X1 U67 ( .B1(n50), .B2(n6), .A(n48), .ZN(n70) );
  OAI21_X1 U68 ( .B1(n50), .B2(n7), .A(n48), .ZN(n71) );
  OAI21_X1 U69 ( .B1(n50), .B2(n8), .A(n48), .ZN(n72) );
  OAI21_X1 U70 ( .B1(n50), .B2(n9), .A(n48), .ZN(n73) );
endmodule


module layer3_16_12_16_16_B_rom_5 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b1;
  assign z[14] = 1'b1;
  assign z[13] = 1'b1;
  assign z[12] = 1'b1;
  assign z[11] = 1'b1;
  assign z[10] = 1'b1;
  assign z[9] = 1'b1;
  assign z[8] = 1'b1;
  assign z[7] = 1'b1;
  assign z[6] = 1'b0;
  assign z[5] = 1'b0;
  assign z[4] = 1'b1;
  assign z[3] = 1'b1;
  assign z[2] = 1'b1;
  assign z[1] = 1'b0;
  assign z[0] = 1'b1;

endmodule


module layer3_16_12_16_16_W_rom_6 ( clk, addr, z );
  input [3:0] addr;
  output [15:0] z;
  input clk;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n19, n23, n24,
         n25, n33, n34, n36, n37, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n14, n15, n16, n17, n18,
         n20, n21, n22, n26, n27, n28, n29, n30, n31, n32, n35, n38, n39, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69;
  assign z[4] = 1'b1;

  DFF_X1 \z_reg[15]  ( .D(n57), .CK(clk), .Q(z[15]), .QN(n1) );
  DFF_X1 \z_reg[14]  ( .D(n56), .CK(clk), .Q(z[14]), .QN(n2) );
  DFF_X1 \z_reg[13]  ( .D(n55), .CK(clk), .Q(z[13]), .QN(n3) );
  DFF_X1 \z_reg[12]  ( .D(n54), .CK(clk), .Q(z[12]), .QN(n4) );
  DFF_X1 \z_reg[11]  ( .D(n53), .CK(clk), .Q(z[11]), .QN(n5) );
  DFF_X1 \z_reg[10]  ( .D(n52), .CK(clk), .Q(z[10]), .QN(n6) );
  DFF_X1 \z_reg[9]  ( .D(n51), .CK(clk), .Q(z[9]), .QN(n7) );
  DFF_X1 \z_reg[8]  ( .D(n50), .CK(clk), .Q(z[8]), .QN(n8) );
  DFF_X1 \z_reg[7]  ( .D(n49), .CK(clk), .Q(z[7]), .QN(n9) );
  DFF_X1 \z_reg[6]  ( .D(n48), .CK(clk), .Q(z[6]), .QN(n10) );
  DFF_X1 \z_reg[5]  ( .D(n47), .CK(clk), .Q(z[5]), .QN(n11) );
  DFF_X1 \z_reg[3]  ( .D(n46), .CK(clk), .Q(z[3]) );
  DFF_X1 \z_reg[2]  ( .D(n45), .CK(clk), .Q(z[2]), .QN(n14) );
  DFF_X1 \z_reg[1]  ( .D(n44), .CK(clk), .Q(z[1]), .QN(n12) );
  DFF_X1 \z_reg[0]  ( .D(n43), .CK(clk), .Q(z[0]), .QN(n13) );
  NAND3_X1 U45 ( .A1(n42), .A2(n69), .A3(addr[2]), .ZN(n23) );
  NAND3_X1 U46 ( .A1(addr[3]), .A2(addr[1]), .A3(n41), .ZN(n24) );
  NAND3_X1 U47 ( .A1(n42), .A2(addr[0]), .A3(addr[2]), .ZN(n34) );
  AND4_X1 U4 ( .A1(n36), .A2(n33), .A3(n23), .A4(n26), .ZN(n15) );
  AND3_X1 U5 ( .A1(n23), .A2(n25), .A3(n24), .ZN(n16) );
  INV_X1 U6 ( .A(n66), .ZN(n67) );
  NAND3_X1 U7 ( .A1(n34), .A2(n24), .A3(n15), .ZN(n19) );
  NAND2_X1 U8 ( .A1(n42), .A2(n40), .ZN(n25) );
  NAND2_X1 U9 ( .A1(n40), .A2(n68), .ZN(n33) );
  NAND2_X1 U10 ( .A1(n37), .A2(n41), .ZN(n36) );
  NOR2_X1 U11 ( .A1(n69), .A2(addr[2]), .ZN(n40) );
  NOR2_X1 U12 ( .A1(addr[2]), .A2(addr[0]), .ZN(n41) );
  NOR2_X1 U13 ( .A1(addr[3]), .A2(addr[1]), .ZN(n37) );
  NOR2_X1 U14 ( .A1(n68), .A2(addr[3]), .ZN(n42) );
  OAI21_X1 U15 ( .B1(n19), .B2(n4), .A(n67), .ZN(n54) );
  OAI21_X1 U16 ( .B1(n19), .B2(n3), .A(n67), .ZN(n55) );
  OAI21_X1 U17 ( .B1(n19), .B2(n2), .A(n67), .ZN(n56) );
  OAI21_X1 U18 ( .B1(n19), .B2(n1), .A(n67), .ZN(n57) );
  INV_X1 U19 ( .A(addr[0]), .ZN(n69) );
  NAND2_X1 U20 ( .A1(n37), .A2(addr[2]), .ZN(n17) );
  AND2_X1 U21 ( .A1(n34), .A2(n31), .ZN(n61) );
  NAND3_X1 U22 ( .A1(n40), .A2(addr[3]), .A3(addr[1]), .ZN(n27) );
  INV_X1 U23 ( .A(n27), .ZN(n58) );
  INV_X1 U24 ( .A(n40), .ZN(n22) );
  INV_X1 U25 ( .A(n37), .ZN(n21) );
  INV_X1 U26 ( .A(n41), .ZN(n20) );
  INV_X1 U27 ( .A(n42), .ZN(n18) );
  OAI22_X1 U28 ( .A1(n22), .A2(n21), .B1(n20), .B2(n18), .ZN(n32) );
  INV_X1 U29 ( .A(addr[1]), .ZN(n68) );
  NAND3_X1 U30 ( .A1(n41), .A2(addr[3]), .A3(n68), .ZN(n64) );
  NAND3_X1 U31 ( .A1(n25), .A2(n64), .A3(n17), .ZN(n66) );
  NOR3_X1 U32 ( .A1(n58), .A2(n32), .A3(n66), .ZN(n26) );
  OAI211_X1 U33 ( .C1(n13), .C2(n19), .A(n16), .B(n27), .ZN(n43) );
  INV_X1 U34 ( .A(n34), .ZN(n29) );
  INV_X1 U35 ( .A(n32), .ZN(n28) );
  NAND3_X1 U36 ( .A1(n28), .A2(n33), .A3(n64), .ZN(n39) );
  NOR2_X1 U37 ( .A1(n29), .A2(n39), .ZN(n30) );
  OAI211_X1 U38 ( .C1(n12), .C2(n19), .A(n16), .B(n30), .ZN(n44) );
  NAND3_X1 U39 ( .A1(n37), .A2(addr[0]), .A3(addr[2]), .ZN(n31) );
  NAND3_X1 U40 ( .A1(n36), .A2(n24), .A3(n61), .ZN(n63) );
  INV_X1 U41 ( .A(n25), .ZN(n35) );
  NOR3_X1 U42 ( .A1(n63), .A2(n35), .A3(n32), .ZN(n38) );
  OAI211_X1 U43 ( .C1(n19), .C2(n14), .A(n17), .B(n38), .ZN(n45) );
  INV_X1 U44 ( .A(n39), .ZN(n62) );
  INV_X1 U48 ( .A(n19), .ZN(n59) );
  AOI21_X1 U49 ( .B1(z[3]), .B2(n59), .A(n58), .ZN(n60) );
  NAND3_X1 U50 ( .A1(n62), .A2(n61), .A3(n60), .ZN(n46) );
  OAI21_X1 U51 ( .B1(n11), .B2(n19), .A(n15), .ZN(n47) );
  INV_X1 U52 ( .A(n63), .ZN(n65) );
  OAI211_X1 U53 ( .C1(n10), .C2(n19), .A(n65), .B(n64), .ZN(n48) );
  OAI21_X1 U54 ( .B1(n9), .B2(n19), .A(n67), .ZN(n49) );
  OAI21_X1 U55 ( .B1(n8), .B2(n19), .A(n67), .ZN(n50) );
  OAI21_X1 U56 ( .B1(n7), .B2(n19), .A(n67), .ZN(n51) );
  OAI21_X1 U57 ( .B1(n6), .B2(n19), .A(n67), .ZN(n52) );
  OAI21_X1 U58 ( .B1(n5), .B2(n19), .A(n67), .ZN(n53) );
endmodule


module layer3_16_12_16_16_B_rom_6 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b1;
  assign z[14] = 1'b1;
  assign z[13] = 1'b1;
  assign z[12] = 1'b1;
  assign z[11] = 1'b1;
  assign z[10] = 1'b1;
  assign z[9] = 1'b1;
  assign z[8] = 1'b1;
  assign z[7] = 1'b1;
  assign z[6] = 1'b0;
  assign z[5] = 1'b0;
  assign z[4] = 1'b1;
  assign z[3] = 1'b0;
  assign z[2] = 1'b0;
  assign z[1] = 1'b1;
  assign z[0] = 1'b1;

endmodule


module layer3_16_12_16_16_W_rom_7 ( clk, addr, z );
  input [3:0] addr;
  output [15:0] z;
  input clk;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n21, n28, n30,
         n36, n42, n43, n44, n45, n46, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n14, n15, n16, n17, n18, n19,
         n20, n22, n23, n24, n25, n26, n27, n29, n31, n32, n33, n34, n35, n37,
         n38, n39, n40, n41, n47, n64, n65, n66, n67, n68, n69;

  DFF_X1 \z_reg[15]  ( .D(n63), .CK(clk), .Q(z[15]), .QN(n1) );
  DFF_X1 \z_reg[14]  ( .D(n62), .CK(clk), .Q(z[14]), .QN(n2) );
  DFF_X1 \z_reg[13]  ( .D(n61), .CK(clk), .Q(z[13]), .QN(n3) );
  DFF_X1 \z_reg[12]  ( .D(n60), .CK(clk), .Q(z[12]), .QN(n4) );
  DFF_X1 \z_reg[11]  ( .D(n59), .CK(clk), .Q(z[11]), .QN(n5) );
  DFF_X1 \z_reg[10]  ( .D(n58), .CK(clk), .Q(z[10]), .QN(n6) );
  DFF_X1 \z_reg[9]  ( .D(n57), .CK(clk), .Q(z[9]), .QN(n7) );
  DFF_X1 \z_reg[8]  ( .D(n56), .CK(clk), .Q(z[8]), .QN(n8) );
  DFF_X1 \z_reg[7]  ( .D(n55), .CK(clk), .Q(z[7]), .QN(n9) );
  DFF_X1 \z_reg[6]  ( .D(n54), .CK(clk), .Q(z[6]), .QN(n10) );
  DFF_X1 \z_reg[5]  ( .D(n53), .CK(clk), .Q(z[5]) );
  DFF_X1 \z_reg[4]  ( .D(n52), .CK(clk), .Q(z[4]), .QN(n19) );
  DFF_X1 \z_reg[3]  ( .D(n51), .CK(clk), .Q(z[3]), .QN(n11) );
  DFF_X1 \z_reg[2]  ( .D(n50), .CK(clk), .Q(z[2]), .QN(n15) );
  DFF_X1 \z_reg[1]  ( .D(n49), .CK(clk), .Q(z[1]), .QN(n12) );
  NAND3_X1 U48 ( .A1(addr[3]), .A2(n68), .A3(n46), .ZN(n28) );
  NAND3_X1 U50 ( .A1(addr[3]), .A2(n44), .A3(addr[0]), .ZN(n42) );
  NAND3_X1 U52 ( .A1(addr[1]), .A2(addr[2]), .A3(n43), .ZN(n36) );
  DFF_X1 \z_reg[0]  ( .D(n48), .CK(clk), .Q(z[0]), .QN(n13) );
  AND4_X1 U3 ( .A1(n16), .A2(n28), .A3(n39), .A4(n65), .ZN(n14) );
  AND4_X1 U4 ( .A1(n36), .A2(n30), .A3(n38), .A4(n24), .ZN(n16) );
  AND2_X1 U5 ( .A1(addr[2]), .A2(n45), .ZN(n17) );
  AND3_X1 U6 ( .A1(n42), .A2(n28), .A3(n32), .ZN(n18) );
  AND2_X1 U7 ( .A1(n18), .A2(n38), .ZN(n20) );
  NAND4_X1 U8 ( .A1(n14), .A2(n32), .A3(n64), .A4(n66), .ZN(n21) );
  AND3_X1 U9 ( .A1(n66), .A2(n65), .A3(n20), .ZN(n22) );
  NAND2_X1 U10 ( .A1(n43), .A2(n46), .ZN(n30) );
  INV_X1 U11 ( .A(n42), .ZN(n69) );
  NOR2_X1 U12 ( .A1(n67), .A2(addr[2]), .ZN(n46) );
  NOR2_X1 U13 ( .A1(addr[3]), .A2(addr[0]), .ZN(n43) );
  NOR2_X1 U14 ( .A1(addr[2]), .A2(addr[1]), .ZN(n44) );
  NOR2_X1 U15 ( .A1(n68), .A2(addr[3]), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n21), .B2(n4), .A(n22), .ZN(n60) );
  OAI21_X1 U17 ( .B1(n21), .B2(n3), .A(n22), .ZN(n61) );
  OAI21_X1 U18 ( .B1(n21), .B2(n2), .A(n22), .ZN(n62) );
  OAI21_X1 U19 ( .B1(n21), .B2(n1), .A(n22), .ZN(n63) );
  NAND2_X1 U20 ( .A1(n17), .A2(addr[1]), .ZN(n38) );
  NAND2_X1 U21 ( .A1(n46), .A2(n45), .ZN(n31) );
  INV_X1 U22 ( .A(n31), .ZN(n23) );
  AOI211_X1 U23 ( .C1(n44), .C2(n45), .A(n69), .B(n23), .ZN(n24) );
  NAND3_X1 U24 ( .A1(n46), .A2(addr[3]), .A3(addr[0]), .ZN(n39) );
  INV_X1 U25 ( .A(addr[0]), .ZN(n68) );
  NAND3_X1 U26 ( .A1(addr[3]), .A2(n44), .A3(n68), .ZN(n65) );
  INV_X1 U27 ( .A(addr[1]), .ZN(n67) );
  NAND2_X1 U28 ( .A1(n17), .A2(n67), .ZN(n32) );
  NAND3_X1 U29 ( .A1(n43), .A2(addr[2]), .A3(n67), .ZN(n64) );
  NAND2_X1 U30 ( .A1(n43), .A2(n44), .ZN(n66) );
  OAI211_X1 U31 ( .C1(n13), .C2(n21), .A(n18), .B(n65), .ZN(n48) );
  NAND3_X1 U32 ( .A1(n30), .A2(n28), .A3(n64), .ZN(n26) );
  INV_X1 U33 ( .A(n26), .ZN(n25) );
  OAI211_X1 U34 ( .C1(n12), .C2(n21), .A(n25), .B(n65), .ZN(n49) );
  INV_X1 U35 ( .A(n66), .ZN(n35) );
  INV_X1 U36 ( .A(n38), .ZN(n27) );
  NOR3_X1 U37 ( .A1(n35), .A2(n27), .A3(n26), .ZN(n29) );
  OAI211_X1 U38 ( .C1(n21), .C2(n15), .A(n31), .B(n29), .ZN(n50) );
  OAI211_X1 U39 ( .C1(n11), .C2(n21), .A(n16), .B(n32), .ZN(n51) );
  INV_X1 U40 ( .A(n65), .ZN(n34) );
  INV_X1 U41 ( .A(n36), .ZN(n33) );
  NOR3_X1 U42 ( .A1(n35), .A2(n34), .A3(n33), .ZN(n37) );
  OAI211_X1 U43 ( .C1(n21), .C2(n19), .A(n39), .B(n37), .ZN(n52) );
  INV_X1 U44 ( .A(n21), .ZN(n41) );
  INV_X1 U45 ( .A(n39), .ZN(n40) );
  AOI21_X1 U46 ( .B1(z[5]), .B2(n41), .A(n40), .ZN(n47) );
  NAND3_X1 U47 ( .A1(n20), .A2(n64), .A3(n47), .ZN(n53) );
  OAI21_X1 U49 ( .B1(n10), .B2(n21), .A(n14), .ZN(n54) );
  OAI21_X1 U51 ( .B1(n9), .B2(n21), .A(n22), .ZN(n55) );
  OAI21_X1 U53 ( .B1(n8), .B2(n21), .A(n22), .ZN(n56) );
  OAI21_X1 U54 ( .B1(n7), .B2(n21), .A(n22), .ZN(n57) );
  OAI21_X1 U55 ( .B1(n6), .B2(n21), .A(n22), .ZN(n58) );
  OAI21_X1 U56 ( .B1(n5), .B2(n21), .A(n22), .ZN(n59) );
endmodule


module layer3_16_12_16_16_B_rom_7 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b1;
  assign z[14] = 1'b1;
  assign z[13] = 1'b1;
  assign z[12] = 1'b1;
  assign z[11] = 1'b1;
  assign z[10] = 1'b1;
  assign z[9] = 1'b1;
  assign z[8] = 1'b1;
  assign z[7] = 1'b1;
  assign z[6] = 1'b0;
  assign z[5] = 1'b1;
  assign z[4] = 1'b0;
  assign z[3] = 1'b1;
  assign z[2] = 1'b1;
  assign z[1] = 1'b0;
  assign z[0] = 1'b0;

endmodule


module layer3_16_12_16_16_W_rom_8 ( clk, addr, z );
  input [3:0] addr;
  output [15:0] z;
  input clk;
  wire   n50, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n51, n52, n53, n54, n68;

  DFF_X1 \z_reg[15]  ( .D(n45), .CK(clk), .Q(z[15]) );
  DFF_X1 \z_reg[14]  ( .D(n46), .CK(clk), .Q(z[14]) );
  DFF_X1 \z_reg[13]  ( .D(n47), .CK(clk), .Q(z[13]) );
  DFF_X1 \z_reg[12]  ( .D(n48), .CK(clk), .Q(z[12]) );
  DFF_X1 \z_reg[11]  ( .D(n49), .CK(clk), .Q(z[11]), .QN(n8) );
  DFF_X1 \z_reg[10]  ( .D(n51), .CK(clk), .Q(z[10]), .QN(n7) );
  DFF_X1 \z_reg[9]  ( .D(n52), .CK(clk), .Q(z[9]), .QN(n6) );
  DFF_X1 \z_reg[8]  ( .D(n53), .CK(clk), .Q(z[8]), .QN(n5) );
  DFF_X1 \z_reg[7]  ( .D(n54), .CK(clk), .Q(z[7]), .QN(n4) );
  DFF_X1 \z_reg[6]  ( .D(n68), .CK(clk), .Q(z[6]), .QN(n3) );
  DFF_X1 \z_reg[5]  ( .D(n67), .CK(clk), .Q(z[5]) );
  DFF_X1 \z_reg[4]  ( .D(n66), .CK(clk), .Q(z[4]) );
  DFF_X1 \z_reg[3]  ( .D(n65), .CK(clk), .Q(z[3]) );
  DFF_X1 \z_reg[2]  ( .D(n64), .CK(clk), .Q(z[2]), .QN(n2) );
  DFF_X1 \z_reg[1]  ( .D(n63), .CK(clk), .Q(z[1]), .QN(n1) );
  DFF_X1 \z_reg[0]  ( .D(n62), .CK(clk), .Q(z[0]) );
  AND3_X1 U3 ( .A1(n34), .A2(n21), .A3(n35), .ZN(n9) );
  AND2_X1 U4 ( .A1(n59), .A2(n32), .ZN(n10) );
  NOR2_X1 U5 ( .A1(addr[0]), .A2(addr[1]), .ZN(n61) );
  NOR2_X1 U6 ( .A1(n43), .A2(addr[2]), .ZN(n60) );
  NOR2_X1 U7 ( .A1(n44), .A2(addr[3]), .ZN(n59) );
  AND2_X1 U8 ( .A1(addr[1]), .A2(n17), .ZN(n11) );
  INV_X1 U9 ( .A(n55), .ZN(n48) );
  AOI21_X1 U10 ( .B1(z[12]), .B2(n42), .A(n50), .ZN(n55) );
  INV_X1 U11 ( .A(n56), .ZN(n47) );
  AOI21_X1 U12 ( .B1(z[13]), .B2(n42), .A(n50), .ZN(n56) );
  INV_X1 U13 ( .A(n57), .ZN(n46) );
  AOI21_X1 U14 ( .B1(z[14]), .B2(n42), .A(n50), .ZN(n57) );
  INV_X1 U15 ( .A(n58), .ZN(n45) );
  AOI21_X1 U16 ( .B1(z[15]), .B2(n42), .A(n50), .ZN(n58) );
  INV_X1 U17 ( .A(n59), .ZN(n13) );
  INV_X1 U18 ( .A(addr[1]), .ZN(n16) );
  NAND2_X1 U19 ( .A1(addr[0]), .A2(n16), .ZN(n12) );
  NAND2_X1 U20 ( .A1(addr[0]), .A2(addr[1]), .ZN(n23) );
  INV_X1 U21 ( .A(addr[2]), .ZN(n44) );
  INV_X1 U22 ( .A(addr[3]), .ZN(n43) );
  NAND2_X1 U23 ( .A1(n44), .A2(n43), .ZN(n30) );
  INV_X1 U24 ( .A(n12), .ZN(n26) );
  NAND2_X1 U25 ( .A1(n26), .A2(n60), .ZN(n21) );
  OAI221_X1 U26 ( .B1(n13), .B2(n12), .C1(n23), .C2(n30), .A(n21), .ZN(n14) );
  INV_X1 U27 ( .A(n14), .ZN(n39) );
  INV_X1 U28 ( .A(n23), .ZN(n32) );
  INV_X1 U29 ( .A(addr[0]), .ZN(n17) );
  OAI21_X1 U30 ( .B1(n32), .B2(n11), .A(n60), .ZN(n22) );
  INV_X1 U31 ( .A(n30), .ZN(n15) );
  NAND2_X1 U32 ( .A1(n15), .A2(n16), .ZN(n18) );
  NAND3_X1 U33 ( .A1(n39), .A2(n22), .A3(n18), .ZN(n50) );
  NAND2_X1 U34 ( .A1(n11), .A2(n59), .ZN(n38) );
  AOI221_X1 U35 ( .B1(n11), .B2(n15), .C1(n61), .C2(n60), .A(n10), .ZN(n34) );
  INV_X1 U36 ( .A(n50), .ZN(n40) );
  NAND3_X1 U37 ( .A1(n59), .A2(n17), .A3(n16), .ZN(n35) );
  NAND4_X1 U38 ( .A1(n34), .A2(n40), .A3(n35), .A4(n38), .ZN(n41) );
  INV_X1 U39 ( .A(n41), .ZN(n42) );
  INV_X1 U40 ( .A(n18), .ZN(n19) );
  AOI21_X1 U41 ( .B1(z[0]), .B2(n42), .A(n19), .ZN(n20) );
  NAND3_X1 U42 ( .A1(n38), .A2(n21), .A3(n20), .ZN(n62) );
  OAI211_X1 U43 ( .C1(n41), .C2(n1), .A(n9), .B(n22), .ZN(n63) );
  NOR2_X1 U44 ( .A1(z[2]), .A2(n44), .ZN(n28) );
  NOR2_X1 U45 ( .A1(n44), .A2(n2), .ZN(n25) );
  NAND2_X1 U46 ( .A1(n23), .A2(n44), .ZN(n29) );
  INV_X1 U47 ( .A(n29), .ZN(n24) );
  AOI211_X1 U48 ( .C1(n25), .C2(n32), .A(n10), .B(n24), .ZN(n27) );
  OAI33_X1 U49 ( .A1(n28), .A2(n43), .A3(n32), .B1(n27), .B2(n11), .B3(n26), 
        .ZN(n64) );
  NAND3_X1 U50 ( .A1(z[3]), .A2(addr[3]), .A3(addr[2]), .ZN(n31) );
  NAND3_X1 U51 ( .A1(n31), .A2(n30), .A3(n29), .ZN(n65) );
  AOI22_X1 U52 ( .A1(n60), .A2(n32), .B1(z[4]), .B2(n42), .ZN(n33) );
  NAND3_X1 U53 ( .A1(n34), .A2(n38), .A3(n33), .ZN(n66) );
  INV_X1 U54 ( .A(n35), .ZN(n36) );
  AOI21_X1 U55 ( .B1(z[5]), .B2(n42), .A(n36), .ZN(n37) );
  NAND3_X1 U56 ( .A1(n39), .A2(n38), .A3(n37), .ZN(n67) );
  OAI21_X1 U57 ( .B1(n41), .B2(n3), .A(n9), .ZN(n68) );
  OAI21_X1 U58 ( .B1(n41), .B2(n4), .A(n40), .ZN(n54) );
  OAI21_X1 U59 ( .B1(n41), .B2(n5), .A(n40), .ZN(n53) );
  OAI21_X1 U60 ( .B1(n41), .B2(n6), .A(n40), .ZN(n52) );
  OAI21_X1 U61 ( .B1(n41), .B2(n7), .A(n40), .ZN(n51) );
  OAI21_X1 U62 ( .B1(n41), .B2(n8), .A(n40), .ZN(n49) );
endmodule


module layer3_16_12_16_16_B_rom_8 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b1;
  assign z[14] = 1'b1;
  assign z[13] = 1'b1;
  assign z[12] = 1'b1;
  assign z[11] = 1'b1;
  assign z[10] = 1'b1;
  assign z[9] = 1'b1;
  assign z[8] = 1'b1;
  assign z[7] = 1'b1;
  assign z[6] = 1'b1;
  assign z[5] = 1'b0;
  assign z[4] = 1'b0;
  assign z[3] = 1'b1;
  assign z[2] = 1'b1;
  assign z[1] = 1'b1;
  assign z[0] = 1'b0;

endmodule


module layer3_16_12_16_16_W_rom_9 ( clk, addr, z );
  input [3:0] addr;
  output [15:0] z;
  input clk;
  wire   n11, n34, n35, n39, n40, n44, n50, n52, n57, n58, n59, n60, n62, n63,
         n65, n66, n67, n68, n69, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n36, n37, n38, n41, n42, n43, n45,
         n46, n47, n48, n49, n51, n53, n54, n55, n56, n61, n64, n70, n71, n72,
         n73;

  DFF_X1 \z_reg[15]  ( .D(n72), .CK(clk), .Q(z[15]) );
  DFF_X1 \z_reg[14]  ( .D(n71), .CK(clk), .Q(z[14]) );
  DFF_X1 \z_reg[13]  ( .D(n70), .CK(clk), .Q(z[13]) );
  DFF_X1 \z_reg[12]  ( .D(n64), .CK(clk), .Q(z[12]) );
  DFF_X1 \z_reg[11]  ( .D(n61), .CK(clk), .Q(z[11]), .QN(n6) );
  DFF_X1 \z_reg[10]  ( .D(n56), .CK(clk), .Q(z[10]), .QN(n5) );
  DFF_X1 \z_reg[9]  ( .D(n55), .CK(clk), .Q(z[9]), .QN(n4) );
  DFF_X1 \z_reg[8]  ( .D(n54), .CK(clk), .Q(z[8]), .QN(n3) );
  DFF_X1 \z_reg[7]  ( .D(n53), .CK(clk), .Q(z[7]), .QN(n2) );
  DFF_X1 \z_reg[6]  ( .D(n69), .CK(clk), .Q(z[6]) );
  DFF_X1 \z_reg[5]  ( .D(n51), .CK(clk), .Q(z[5]) );
  DFF_X1 \z_reg[4]  ( .D(n68), .CK(clk), .Q(z[4]) );
  DFF_X1 \z_reg[3]  ( .D(n67), .CK(clk), .Q(z[3]) );
  DFF_X1 \z_reg[2]  ( .D(n66), .CK(clk), .Q(z[2]), .QN(n1) );
  DFF_X1 \z_reg[1]  ( .D(n65), .CK(clk), .Q(z[1]), .QN(n11) );
  DFF_X1 \z_reg[0]  ( .D(n49), .CK(clk), .Q(z[0]) );
  NAND3_X1 U65 ( .A1(n63), .A2(n47), .A3(addr[0]), .ZN(n62) );
  NAND3_X1 U66 ( .A1(addr[0]), .A2(n47), .A3(n34), .ZN(n44) );
  NAND3_X1 U67 ( .A1(n48), .A2(n47), .A3(n34), .ZN(n39) );
  NAND3_X1 U69 ( .A1(n63), .A2(n48), .A3(addr[1]), .ZN(n40) );
  AND2_X1 U3 ( .A1(n8), .A2(n27), .ZN(n7) );
  AND2_X1 U4 ( .A1(n50), .A2(n12), .ZN(n8) );
  INV_X1 U5 ( .A(n39), .ZN(n73) );
  NAND2_X1 U6 ( .A1(n45), .A2(n47), .ZN(n50) );
  AND3_X1 U7 ( .A1(n50), .A2(n40), .A3(n27), .ZN(n9) );
  NAND2_X1 U8 ( .A1(n48), .A2(n47), .ZN(n35) );
  NOR2_X1 U9 ( .A1(n46), .A2(addr[2]), .ZN(n34) );
  NOR2_X1 U10 ( .A1(addr[3]), .A2(addr[2]), .ZN(n63) );
  AND2_X1 U11 ( .A1(addr[2]), .A2(n46), .ZN(n10) );
  INV_X1 U12 ( .A(n57), .ZN(n64) );
  AOI21_X1 U13 ( .B1(n43), .B2(z[12]), .A(n52), .ZN(n57) );
  INV_X1 U14 ( .A(n58), .ZN(n70) );
  AOI21_X1 U15 ( .B1(n43), .B2(z[13]), .A(n52), .ZN(n58) );
  INV_X1 U16 ( .A(n59), .ZN(n71) );
  AOI21_X1 U17 ( .B1(n43), .B2(z[14]), .A(n52), .ZN(n59) );
  INV_X1 U18 ( .A(n60), .ZN(n72) );
  AOI21_X1 U19 ( .B1(n43), .B2(z[15]), .A(n52), .ZN(n60) );
  INV_X1 U20 ( .A(addr[1]), .ZN(n47) );
  INV_X1 U21 ( .A(addr[3]), .ZN(n46) );
  INV_X1 U22 ( .A(addr[0]), .ZN(n48) );
  NAND2_X1 U23 ( .A1(n10), .A2(n48), .ZN(n42) );
  NAND2_X1 U24 ( .A1(addr[0]), .A2(addr[1]), .ZN(n19) );
  INV_X1 U25 ( .A(n19), .ZN(n24) );
  NAND2_X1 U26 ( .A1(n34), .A2(n24), .ZN(n29) );
  OAI21_X1 U27 ( .B1(n47), .B2(n42), .A(n29), .ZN(n16) );
  INV_X1 U28 ( .A(n16), .ZN(n12) );
  NAND2_X1 U29 ( .A1(n63), .A2(n24), .ZN(n27) );
  NAND3_X1 U30 ( .A1(n34), .A2(addr[1]), .A3(n48), .ZN(n32) );
  NAND2_X1 U31 ( .A1(n7), .A2(n32), .ZN(n52) );
  INV_X1 U32 ( .A(n52), .ZN(n38) );
  NAND3_X1 U33 ( .A1(n63), .A2(n47), .A3(n48), .ZN(n13) );
  NAND2_X1 U34 ( .A1(n44), .A2(n13), .ZN(n28) );
  NOR3_X1 U35 ( .A1(n73), .A2(n10), .A3(n28), .ZN(n14) );
  NAND4_X1 U36 ( .A1(n40), .A2(n62), .A3(n38), .A4(n14), .ZN(n41) );
  INV_X1 U37 ( .A(n41), .ZN(n43) );
  NAND3_X1 U38 ( .A1(n39), .A2(n40), .A3(n8), .ZN(n23) );
  AOI21_X1 U39 ( .B1(z[0]), .B2(n43), .A(n23), .ZN(n15) );
  NAND3_X1 U40 ( .A1(n44), .A2(n62), .A3(n15), .ZN(n49) );
  OAI21_X1 U41 ( .B1(n11), .B2(n41), .A(n7), .ZN(n65) );
  INV_X1 U42 ( .A(n27), .ZN(n17) );
  NOR3_X1 U43 ( .A1(n17), .A2(n16), .A3(n28), .ZN(n18) );
  OAI211_X1 U44 ( .C1(n41), .C2(n1), .A(n32), .B(n18), .ZN(n66) );
  NAND3_X1 U45 ( .A1(z[3]), .A2(addr[3]), .A3(addr[2]), .ZN(n22) );
  MUX2_X1 U46 ( .A(n46), .B(n34), .S(n35), .Z(n20) );
  OAI21_X1 U47 ( .B1(n10), .B2(n20), .A(n19), .ZN(n21) );
  NAND2_X1 U48 ( .A1(n22), .A2(n21), .ZN(n67) );
  INV_X1 U49 ( .A(n23), .ZN(n26) );
  AOI22_X1 U50 ( .A1(n24), .A2(n10), .B1(z[4]), .B2(n43), .ZN(n25) );
  NAND3_X1 U51 ( .A1(n26), .A2(n32), .A3(n25), .ZN(n68) );
  INV_X1 U52 ( .A(n28), .ZN(n37) );
  INV_X1 U53 ( .A(n29), .ZN(n30) );
  AOI21_X1 U54 ( .B1(z[5]), .B2(n43), .A(n30), .ZN(n31) );
  NAND3_X1 U55 ( .A1(n9), .A2(n37), .A3(n31), .ZN(n51) );
  INV_X1 U56 ( .A(n32), .ZN(n33) );
  AOI221_X1 U57 ( .B1(n10), .B2(n47), .C1(z[6]), .C2(n43), .A(n33), .ZN(n36)
         );
  NAND4_X1 U58 ( .A1(n37), .A2(n62), .A3(n9), .A4(n36), .ZN(n69) );
  OAI21_X1 U59 ( .B1(n41), .B2(n2), .A(n38), .ZN(n53) );
  OAI21_X1 U60 ( .B1(n41), .B2(n3), .A(n38), .ZN(n54) );
  OAI21_X1 U61 ( .B1(n41), .B2(n4), .A(n38), .ZN(n55) );
  OAI21_X1 U62 ( .B1(n41), .B2(n5), .A(n38), .ZN(n56) );
  OAI21_X1 U63 ( .B1(n41), .B2(n6), .A(n38), .ZN(n61) );
  INV_X1 U64 ( .A(n42), .ZN(n45) );
endmodule


module layer3_16_12_16_16_B_rom_9 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b0;
  assign z[14] = 1'b0;
  assign z[13] = 1'b0;
  assign z[12] = 1'b0;
  assign z[11] = 1'b0;
  assign z[10] = 1'b0;
  assign z[9] = 1'b0;
  assign z[8] = 1'b0;
  assign z[7] = 1'b0;
  assign z[6] = 1'b0;
  assign z[5] = 1'b1;
  assign z[4] = 1'b1;
  assign z[3] = 1'b1;
  assign z[2] = 1'b1;
  assign z[1] = 1'b1;
  assign z[0] = 1'b1;

endmodule


module layer3_16_12_16_16_W_rom_10 ( clk, addr, z );
  input [3:0] addr;
  output [15:0] z;
  input clk;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n21, n38, n39, n41,
         n46, n47, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n13, n14, n15, n16, n17, n18, n19, n20, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n40, n42, n43, n44, n45, n48, n49, n50, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80;

  DFF_X1 \z_reg[15]  ( .D(n66), .CK(clk), .Q(z[15]), .QN(n1) );
  DFF_X1 \z_reg[13]  ( .D(n64), .CK(clk), .Q(z[13]), .QN(n3) );
  DFF_X1 \z_reg[12]  ( .D(n63), .CK(clk), .Q(z[12]), .QN(n4) );
  DFF_X1 \z_reg[11]  ( .D(n62), .CK(clk), .Q(z[11]), .QN(n5) );
  DFF_X1 \z_reg[10]  ( .D(n61), .CK(clk), .Q(z[10]), .QN(n6) );
  DFF_X1 \z_reg[9]  ( .D(n60), .CK(clk), .Q(z[9]), .QN(n7) );
  DFF_X1 \z_reg[8]  ( .D(n59), .CK(clk), .Q(z[8]), .QN(n8) );
  DFF_X1 \z_reg[7]  ( .D(n58), .CK(clk), .Q(z[7]), .QN(n9) );
  DFF_X1 \z_reg[6]  ( .D(n57), .CK(clk), .Q(z[6]), .QN(n10) );
  DFF_X1 \z_reg[5]  ( .D(n56), .CK(clk), .Q(z[5]) );
  DFF_X1 \z_reg[4]  ( .D(n55), .CK(clk), .Q(z[4]), .QN(n11) );
  DFF_X1 \z_reg[3]  ( .D(n54), .CK(clk), .Q(z[3]), .QN(n15) );
  DFF_X1 \z_reg[2]  ( .D(n53), .CK(clk), .Q(z[2]), .QN(n13) );
  DFF_X1 \z_reg[1]  ( .D(n52), .CK(clk), .Q(z[1]), .QN(n14) );
  DFF_X1 \z_reg[0]  ( .D(n51), .CK(clk), .Q(z[0]), .QN(n12) );
  DFF_X1 \z_reg[14]  ( .D(n65), .CK(clk), .Q(z[14]), .QN(n2) );
  AND2_X1 U3 ( .A1(n42), .A2(n50), .ZN(n16) );
  NAND3_X1 U4 ( .A1(n42), .A2(n35), .A3(n26), .ZN(n21) );
  INV_X1 U5 ( .A(n76), .ZN(n77) );
  NAND2_X1 U6 ( .A1(n47), .A2(n39), .ZN(n41) );
  NOR2_X1 U7 ( .A1(addr[3]), .A2(addr[2]), .ZN(n46) );
  NOR2_X1 U8 ( .A1(n78), .A2(addr[0]), .ZN(n47) );
  NOR2_X1 U9 ( .A1(n79), .A2(addr[1]), .ZN(n38) );
  OAI21_X1 U10 ( .B1(n21), .B2(n4), .A(n77), .ZN(n63) );
  OAI21_X1 U11 ( .B1(n21), .B2(n3), .A(n77), .ZN(n64) );
  OAI21_X1 U12 ( .B1(n21), .B2(n2), .A(n77), .ZN(n65) );
  OAI21_X1 U13 ( .B1(n21), .B2(n1), .A(n77), .ZN(n66) );
  AND2_X1 U14 ( .A1(addr[3]), .A2(n80), .ZN(n39) );
  NAND2_X1 U15 ( .A1(n47), .A2(n46), .ZN(n42) );
  NAND2_X1 U16 ( .A1(addr[1]), .A2(addr[0]), .ZN(n45) );
  INV_X1 U17 ( .A(n45), .ZN(n18) );
  INV_X1 U18 ( .A(addr[3]), .ZN(n17) );
  NAND2_X1 U19 ( .A1(addr[2]), .A2(n17), .ZN(n44) );
  INV_X1 U20 ( .A(n44), .ZN(n20) );
  NAND2_X1 U21 ( .A1(n18), .A2(n20), .ZN(n35) );
  NAND3_X1 U22 ( .A1(n39), .A2(addr[1]), .A3(addr[0]), .ZN(n75) );
  INV_X1 U23 ( .A(addr[0]), .ZN(n79) );
  INV_X1 U24 ( .A(addr[1]), .ZN(n78) );
  NAND3_X1 U25 ( .A1(n79), .A2(n78), .A3(n20), .ZN(n19) );
  NAND2_X1 U26 ( .A1(n75), .A2(n19), .ZN(n27) );
  NAND2_X1 U27 ( .A1(n38), .A2(n20), .ZN(n40) );
  NAND3_X1 U28 ( .A1(n46), .A2(addr[1]), .A3(addr[0]), .ZN(n71) );
  NAND2_X1 U29 ( .A1(n38), .A2(n46), .ZN(n50) );
  INV_X1 U30 ( .A(n50), .ZN(n24) );
  NAND2_X1 U31 ( .A1(n47), .A2(n20), .ZN(n34) );
  INV_X1 U32 ( .A(n34), .ZN(n23) );
  INV_X1 U33 ( .A(n39), .ZN(n22) );
  NAND3_X1 U34 ( .A1(n46), .A2(n79), .A3(n78), .ZN(n33) );
  OAI21_X1 U35 ( .B1(addr[1]), .B2(n22), .A(n33), .ZN(n28) );
  NOR3_X1 U36 ( .A1(n24), .A2(n23), .A3(n28), .ZN(n25) );
  NAND3_X1 U37 ( .A1(n40), .A2(n71), .A3(n25), .ZN(n76) );
  INV_X1 U38 ( .A(n41), .ZN(n31) );
  NOR3_X1 U39 ( .A1(n27), .A2(n76), .A3(n31), .ZN(n26) );
  INV_X1 U40 ( .A(n27), .ZN(n30) );
  INV_X1 U41 ( .A(n28), .ZN(n29) );
  NAND2_X1 U42 ( .A1(n30), .A2(n29), .ZN(n48) );
  NOR2_X1 U43 ( .A1(n31), .A2(n48), .ZN(n32) );
  OAI211_X1 U44 ( .C1(n12), .C2(n21), .A(n40), .B(n32), .ZN(n51) );
  INV_X1 U45 ( .A(n33), .ZN(n36) );
  NAND2_X1 U46 ( .A1(n41), .A2(n34), .ZN(n72) );
  NAND3_X1 U47 ( .A1(n35), .A2(n71), .A3(n75), .ZN(n67) );
  NOR3_X1 U48 ( .A1(n36), .A2(n72), .A3(n67), .ZN(n37) );
  OAI211_X1 U49 ( .C1(n21), .C2(n14), .A(n40), .B(n37), .ZN(n52) );
  INV_X1 U50 ( .A(n48), .ZN(n43) );
  OAI211_X1 U51 ( .C1(n21), .C2(n13), .A(n43), .B(n16), .ZN(n53) );
  INV_X1 U52 ( .A(addr[2]), .ZN(n80) );
  OAI221_X1 U53 ( .B1(addr[3]), .B2(n45), .C1(n80), .C2(n15), .A(n44), .ZN(n54) );
  NOR2_X1 U54 ( .A1(n72), .A2(n48), .ZN(n49) );
  OAI211_X1 U55 ( .C1(n11), .C2(n21), .A(n50), .B(n49), .ZN(n55) );
  INV_X1 U56 ( .A(n67), .ZN(n70) );
  INV_X1 U57 ( .A(n21), .ZN(n68) );
  AOI22_X1 U58 ( .A1(z[5]), .A2(n68), .B1(n38), .B2(n39), .ZN(n69) );
  NAND3_X1 U59 ( .A1(n70), .A2(n16), .A3(n69), .ZN(n56) );
  INV_X1 U60 ( .A(n71), .ZN(n73) );
  NOR2_X1 U61 ( .A1(n73), .A2(n72), .ZN(n74) );
  OAI211_X1 U62 ( .C1(n10), .C2(n21), .A(n75), .B(n74), .ZN(n57) );
  OAI21_X1 U63 ( .B1(n9), .B2(n21), .A(n77), .ZN(n58) );
  OAI21_X1 U64 ( .B1(n8), .B2(n21), .A(n77), .ZN(n59) );
  OAI21_X1 U65 ( .B1(n7), .B2(n21), .A(n77), .ZN(n60) );
  OAI21_X1 U66 ( .B1(n6), .B2(n21), .A(n77), .ZN(n61) );
  OAI21_X1 U67 ( .B1(n5), .B2(n21), .A(n77), .ZN(n62) );
endmodule


module layer3_16_12_16_16_B_rom_10 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b0;
  assign z[14] = 1'b0;
  assign z[13] = 1'b0;
  assign z[12] = 1'b0;
  assign z[11] = 1'b0;
  assign z[10] = 1'b0;
  assign z[9] = 1'b0;
  assign z[8] = 1'b0;
  assign z[7] = 1'b0;
  assign z[6] = 1'b1;
  assign z[5] = 1'b1;
  assign z[4] = 1'b1;
  assign z[3] = 1'b0;
  assign z[2] = 1'b1;
  assign z[1] = 1'b0;
  assign z[0] = 1'b0;

endmodule


module layer3_16_12_16_16_W_rom_11 ( clk, addr, z );
  input [3:0] addr;
  output [15:0] z;
  input clk;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n18, n33, n37, n39,
         n40, n41, n43, n44, n45, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n13, n14, n15, n16, n17, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n34,
         n35, n36, n38, n42, n46, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77;

  DFF_X1 \z_reg[15]  ( .D(n63), .CK(clk), .Q(z[15]), .QN(n1) );
  DFF_X1 \z_reg[14]  ( .D(n62), .CK(clk), .Q(z[14]), .QN(n2) );
  DFF_X1 \z_reg[13]  ( .D(n61), .CK(clk), .Q(z[13]), .QN(n3) );
  DFF_X1 \z_reg[12]  ( .D(n60), .CK(clk), .Q(z[12]), .QN(n4) );
  DFF_X1 \z_reg[11]  ( .D(n59), .CK(clk), .Q(z[11]), .QN(n5) );
  DFF_X1 \z_reg[10]  ( .D(n58), .CK(clk), .Q(z[10]), .QN(n6) );
  DFF_X1 \z_reg[9]  ( .D(n57), .CK(clk), .Q(z[9]), .QN(n7) );
  DFF_X1 \z_reg[8]  ( .D(n56), .CK(clk), .Q(z[8]), .QN(n8) );
  DFF_X1 \z_reg[7]  ( .D(n55), .CK(clk), .Q(z[7]), .QN(n9) );
  DFF_X1 \z_reg[6]  ( .D(n54), .CK(clk), .Q(z[6]) );
  DFF_X1 \z_reg[5]  ( .D(n53), .CK(clk), .Q(z[5]), .QN(n10) );
  DFF_X1 \z_reg[4]  ( .D(n52), .CK(clk), .Q(z[4]), .QN(n15) );
  DFF_X1 \z_reg[3]  ( .D(n51), .CK(clk), .Q(z[3]) );
  DFF_X1 \z_reg[2]  ( .D(n50), .CK(clk), .Q(z[2]), .QN(n11) );
  DFF_X1 \z_reg[1]  ( .D(n49), .CK(clk), .Q(z[1]), .QN(n13) );
  DFF_X1 \z_reg[0]  ( .D(n48), .CK(clk), .Q(z[0]), .QN(n12) );
  NAND3_X1 U47 ( .A1(addr[0]), .A2(n44), .A3(addr[2]), .ZN(n37) );
  NAND3_X1 U49 ( .A1(n76), .A2(n77), .A3(n45), .ZN(n33) );
  NAND3_X1 U50 ( .A1(n44), .A2(n76), .A3(addr[2]), .ZN(n39) );
  NAND3_X1 U52 ( .A1(addr[0]), .A2(n77), .A3(n45), .ZN(n41) );
  AND2_X1 U3 ( .A1(addr[1]), .A2(n45), .ZN(n14) );
  AND2_X1 U4 ( .A1(n39), .A2(n40), .ZN(n16) );
  NAND3_X1 U5 ( .A1(n24), .A2(n31), .A3(n20), .ZN(n18) );
  AND3_X1 U6 ( .A1(n41), .A2(n16), .A3(n74), .ZN(n17) );
  NAND2_X1 U7 ( .A1(n47), .A2(n76), .ZN(n40) );
  NOR3_X1 U8 ( .A1(addr[2]), .A2(addr[3]), .A3(addr[1]), .ZN(n47) );
  NOR3_X1 U9 ( .A1(addr[1]), .A2(addr[3]), .A3(n75), .ZN(n43) );
  NOR2_X1 U10 ( .A1(n77), .A2(addr[3]), .ZN(n44) );
  OAI21_X1 U11 ( .B1(n18), .B2(n4), .A(n17), .ZN(n60) );
  OAI21_X1 U12 ( .B1(n18), .B2(n3), .A(n17), .ZN(n61) );
  OAI21_X1 U13 ( .B1(n18), .B2(n2), .A(n17), .ZN(n62) );
  OAI21_X1 U14 ( .B1(n18), .B2(n1), .A(n17), .ZN(n63) );
  INV_X1 U15 ( .A(addr[1]), .ZN(n77) );
  AND2_X1 U16 ( .A1(addr[3]), .A2(n75), .ZN(n45) );
  INV_X1 U17 ( .A(addr[2]), .ZN(n75) );
  NAND3_X1 U18 ( .A1(n44), .A2(addr[0]), .A3(n75), .ZN(n21) );
  NAND2_X1 U19 ( .A1(n43), .A2(addr[0]), .ZN(n28) );
  NAND3_X1 U20 ( .A1(n41), .A2(n21), .A3(n28), .ZN(n32) );
  INV_X1 U21 ( .A(n32), .ZN(n24) );
  NAND2_X1 U22 ( .A1(n14), .A2(addr[0]), .ZN(n70) );
  NAND2_X1 U23 ( .A1(n33), .A2(n70), .ZN(n35) );
  INV_X1 U24 ( .A(n35), .ZN(n31) );
  INV_X1 U25 ( .A(addr[0]), .ZN(n76) );
  NAND3_X1 U26 ( .A1(n44), .A2(n75), .A3(n76), .ZN(n30) );
  NAND2_X1 U27 ( .A1(n16), .A2(n30), .ZN(n22) );
  INV_X1 U28 ( .A(n22), .ZN(n19) );
  NAND2_X1 U29 ( .A1(n14), .A2(n76), .ZN(n69) );
  NAND2_X1 U30 ( .A1(n43), .A2(n76), .ZN(n64) );
  NAND3_X1 U31 ( .A1(n19), .A2(n69), .A3(n64), .ZN(n25) );
  INV_X1 U32 ( .A(n37), .ZN(n38) );
  NOR3_X1 U33 ( .A1(n25), .A2(n38), .A3(n47), .ZN(n20) );
  INV_X1 U34 ( .A(n21), .ZN(n73) );
  NOR2_X1 U35 ( .A1(n73), .A2(n22), .ZN(n23) );
  OAI211_X1 U36 ( .C1(n12), .C2(n18), .A(n28), .B(n23), .ZN(n48) );
  OAI211_X1 U37 ( .C1(n18), .C2(n13), .A(n24), .B(n69), .ZN(n49) );
  INV_X1 U38 ( .A(n25), .ZN(n68) );
  INV_X1 U39 ( .A(n41), .ZN(n42) );
  INV_X1 U40 ( .A(n33), .ZN(n26) );
  NOR3_X1 U41 ( .A1(n47), .A2(n42), .A3(n26), .ZN(n27) );
  OAI211_X1 U42 ( .C1(n11), .C2(n18), .A(n68), .B(n27), .ZN(n50) );
  INV_X1 U43 ( .A(n18), .ZN(n66) );
  INV_X1 U44 ( .A(n28), .ZN(n65) );
  AOI21_X1 U45 ( .B1(z[3]), .B2(n66), .A(n65), .ZN(n29) );
  NAND3_X1 U46 ( .A1(n31), .A2(n30), .A3(n29), .ZN(n51) );
  INV_X1 U48 ( .A(n40), .ZN(n34) );
  NOR3_X1 U51 ( .A1(n35), .A2(n34), .A3(n32), .ZN(n36) );
  OAI211_X1 U53 ( .C1(n18), .C2(n15), .A(n64), .B(n36), .ZN(n52) );
  NOR3_X1 U54 ( .A1(n73), .A2(n42), .A3(n38), .ZN(n46) );
  OAI211_X1 U55 ( .C1(n10), .C2(n18), .A(n64), .B(n46), .ZN(n53) );
  AOI21_X1 U56 ( .B1(z[6]), .B2(n66), .A(n65), .ZN(n67) );
  NAND3_X1 U57 ( .A1(n68), .A2(n37), .A3(n67), .ZN(n54) );
  INV_X1 U58 ( .A(n69), .ZN(n72) );
  INV_X1 U59 ( .A(n70), .ZN(n71) );
  NOR3_X1 U60 ( .A1(n73), .A2(n72), .A3(n71), .ZN(n74) );
  OAI21_X1 U61 ( .B1(n9), .B2(n18), .A(n17), .ZN(n55) );
  OAI21_X1 U62 ( .B1(n8), .B2(n18), .A(n17), .ZN(n56) );
  OAI21_X1 U63 ( .B1(n7), .B2(n18), .A(n17), .ZN(n57) );
  OAI21_X1 U64 ( .B1(n6), .B2(n18), .A(n17), .ZN(n58) );
  OAI21_X1 U65 ( .B1(n5), .B2(n18), .A(n17), .ZN(n59) );
endmodule


module layer3_16_12_16_16_B_rom_11 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b0;
  assign z[14] = 1'b0;
  assign z[13] = 1'b0;
  assign z[12] = 1'b0;
  assign z[11] = 1'b0;
  assign z[10] = 1'b0;
  assign z[9] = 1'b0;
  assign z[8] = 1'b0;
  assign z[7] = 1'b0;
  assign z[6] = 1'b0;
  assign z[5] = 1'b1;
  assign z[4] = 1'b1;
  assign z[3] = 1'b0;
  assign z[2] = 1'b1;
  assign z[1] = 1'b0;
  assign z[0] = 1'b1;

endmodule


module layer3_16_12_16_16_W_rom_12 ( clk, addr, z );
  input [3:0] addr;
  output [15:0] z;
  input clk;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n20, n27,
         n29, n36, n37, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n15, n16, n17, n18, n19, n21, n22, n23, n24, n25, n26, n28, n30,
         n31, n32, n33, n34, n35, n38, n39, n66, n67, n68, n69, n70;

  DFF_X1 \z_reg[15]  ( .D(n65), .CK(clk), .Q(z[15]), .QN(n1) );
  DFF_X1 \z_reg[14]  ( .D(n64), .CK(clk), .Q(z[14]), .QN(n2) );
  DFF_X1 \z_reg[13]  ( .D(n63), .CK(clk), .Q(z[13]), .QN(n3) );
  DFF_X1 \z_reg[12]  ( .D(n62), .CK(clk), .Q(z[12]), .QN(n4) );
  DFF_X1 \z_reg[11]  ( .D(n61), .CK(clk), .Q(z[11]), .QN(n5) );
  DFF_X1 \z_reg[10]  ( .D(n60), .CK(clk), .Q(z[10]), .QN(n6) );
  DFF_X1 \z_reg[9]  ( .D(n59), .CK(clk), .Q(z[9]), .QN(n7) );
  DFF_X1 \z_reg[8]  ( .D(n58), .CK(clk), .Q(z[8]), .QN(n8) );
  DFF_X1 \z_reg[7]  ( .D(n57), .CK(clk), .Q(z[7]), .QN(n9) );
  DFF_X1 \z_reg[6]  ( .D(n56), .CK(clk), .Q(z[6]), .QN(n10) );
  DFF_X1 \z_reg[5]  ( .D(n55), .CK(clk), .Q(z[5]), .QN(n11) );
  DFF_X1 \z_reg[4]  ( .D(n54), .CK(clk), .Q(z[4]), .QN(n21) );
  DFF_X1 \z_reg[3]  ( .D(n53), .CK(clk), .Q(z[3]), .QN(n12) );
  DFF_X1 \z_reg[2]  ( .D(n52), .CK(clk), .Q(z[2]), .QN(n17) );
  DFF_X1 \z_reg[1]  ( .D(n51), .CK(clk), .Q(z[1]), .QN(n13) );
  DFF_X1 \z_reg[0]  ( .D(n50), .CK(clk), .Q(z[0]), .QN(n14) );
  NAND3_X1 U47 ( .A1(n68), .A2(n67), .A3(n45), .ZN(n36) );
  NAND3_X1 U48 ( .A1(addr[1]), .A2(n68), .A3(addr[0]), .ZN(n48) );
  NAND3_X1 U49 ( .A1(n70), .A2(n69), .A3(n49), .ZN(n37) );
  NAND3_X1 U50 ( .A1(n68), .A2(n67), .A3(n46), .ZN(n43) );
  NAND3_X1 U51 ( .A1(n47), .A2(addr[1]), .A3(addr[0]), .ZN(n40) );
  NAND3_X1 U52 ( .A1(addr[0]), .A2(addr[1]), .A3(n49), .ZN(n27) );
  NAND3_X1 U53 ( .A1(n70), .A2(n69), .A3(n47), .ZN(n41) );
  AND3_X1 U3 ( .A1(n29), .A2(n22), .A3(n66), .ZN(n15) );
  AND3_X1 U4 ( .A1(n48), .A2(n37), .A3(n19), .ZN(n16) );
  AND3_X1 U5 ( .A1(n40), .A2(n66), .A3(n39), .ZN(n18) );
  AND3_X1 U6 ( .A1(n27), .A2(n41), .A3(n33), .ZN(n19) );
  AND3_X1 U7 ( .A1(n43), .A2(n42), .A3(n40), .ZN(n22) );
  AND4_X1 U8 ( .A1(n37), .A2(n44), .A3(n41), .A4(n22), .ZN(n23) );
  NAND4_X1 U9 ( .A1(n36), .A2(n44), .A3(n15), .A4(n16), .ZN(n20) );
  NAND2_X1 U10 ( .A1(n46), .A2(n47), .ZN(n44) );
  NAND2_X1 U11 ( .A1(n49), .A2(n46), .ZN(n42) );
  NAND2_X1 U12 ( .A1(n45), .A2(n47), .ZN(n29) );
  NOR2_X1 U13 ( .A1(n68), .A2(addr[3]), .ZN(n47) );
  NOR2_X1 U14 ( .A1(n67), .A2(addr[2]), .ZN(n49) );
  NOR2_X1 U15 ( .A1(n70), .A2(addr[1]), .ZN(n46) );
  NOR2_X1 U16 ( .A1(n69), .A2(addr[0]), .ZN(n45) );
  OAI21_X1 U17 ( .B1(n20), .B2(n4), .A(n23), .ZN(n62) );
  OAI21_X1 U18 ( .B1(n20), .B2(n3), .A(n23), .ZN(n63) );
  OAI21_X1 U19 ( .B1(n20), .B2(n2), .A(n23), .ZN(n64) );
  OAI21_X1 U20 ( .B1(n20), .B2(n1), .A(n23), .ZN(n65) );
  INV_X1 U21 ( .A(addr[0]), .ZN(n70) );
  INV_X1 U22 ( .A(addr[2]), .ZN(n68) );
  INV_X1 U23 ( .A(addr[1]), .ZN(n69) );
  INV_X1 U24 ( .A(addr[3]), .ZN(n67) );
  NAND4_X1 U25 ( .A1(n70), .A2(n68), .A3(n69), .A4(n67), .ZN(n66) );
  NAND2_X1 U26 ( .A1(n49), .A2(n45), .ZN(n33) );
  OAI21_X1 U27 ( .B1(n14), .B2(n20), .A(n15), .ZN(n50) );
  NAND3_X1 U28 ( .A1(n27), .A2(n29), .A3(n66), .ZN(n31) );
  INV_X1 U29 ( .A(n31), .ZN(n26) );
  INV_X1 U30 ( .A(n42), .ZN(n35) );
  INV_X1 U31 ( .A(n41), .ZN(n24) );
  NOR2_X1 U32 ( .A1(n35), .A2(n24), .ZN(n25) );
  OAI211_X1 U33 ( .C1(n13), .C2(n20), .A(n26), .B(n25), .ZN(n51) );
  INV_X1 U34 ( .A(n44), .ZN(n30) );
  INV_X1 U35 ( .A(n43), .ZN(n28) );
  NOR3_X1 U36 ( .A1(n31), .A2(n30), .A3(n28), .ZN(n32) );
  OAI211_X1 U37 ( .C1(n20), .C2(n17), .A(n33), .B(n32), .ZN(n52) );
  INV_X1 U38 ( .A(n37), .ZN(n38) );
  INV_X1 U39 ( .A(n36), .ZN(n34) );
  NOR3_X1 U40 ( .A1(n38), .A2(n35), .A3(n34), .ZN(n39) );
  OAI21_X1 U41 ( .B1(n12), .B2(n20), .A(n18), .ZN(n53) );
  OAI211_X1 U42 ( .C1(n20), .C2(n21), .A(n16), .B(n66), .ZN(n54) );
  OAI211_X1 U43 ( .C1(n11), .C2(n20), .A(n18), .B(n43), .ZN(n55) );
  OAI211_X1 U44 ( .C1(n10), .C2(n20), .A(n15), .B(n19), .ZN(n56) );
  OAI21_X1 U45 ( .B1(n9), .B2(n20), .A(n23), .ZN(n57) );
  OAI21_X1 U46 ( .B1(n8), .B2(n20), .A(n23), .ZN(n58) );
  OAI21_X1 U54 ( .B1(n7), .B2(n20), .A(n23), .ZN(n59) );
  OAI21_X1 U55 ( .B1(n6), .B2(n20), .A(n23), .ZN(n60) );
  OAI21_X1 U56 ( .B1(n5), .B2(n20), .A(n23), .ZN(n61) );
endmodule


module layer3_16_12_16_16_B_rom_12 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b0;
  assign z[14] = 1'b0;
  assign z[13] = 1'b0;
  assign z[12] = 1'b0;
  assign z[11] = 1'b0;
  assign z[10] = 1'b0;
  assign z[9] = 1'b0;
  assign z[8] = 1'b0;
  assign z[7] = 1'b0;
  assign z[6] = 1'b0;
  assign z[5] = 1'b1;
  assign z[4] = 1'b1;
  assign z[3] = 1'b0;
  assign z[2] = 1'b0;
  assign z[1] = 1'b0;
  assign z[0] = 1'b1;

endmodule


module layer3_16_12_16_16_W_rom_13 ( clk, addr, z );
  input [3:0] addr;
  output [15:0] z;
  input clk;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n23, n40, n41,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n42, n63, n64, n65, n66, n67, n68, n69, n70, n71;

  DFF_X1 \z_reg[15]  ( .D(n62), .CK(clk), .Q(z[15]), .QN(n1) );
  DFF_X1 \z_reg[14]  ( .D(n61), .CK(clk), .Q(z[14]), .QN(n2) );
  DFF_X1 \z_reg[13]  ( .D(n60), .CK(clk), .Q(z[13]), .QN(n3) );
  DFF_X1 \z_reg[12]  ( .D(n59), .CK(clk), .Q(z[12]), .QN(n4) );
  DFF_X1 \z_reg[11]  ( .D(n58), .CK(clk), .Q(z[11]), .QN(n5) );
  DFF_X1 \z_reg[10]  ( .D(n57), .CK(clk), .Q(z[10]), .QN(n6) );
  DFF_X1 \z_reg[9]  ( .D(n56), .CK(clk), .Q(z[9]), .QN(n7) );
  DFF_X1 \z_reg[8]  ( .D(n55), .CK(clk), .Q(z[8]), .QN(n8) );
  DFF_X1 \z_reg[7]  ( .D(n54), .CK(clk), .Q(z[7]), .QN(n9) );
  DFF_X1 \z_reg[6]  ( .D(n53), .CK(clk), .Q(z[6]), .QN(n20) );
  DFF_X1 \z_reg[5]  ( .D(n52), .CK(clk), .Q(z[5]) );
  DFF_X1 \z_reg[4]  ( .D(n51), .CK(clk), .Q(z[4]), .QN(n18) );
  DFF_X1 \z_reg[3]  ( .D(n50), .CK(clk), .Q(z[3]), .QN(n10) );
  DFF_X1 \z_reg[2]  ( .D(n49), .CK(clk), .Q(z[2]), .QN(n11) );
  DFF_X1 \z_reg[1]  ( .D(n48), .CK(clk), .Q(z[1]), .QN(n12) );
  DFF_X1 \z_reg[0]  ( .D(n47), .CK(clk), .Q(z[0]), .QN(n13) );
  NAND3_X1 U45 ( .A1(n46), .A2(n69), .A3(addr[1]), .ZN(n41) );
  NAND3_X1 U47 ( .A1(n69), .A2(n71), .A3(addr[2]), .ZN(n43) );
  NAND3_X1 U51 ( .A1(n67), .A2(n71), .A3(n69), .ZN(n44) );
  AND2_X1 U3 ( .A1(n26), .A2(n30), .ZN(n14) );
  AND4_X1 U4 ( .A1(n41), .A2(n31), .A3(n36), .A4(n32), .ZN(n15) );
  AND2_X1 U5 ( .A1(n45), .A2(addr[2]), .ZN(n16) );
  AND2_X1 U6 ( .A1(n29), .A2(n43), .ZN(n17) );
  AND2_X1 U7 ( .A1(n41), .A2(n40), .ZN(n19) );
  NAND4_X1 U8 ( .A1(n44), .A2(n43), .A3(n21), .A4(n15), .ZN(n23) );
  AND4_X1 U9 ( .A1(n40), .A2(n14), .A3(n27), .A4(n33), .ZN(n21) );
  NAND2_X1 U10 ( .A1(n70), .A2(n68), .ZN(n40) );
  NOR2_X1 U11 ( .A1(n71), .A2(addr[2]), .ZN(n46) );
  NOR2_X1 U12 ( .A1(n69), .A2(addr[3]), .ZN(n45) );
  OAI21_X1 U13 ( .B1(n23), .B2(n4), .A(n21), .ZN(n59) );
  OAI21_X1 U14 ( .B1(n23), .B2(n3), .A(n21), .ZN(n60) );
  OAI21_X1 U15 ( .B1(n23), .B2(n2), .A(n21), .ZN(n61) );
  OAI21_X1 U16 ( .B1(n23), .B2(n1), .A(n21), .ZN(n62) );
  INV_X1 U17 ( .A(addr[3]), .ZN(n71) );
  INV_X1 U18 ( .A(addr[1]), .ZN(n68) );
  INV_X1 U19 ( .A(n44), .ZN(n22) );
  NAND2_X1 U20 ( .A1(n68), .A2(n22), .ZN(n26) );
  INV_X1 U21 ( .A(addr[2]), .ZN(n67) );
  NAND3_X1 U22 ( .A1(n45), .A2(n68), .A3(n67), .ZN(n30) );
  NAND2_X1 U23 ( .A1(n16), .A2(n68), .ZN(n27) );
  NAND3_X1 U24 ( .A1(n46), .A2(addr[0]), .A3(n68), .ZN(n33) );
  INV_X1 U25 ( .A(n45), .ZN(n24) );
  NAND3_X1 U26 ( .A1(n46), .A2(addr[1]), .A3(addr[0]), .ZN(n66) );
  OAI21_X1 U27 ( .B1(addr[2]), .B2(n24), .A(n66), .ZN(n25) );
  INV_X1 U28 ( .A(n25), .ZN(n31) );
  NAND2_X1 U29 ( .A1(n16), .A2(addr[1]), .ZN(n36) );
  INV_X1 U30 ( .A(addr[0]), .ZN(n69) );
  NAND3_X1 U31 ( .A1(n46), .A2(n68), .A3(n69), .ZN(n32) );
  NAND2_X1 U32 ( .A1(n27), .A2(n26), .ZN(n34) );
  INV_X1 U33 ( .A(n34), .ZN(n28) );
  NAND2_X1 U34 ( .A1(n19), .A2(n28), .ZN(n42) );
  INV_X1 U35 ( .A(n42), .ZN(n29) );
  OAI21_X1 U36 ( .B1(n13), .B2(n23), .A(n17), .ZN(n47) );
  OAI211_X1 U37 ( .C1(n12), .C2(n23), .A(n30), .B(n17), .ZN(n48) );
  OAI211_X1 U38 ( .C1(n11), .C2(n23), .A(n31), .B(n14), .ZN(n49) );
  OAI21_X1 U39 ( .B1(n10), .B2(n23), .A(n15), .ZN(n50) );
  INV_X1 U40 ( .A(n32), .ZN(n64) );
  INV_X1 U41 ( .A(n33), .ZN(n63) );
  NOR3_X1 U42 ( .A1(n64), .A2(n63), .A3(n34), .ZN(n35) );
  OAI211_X1 U43 ( .C1(n23), .C2(n18), .A(n36), .B(n35), .ZN(n51) );
  INV_X1 U44 ( .A(n23), .ZN(n38) );
  INV_X1 U46 ( .A(n36), .ZN(n37) );
  AOI21_X1 U48 ( .B1(z[5]), .B2(n38), .A(n37), .ZN(n39) );
  NAND3_X1 U49 ( .A1(n19), .A2(n14), .A3(n39), .ZN(n52) );
  NOR3_X1 U50 ( .A1(n64), .A2(n63), .A3(n42), .ZN(n65) );
  OAI211_X1 U52 ( .C1(n23), .C2(n20), .A(n66), .B(n65), .ZN(n53) );
  OAI21_X1 U53 ( .B1(n9), .B2(n23), .A(n21), .ZN(n54) );
  OAI21_X1 U54 ( .B1(n8), .B2(n23), .A(n21), .ZN(n55) );
  OAI21_X1 U55 ( .B1(n7), .B2(n23), .A(n21), .ZN(n56) );
  OAI21_X1 U56 ( .B1(n6), .B2(n23), .A(n21), .ZN(n57) );
  OAI21_X1 U57 ( .B1(n5), .B2(n23), .A(n21), .ZN(n58) );
  INV_X1 U58 ( .A(n43), .ZN(n70) );
endmodule


module layer3_16_12_16_16_B_rom_13 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b0;
  assign z[14] = 1'b0;
  assign z[13] = 1'b0;
  assign z[12] = 1'b0;
  assign z[11] = 1'b0;
  assign z[10] = 1'b0;
  assign z[9] = 1'b0;
  assign z[8] = 1'b0;
  assign z[7] = 1'b0;
  assign z[6] = 1'b1;
  assign z[5] = 1'b0;
  assign z[4] = 1'b1;
  assign z[3] = 1'b0;
  assign z[2] = 1'b1;
  assign z[1] = 1'b0;
  assign z[0] = 1'b1;

endmodule


module layer3_16_12_16_16_W_rom_14 ( clk, addr, z );
  input [3:0] addr;
  output [15:0] z;
  input clk;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n19, n35,
         n36, n37, n38, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n15, n16, n17, n18,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n39, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72;

  DFF_X1 \z_reg[15]  ( .D(n60), .CK(clk), .Q(z[15]), .QN(n1) );
  DFF_X1 \z_reg[14]  ( .D(n59), .CK(clk), .Q(z[14]), .QN(n2) );
  DFF_X1 \z_reg[13]  ( .D(n58), .CK(clk), .Q(z[13]), .QN(n3) );
  DFF_X1 \z_reg[12]  ( .D(n57), .CK(clk), .Q(z[12]), .QN(n4) );
  DFF_X1 \z_reg[11]  ( .D(n56), .CK(clk), .Q(z[11]), .QN(n5) );
  DFF_X1 \z_reg[10]  ( .D(n55), .CK(clk), .Q(z[10]), .QN(n6) );
  DFF_X1 \z_reg[9]  ( .D(n54), .CK(clk), .Q(z[9]), .QN(n7) );
  DFF_X1 \z_reg[8]  ( .D(n53), .CK(clk), .Q(z[8]), .QN(n8) );
  DFF_X1 \z_reg[7]  ( .D(n52), .CK(clk), .Q(z[7]), .QN(n9) );
  DFF_X1 \z_reg[6]  ( .D(n51), .CK(clk), .Q(z[6]) );
  DFF_X1 \z_reg[5]  ( .D(n50), .CK(clk), .Q(z[5]), .QN(n10) );
  DFF_X1 \z_reg[4]  ( .D(n49), .CK(clk), .Q(z[4]), .QN(n11) );
  DFF_X1 \z_reg[3]  ( .D(n48), .CK(clk), .Q(z[3]), .QN(n12) );
  DFF_X1 \z_reg[2]  ( .D(n47), .CK(clk), .Q(z[2]), .QN(n16) );
  DFF_X1 \z_reg[1]  ( .D(n46), .CK(clk), .Q(z[1]), .QN(n13) );
  DFF_X1 \z_reg[0]  ( .D(n45), .CK(clk), .Q(z[0]), .QN(n14) );
  NAND3_X1 U40 ( .A1(n41), .A2(n71), .A3(addr[2]), .ZN(n38) );
  NAND3_X1 U42 ( .A1(addr[2]), .A2(addr[1]), .A3(n42), .ZN(n37) );
  NAND3_X1 U45 ( .A1(n43), .A2(n72), .A3(addr[3]), .ZN(n36) );
  NAND3_X1 U46 ( .A1(n71), .A2(n70), .A3(n42), .ZN(n40) );
  NAND3_X1 U47 ( .A1(addr[2]), .A2(n71), .A3(n42), .ZN(n35) );
  NAND3_X1 U48 ( .A1(addr[0]), .A2(n70), .A3(addr[3]), .ZN(n44) );
  AND3_X1 U3 ( .A1(n36), .A2(n69), .A3(n18), .ZN(n15) );
  AND4_X1 U4 ( .A1(n36), .A2(n37), .A3(n40), .A4(n24), .ZN(n17) );
  AND2_X1 U5 ( .A1(n37), .A2(n38), .ZN(n18) );
  NAND4_X1 U6 ( .A1(n44), .A2(n17), .A3(n29), .A4(n69), .ZN(n19) );
  AND4_X1 U7 ( .A1(n40), .A2(n18), .A3(n69), .A4(n68), .ZN(n20) );
  NOR2_X1 U8 ( .A1(n72), .A2(addr[3]), .ZN(n42) );
  NOR2_X1 U9 ( .A1(n71), .A2(addr[2]), .ZN(n43) );
  OAI21_X1 U10 ( .B1(n19), .B2(n4), .A(n20), .ZN(n57) );
  OAI21_X1 U11 ( .B1(n19), .B2(n3), .A(n20), .ZN(n58) );
  OAI21_X1 U12 ( .B1(n19), .B2(n2), .A(n20), .ZN(n59) );
  OAI21_X1 U13 ( .B1(n19), .B2(n1), .A(n20), .ZN(n60) );
  NOR2_X1 U14 ( .A1(addr[3]), .A2(addr[0]), .ZN(n41) );
  NAND3_X1 U15 ( .A1(n43), .A2(addr[3]), .A3(addr[0]), .ZN(n33) );
  INV_X1 U16 ( .A(n33), .ZN(n23) );
  INV_X1 U17 ( .A(n41), .ZN(n22) );
  INV_X1 U18 ( .A(n43), .ZN(n21) );
  INV_X1 U19 ( .A(addr[1]), .ZN(n71) );
  INV_X1 U20 ( .A(addr[2]), .ZN(n70) );
  NAND3_X1 U21 ( .A1(n41), .A2(n71), .A3(n70), .ZN(n68) );
  OAI21_X1 U22 ( .B1(n22), .B2(n21), .A(n68), .ZN(n31) );
  OAI21_X1 U23 ( .B1(n70), .B2(n22), .A(n35), .ZN(n63) );
  NOR3_X1 U24 ( .A1(n23), .A2(n31), .A3(n63), .ZN(n24) );
  NAND2_X1 U25 ( .A1(n42), .A2(n43), .ZN(n29) );
  INV_X1 U26 ( .A(addr[0]), .ZN(n72) );
  NAND4_X1 U27 ( .A1(addr[3]), .A2(n71), .A3(n72), .A4(n70), .ZN(n69) );
  INV_X1 U28 ( .A(n69), .ZN(n26) );
  INV_X1 U29 ( .A(n38), .ZN(n25) );
  INV_X1 U30 ( .A(n40), .ZN(n39) );
  NOR3_X1 U31 ( .A1(n26), .A2(n25), .A3(n39), .ZN(n27) );
  OAI211_X1 U32 ( .C1(n14), .C2(n19), .A(n33), .B(n27), .ZN(n45) );
  OAI211_X1 U33 ( .C1(n13), .C2(n19), .A(n15), .B(n35), .ZN(n46) );
  INV_X1 U34 ( .A(n31), .ZN(n28) );
  OAI211_X1 U35 ( .C1(n19), .C2(n16), .A(n15), .B(n28), .ZN(n47) );
  INV_X1 U36 ( .A(n29), .ZN(n64) );
  INV_X1 U37 ( .A(n44), .ZN(n30) );
  NOR3_X1 U38 ( .A1(n64), .A2(n31), .A3(n30), .ZN(n32) );
  OAI211_X1 U39 ( .C1(n12), .C2(n19), .A(n33), .B(n32), .ZN(n48) );
  INV_X1 U41 ( .A(n35), .ZN(n61) );
  INV_X1 U43 ( .A(n36), .ZN(n34) );
  NOR3_X1 U44 ( .A1(n61), .A2(n39), .A3(n34), .ZN(n62) );
  OAI211_X1 U49 ( .C1(n11), .C2(n19), .A(n69), .B(n62), .ZN(n49) );
  OAI21_X1 U50 ( .B1(n10), .B2(n19), .A(n17), .ZN(n50) );
  INV_X1 U51 ( .A(n63), .ZN(n67) );
  INV_X1 U52 ( .A(n19), .ZN(n65) );
  AOI21_X1 U53 ( .B1(z[6]), .B2(n65), .A(n64), .ZN(n66) );
  NAND3_X1 U54 ( .A1(n15), .A2(n67), .A3(n66), .ZN(n51) );
  OAI21_X1 U55 ( .B1(n9), .B2(n19), .A(n20), .ZN(n52) );
  OAI21_X1 U56 ( .B1(n8), .B2(n19), .A(n20), .ZN(n53) );
  OAI21_X1 U57 ( .B1(n7), .B2(n19), .A(n20), .ZN(n54) );
  OAI21_X1 U58 ( .B1(n6), .B2(n19), .A(n20), .ZN(n55) );
  OAI21_X1 U59 ( .B1(n5), .B2(n19), .A(n20), .ZN(n56) );
endmodule


module layer3_16_12_16_16_B_rom_14 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b1;
  assign z[14] = 1'b1;
  assign z[13] = 1'b1;
  assign z[12] = 1'b1;
  assign z[11] = 1'b1;
  assign z[10] = 1'b1;
  assign z[9] = 1'b1;
  assign z[8] = 1'b1;
  assign z[7] = 1'b1;
  assign z[6] = 1'b0;
  assign z[5] = 1'b0;
  assign z[4] = 1'b1;
  assign z[3] = 1'b1;
  assign z[2] = 1'b1;
  assign z[1] = 1'b0;
  assign z[0] = 1'b0;

endmodule


module layer3_16_12_16_16_W_rom_15 ( clk, addr, z );
  input [3:0] addr;
  output [15:0] z;
  input clk;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n19, n30, n34,
         n35, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n12, n15, n16, n17,
         n18, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n31, n32, n33,
         n36, n37, n38, n39, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77;

  DFF_X1 \z_reg[15]  ( .D(n62), .CK(clk), .Q(z[15]), .QN(n1) );
  DFF_X1 \z_reg[14]  ( .D(n61), .CK(clk), .Q(z[14]), .QN(n2) );
  DFF_X1 \z_reg[13]  ( .D(n60), .CK(clk), .Q(z[13]), .QN(n3) );
  DFF_X1 \z_reg[12]  ( .D(n59), .CK(clk), .Q(z[12]), .QN(n4) );
  DFF_X1 \z_reg[11]  ( .D(n58), .CK(clk), .Q(z[11]), .QN(n5) );
  DFF_X1 \z_reg[10]  ( .D(n57), .CK(clk), .Q(z[10]), .QN(n6) );
  DFF_X1 \z_reg[9]  ( .D(n56), .CK(clk), .Q(z[9]), .QN(n7) );
  DFF_X1 \z_reg[8]  ( .D(n55), .CK(clk), .Q(z[8]), .QN(n8) );
  DFF_X1 \z_reg[7]  ( .D(n54), .CK(clk), .Q(z[7]), .QN(n9) );
  DFF_X1 \z_reg[6]  ( .D(n53), .CK(clk), .Q(z[6]), .QN(n10) );
  DFF_X1 \z_reg[5]  ( .D(n52), .CK(clk), .Q(z[5]) );
  DFF_X1 \z_reg[4]  ( .D(n51), .CK(clk), .Q(z[4]), .QN(n11) );
  DFF_X1 \z_reg[3]  ( .D(n50), .CK(clk), .Q(z[3]) );
  DFF_X1 \z_reg[2]  ( .D(n49), .CK(clk), .Q(z[2]), .QN(n13) );
  DFF_X1 \z_reg[1]  ( .D(n48), .CK(clk), .Q(z[1]), .QN(n12) );
  DFF_X1 \z_reg[0]  ( .D(n47), .CK(clk), .Q(z[0]), .QN(n14) );
  NAND3_X1 U45 ( .A1(n44), .A2(addr[2]), .A3(addr[0]), .ZN(n43) );
  NAND3_X1 U46 ( .A1(addr[2]), .A2(n77), .A3(n44), .ZN(n35) );
  NAND3_X1 U47 ( .A1(n42), .A2(n77), .A3(addr[2]), .ZN(n40) );
  NAND3_X1 U48 ( .A1(n45), .A2(n76), .A3(addr[3]), .ZN(n34) );
  AND3_X1 U3 ( .A1(n34), .A2(n40), .A3(n35), .ZN(n46) );
  AND2_X1 U4 ( .A1(addr[3]), .A2(n41), .ZN(n15) );
  AND2_X1 U5 ( .A1(n69), .A2(n25), .ZN(n16) );
  NAND3_X1 U6 ( .A1(n43), .A2(n24), .A3(n18), .ZN(n19) );
  AND3_X1 U7 ( .A1(n16), .A2(n75), .A3(n74), .ZN(n17) );
  AND4_X1 U8 ( .A1(n46), .A2(n70), .A3(n32), .A4(n16), .ZN(n18) );
  NAND2_X1 U9 ( .A1(n45), .A2(n42), .ZN(n30) );
  NOR2_X1 U10 ( .A1(addr[3]), .A2(addr[1]), .ZN(n42) );
  NOR2_X1 U11 ( .A1(n77), .A2(addr[2]), .ZN(n45) );
  NOR2_X1 U12 ( .A1(n76), .A2(addr[3]), .ZN(n44) );
  NOR2_X1 U13 ( .A1(addr[2]), .A2(addr[0]), .ZN(n41) );
  OAI21_X1 U14 ( .B1(n19), .B2(n4), .A(n17), .ZN(n59) );
  OAI21_X1 U15 ( .B1(n19), .B2(n3), .A(n17), .ZN(n60) );
  OAI21_X1 U16 ( .B1(n19), .B2(n2), .A(n17), .ZN(n61) );
  OAI21_X1 U17 ( .B1(n19), .B2(n1), .A(n17), .ZN(n62) );
  INV_X1 U18 ( .A(addr[0]), .ZN(n77) );
  INV_X1 U19 ( .A(n41), .ZN(n21) );
  INV_X1 U20 ( .A(n42), .ZN(n20) );
  NAND2_X1 U21 ( .A1(n15), .A2(addr[1]), .ZN(n75) );
  OAI211_X1 U22 ( .C1(n21), .C2(n20), .A(n30), .B(n75), .ZN(n29) );
  INV_X1 U23 ( .A(n29), .ZN(n24) );
  INV_X1 U24 ( .A(n44), .ZN(n23) );
  INV_X1 U25 ( .A(n45), .ZN(n22) );
  NAND3_X1 U26 ( .A1(addr[2]), .A2(n42), .A3(addr[0]), .ZN(n63) );
  OAI21_X1 U27 ( .B1(n23), .B2(n22), .A(n63), .ZN(n27) );
  INV_X1 U28 ( .A(n27), .ZN(n70) );
  INV_X1 U29 ( .A(addr[1]), .ZN(n76) );
  NAND2_X1 U30 ( .A1(n15), .A2(n76), .ZN(n32) );
  NAND3_X1 U31 ( .A1(n45), .A2(addr[3]), .A3(addr[1]), .ZN(n69) );
  NAND2_X1 U32 ( .A1(n44), .A2(n41), .ZN(n25) );
  OAI21_X1 U33 ( .B1(n14), .B2(n19), .A(n18), .ZN(n47) );
  NAND4_X1 U34 ( .A1(n35), .A2(n30), .A3(n34), .A4(n25), .ZN(n33) );
  INV_X1 U35 ( .A(n33), .ZN(n26) );
  OAI211_X1 U36 ( .C1(n19), .C2(n12), .A(n26), .B(n63), .ZN(n48) );
  NOR2_X1 U37 ( .A1(n29), .A2(n27), .ZN(n28) );
  OAI211_X1 U38 ( .C1(n13), .C2(n19), .A(n32), .B(n28), .ZN(n49) );
  INV_X1 U39 ( .A(n19), .ZN(n66) );
  INV_X1 U40 ( .A(n69), .ZN(n39) );
  AOI211_X1 U41 ( .C1(z[3]), .C2(n66), .A(n39), .B(n29), .ZN(n31) );
  NAND4_X1 U42 ( .A1(n35), .A2(n40), .A3(n34), .A4(n31), .ZN(n50) );
  INV_X1 U43 ( .A(n32), .ZN(n73) );
  NOR2_X1 U44 ( .A1(n73), .A2(n33), .ZN(n36) );
  OAI211_X1 U49 ( .C1(n11), .C2(n19), .A(n69), .B(n36), .ZN(n51) );
  INV_X1 U50 ( .A(n40), .ZN(n71) );
  INV_X1 U51 ( .A(n30), .ZN(n38) );
  INV_X1 U52 ( .A(n43), .ZN(n37) );
  NOR4_X1 U53 ( .A1(n39), .A2(n71), .A3(n38), .A4(n37), .ZN(n68) );
  INV_X1 U54 ( .A(n75), .ZN(n65) );
  INV_X1 U55 ( .A(n63), .ZN(n64) );
  AOI211_X1 U56 ( .C1(z[5]), .C2(n66), .A(n65), .B(n64), .ZN(n67) );
  NAND2_X1 U57 ( .A1(n68), .A2(n67), .ZN(n52) );
  OAI211_X1 U58 ( .C1(n10), .C2(n19), .A(n70), .B(n69), .ZN(n53) );
  INV_X1 U59 ( .A(n34), .ZN(n72) );
  NOR3_X1 U60 ( .A1(n73), .A2(n72), .A3(n71), .ZN(n74) );
  OAI21_X1 U61 ( .B1(n9), .B2(n19), .A(n17), .ZN(n54) );
  OAI21_X1 U62 ( .B1(n8), .B2(n19), .A(n17), .ZN(n55) );
  OAI21_X1 U63 ( .B1(n7), .B2(n19), .A(n17), .ZN(n56) );
  OAI21_X1 U64 ( .B1(n6), .B2(n19), .A(n17), .ZN(n57) );
  OAI21_X1 U65 ( .B1(n5), .B2(n19), .A(n17), .ZN(n58) );
endmodule


module layer3_16_12_16_16_B_rom_15 ( clk, addr, z );
  input [0:0] addr;
  output [15:0] z;
  input clk;

  assign z[15] = 1'b1;
  assign z[14] = 1'b1;
  assign z[13] = 1'b1;
  assign z[12] = 1'b1;
  assign z[11] = 1'b1;
  assign z[10] = 1'b1;
  assign z[9] = 1'b1;
  assign z[8] = 1'b1;
  assign z[7] = 1'b1;
  assign z[6] = 1'b0;
  assign z[5] = 1'b0;
  assign z[4] = 1'b0;
  assign z[3] = 1'b1;
  assign z[2] = 1'b0;
  assign z[1] = 1'b0;
  assign z[0] = 1'b0;

endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_0_DW_mult_tc_1 ( a, b, 
        product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n9, n12, n13, n16, n18, n19, n21, n23, n25, n29, n31, n32,
         n34, n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n50, n51,
         n53, n54, n55, n56, n57, n58, n59, n62, n63, n64, n65, n67, n69, n70,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n93, n95, n96, n97, n98, n103, n104,
         n105, n106, n107, n111, n112, n113, n114, n115, n117, n119, n120,
         n122, n125, n126, n127, n135, n139, n141, n142, n143, n145, n146,
         n147, n148, n149, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n247,
         n249, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n418, n419, n420, n421, n422,
         n423, n424, n426, n427, n431, n433, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U150 ( .A(n271), .B(n146), .Z(n147) );
  XOR2_X1 U152 ( .A(n301), .B(n148), .Z(n149) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U161 ( .A(n177), .B(n168), .CI(n166), .CO(n163), .S(n164) );
  FA_X1 U162 ( .A(n170), .B(n172), .CI(n179), .CO(n165), .S(n166) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n263), .CI(n291), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n317), .B(n252), .CO(n173), .S(n174) );
  FA_X1 U170 ( .A(n268), .B(n292), .CI(n274), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U173 ( .A(n199), .B(n201), .CI(n192), .CO(n187), .S(n188) );
  FA_X1 U174 ( .A(n275), .B(n293), .CI(n194), .CO(n189), .S(n190) );
  HA_X1 U176 ( .A(n269), .B(n319), .CO(n193), .S(n194) );
  FA_X1 U177 ( .A(n205), .B(n200), .CI(n198), .CO(n195), .S(n196) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U179 ( .A(n276), .B(n294), .CI(n284), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n306), .B(n270), .CI(n320), .CO(n201), .S(n202) );
  FA_X1 U181 ( .A(n208), .B(n213), .CI(n206), .CO(n203), .S(n204) );
  FA_X1 U182 ( .A(n210), .B(n307), .CI(n215), .CO(n205), .S(n206) );
  FA_X1 U183 ( .A(n295), .B(n285), .CI(n254), .CO(n207), .S(n208) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n322), .B(n278), .CI(n308), .CO(n215), .S(n216) );
  FA_X1 U188 ( .A(n225), .B(n222), .CI(n220), .CO(n217), .S(n218) );
  FA_X1 U189 ( .A(n297), .B(n309), .CI(n255), .CO(n219), .S(n220) );
  HA_X1 U190 ( .A(n287), .B(n323), .CO(n221), .S(n222) );
  FA_X1 U192 ( .A(n288), .B(n324), .CI(n310), .CO(n225), .S(n226) );
  HA_X1 U194 ( .A(n311), .B(n325), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n326), .B(n300), .CI(n312), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  BUF_X1 U414 ( .A(n528), .Z(n490) );
  OR2_X2 U415 ( .A1(n491), .A2(n564), .ZN(n34) );
  XOR2_X1 U416 ( .A(n613), .B(a[10]), .Z(n491) );
  OR2_X1 U417 ( .A1(n218), .A2(n223), .ZN(n492) );
  AND2_X1 U418 ( .A1(n232), .A2(n233), .ZN(n493) );
  INV_X2 U419 ( .A(n570), .ZN(n21) );
  XNOR2_X1 U420 ( .A(n226), .B(n494), .ZN(n224) );
  XNOR2_X1 U421 ( .A(n229), .B(n298), .ZN(n494) );
  BUF_X1 U422 ( .A(n45), .Z(n495) );
  OR2_X1 U423 ( .A1(n550), .A2(n570), .ZN(n540) );
  OR2_X1 U424 ( .A1(n550), .A2(n570), .ZN(n23) );
  CLKBUF_X3 U425 ( .A(n601), .Z(n506) );
  NAND2_X2 U426 ( .A1(n433), .A2(n548), .ZN(n583) );
  INV_X1 U427 ( .A(n613), .ZN(n612) );
  INV_X1 U428 ( .A(n522), .ZN(n37) );
  OR2_X1 U429 ( .A1(n329), .A2(n258), .ZN(n496) );
  INV_X1 U430 ( .A(n575), .ZN(n16) );
  INV_X1 U431 ( .A(n555), .ZN(n497) );
  CLKBUF_X1 U432 ( .A(n7), .Z(n534) );
  XNOR2_X1 U433 ( .A(n498), .B(n178), .ZN(n176) );
  XNOR2_X1 U434 ( .A(n501), .B(n187), .ZN(n498) );
  BUF_X1 U435 ( .A(n562), .Z(n571) );
  XNOR2_X1 U436 ( .A(n45), .B(n499), .ZN(product[12]) );
  AND2_X1 U437 ( .A1(n126), .A2(n79), .ZN(n499) );
  INV_X1 U438 ( .A(n611), .ZN(n500) );
  INV_X1 U439 ( .A(n611), .ZN(n610) );
  XOR2_X1 U440 ( .A(n602), .B(a[2]), .Z(n9) );
  XOR2_X1 U441 ( .A(n526), .B(n551), .Z(n501) );
  OAI22_X1 U442 ( .A1(n23), .A2(n359), .B1(n358), .B2(n21), .ZN(n502) );
  AOI21_X1 U443 ( .B1(n104), .B2(n590), .A(n580), .ZN(n503) );
  XNOR2_X1 U444 ( .A(n214), .B(n504), .ZN(n212) );
  XNOR2_X1 U445 ( .A(n216), .B(n219), .ZN(n504) );
  OAI21_X1 U446 ( .B1(n503), .B2(n97), .A(n98), .ZN(n505) );
  BUF_X2 U447 ( .A(n601), .Z(n507) );
  INV_X1 U448 ( .A(n602), .ZN(n601) );
  XOR2_X1 U449 ( .A(n305), .B(n283), .Z(n508) );
  XOR2_X1 U450 ( .A(n508), .B(n253), .Z(n192) );
  NAND2_X1 U451 ( .A1(n253), .A2(n502), .ZN(n509) );
  NAND2_X1 U452 ( .A1(n253), .A2(n305), .ZN(n510) );
  NAND2_X1 U453 ( .A1(n502), .A2(n305), .ZN(n511) );
  NAND3_X1 U454 ( .A1(n509), .A2(n510), .A3(n511), .ZN(n191) );
  BUF_X1 U455 ( .A(n191), .Z(n526) );
  OR2_X2 U456 ( .A1(n512), .A2(n555), .ZN(n29) );
  XNOR2_X1 U457 ( .A(n610), .B(a[8]), .ZN(n512) );
  INV_X1 U458 ( .A(n532), .ZN(n513) );
  BUF_X2 U459 ( .A(n602), .Z(n532) );
  CLKBUF_X1 U460 ( .A(n85), .Z(n514) );
  XOR2_X1 U461 ( .A(n182), .B(n184), .Z(n515) );
  XOR2_X1 U462 ( .A(n515), .B(n189), .Z(n178) );
  NAND2_X1 U463 ( .A1(n182), .A2(n184), .ZN(n516) );
  NAND2_X1 U464 ( .A1(n182), .A2(n189), .ZN(n517) );
  NAND2_X1 U465 ( .A1(n184), .A2(n189), .ZN(n518) );
  NAND3_X1 U466 ( .A1(n516), .A2(n517), .A3(n518), .ZN(n177) );
  NAND2_X1 U467 ( .A1(n501), .A2(n187), .ZN(n519) );
  NAND2_X1 U468 ( .A1(n501), .A2(n178), .ZN(n520) );
  NAND2_X1 U469 ( .A1(n187), .A2(n178), .ZN(n521) );
  NAND3_X1 U470 ( .A1(n519), .A2(n520), .A3(n521), .ZN(n175) );
  XNOR2_X1 U471 ( .A(n613), .B(a[12]), .ZN(n522) );
  OAI21_X1 U472 ( .B1(n86), .B2(n82), .A(n83), .ZN(n81) );
  XNOR2_X1 U473 ( .A(n536), .B(a[2]), .ZN(n585) );
  CLKBUF_X1 U474 ( .A(n78), .Z(n523) );
  FA_X1 U475 ( .A(n205), .B(n200), .CI(n198), .S(n524) );
  XNOR2_X1 U476 ( .A(n532), .B(n249), .ZN(n525) );
  CLKBUF_X1 U477 ( .A(n104), .Z(n527) );
  XNOR2_X1 U478 ( .A(n607), .B(a[4]), .ZN(n431) );
  INV_X1 U479 ( .A(n607), .ZN(n605) );
  INV_X1 U480 ( .A(n13), .ZN(n607) );
  NAND2_X1 U481 ( .A1(n524), .A2(n203), .ZN(n528) );
  BUF_X1 U482 ( .A(n230), .Z(n529) );
  OR2_X1 U483 ( .A1(n196), .A2(n203), .ZN(n530) );
  INV_X1 U484 ( .A(n575), .ZN(n531) );
  INV_X1 U485 ( .A(n247), .ZN(n533) );
  XOR2_X1 U486 ( .A(n609), .B(a[6]), .Z(n550) );
  CLKBUF_X1 U487 ( .A(n532), .Z(n535) );
  INV_X1 U488 ( .A(n556), .ZN(n73) );
  INV_X1 U489 ( .A(n7), .ZN(n536) );
  INV_X1 U490 ( .A(n7), .ZN(n537) );
  OR2_X1 U491 ( .A1(n204), .A2(n211), .ZN(n538) );
  CLKBUF_X1 U492 ( .A(n32), .Z(n539) );
  CLKBUF_X1 U493 ( .A(n503), .Z(n541) );
  XNOR2_X1 U494 ( .A(n532), .B(n249), .ZN(n433) );
  CLKBUF_X1 U495 ( .A(n115), .Z(n542) );
  BUF_X1 U496 ( .A(n563), .Z(n543) );
  XNOR2_X1 U497 ( .A(n188), .B(n544), .ZN(n186) );
  XNOR2_X1 U498 ( .A(n197), .B(n190), .ZN(n544) );
  NAND2_X1 U499 ( .A1(n188), .A2(n197), .ZN(n545) );
  NAND2_X1 U500 ( .A1(n188), .A2(n190), .ZN(n546) );
  NAND2_X1 U501 ( .A1(n197), .A2(n190), .ZN(n547) );
  NAND3_X1 U502 ( .A1(n545), .A2(n546), .A3(n547), .ZN(n185) );
  XNOR2_X1 U503 ( .A(n612), .B(n420), .ZN(n338) );
  INV_X1 U504 ( .A(n249), .ZN(n548) );
  INV_X2 U505 ( .A(n249), .ZN(n549) );
  BUF_X2 U506 ( .A(n9), .Z(n597) );
  XOR2_X1 U507 ( .A(n193), .B(n282), .Z(n551) );
  NAND2_X1 U508 ( .A1(n191), .A2(n193), .ZN(n552) );
  NAND2_X1 U509 ( .A1(n191), .A2(n282), .ZN(n553) );
  NAND2_X1 U510 ( .A1(n193), .A2(n282), .ZN(n554) );
  NAND3_X1 U511 ( .A1(n552), .A2(n553), .A3(n554), .ZN(n179) );
  XNOR2_X1 U512 ( .A(n609), .B(a[8]), .ZN(n555) );
  INV_X1 U513 ( .A(n564), .ZN(n32) );
  OR2_X1 U514 ( .A1(n78), .A2(n563), .ZN(n556) );
  XOR2_X1 U515 ( .A(n299), .B(n256), .Z(n557) );
  XOR2_X1 U516 ( .A(n230), .B(n557), .Z(n228) );
  NAND2_X1 U517 ( .A1(n529), .A2(n299), .ZN(n558) );
  NAND2_X1 U518 ( .A1(n529), .A2(n256), .ZN(n559) );
  NAND2_X1 U519 ( .A1(n299), .A2(n256), .ZN(n560) );
  NAND3_X1 U520 ( .A1(n558), .A2(n559), .A3(n560), .ZN(n227) );
  XNOR2_X1 U521 ( .A(n571), .B(n561), .ZN(product[9]) );
  AND2_X1 U522 ( .A1(n538), .A2(n90), .ZN(n561) );
  AOI21_X1 U523 ( .B1(n505), .B2(n587), .A(n93), .ZN(n562) );
  NOR2_X1 U524 ( .A1(n164), .A2(n175), .ZN(n563) );
  NOR2_X1 U525 ( .A1(n164), .A2(n175), .ZN(n75) );
  XNOR2_X1 U526 ( .A(n611), .B(a[10]), .ZN(n564) );
  NAND2_X1 U527 ( .A1(n214), .A2(n216), .ZN(n565) );
  NAND2_X1 U528 ( .A1(n214), .A2(n219), .ZN(n566) );
  NAND2_X1 U529 ( .A1(n216), .A2(n219), .ZN(n567) );
  NAND3_X1 U530 ( .A1(n565), .A2(n566), .A3(n567), .ZN(n211) );
  NOR2_X1 U531 ( .A1(n583), .A2(n402), .ZN(n568) );
  NOR2_X1 U532 ( .A1(n401), .A2(n549), .ZN(n569) );
  OR2_X1 U533 ( .A1(n568), .A2(n569), .ZN(n323) );
  XNOR2_X1 U534 ( .A(n607), .B(a[6]), .ZN(n570) );
  AOI21_X1 U535 ( .B1(n96), .B2(n587), .A(n93), .ZN(n91) );
  NAND2_X1 U536 ( .A1(n226), .A2(n229), .ZN(n572) );
  NAND2_X1 U537 ( .A1(n226), .A2(n298), .ZN(n573) );
  NAND2_X1 U538 ( .A1(n229), .A2(n298), .ZN(n574) );
  NAND3_X1 U539 ( .A1(n572), .A2(n573), .A3(n574), .ZN(n223) );
  BUF_X1 U540 ( .A(n12), .Z(n576) );
  XNOR2_X1 U541 ( .A(n604), .B(a[4]), .ZN(n575) );
  BUF_X2 U542 ( .A(n12), .Z(n577) );
  NAND2_X1 U543 ( .A1(n9), .A2(n585), .ZN(n12) );
  INV_X1 U544 ( .A(n580), .ZN(n103) );
  AND2_X1 U545 ( .A1(n224), .A2(n227), .ZN(n580) );
  NOR2_X1 U546 ( .A1(n186), .A2(n195), .ZN(n578) );
  NOR2_X1 U547 ( .A1(n186), .A2(n195), .ZN(n82) );
  CLKBUF_X1 U548 ( .A(n107), .Z(n579) );
  OR2_X1 U549 ( .A1(n228), .A2(n231), .ZN(n581) );
  NAND2_X2 U550 ( .A1(n431), .A2(n531), .ZN(n18) );
  NAND2_X1 U551 ( .A1(n525), .A2(n548), .ZN(n582) );
  NAND2_X1 U552 ( .A1(n525), .A2(n548), .ZN(n6) );
  AOI21_X1 U553 ( .B1(n598), .B2(n80), .A(n81), .ZN(n584) );
  OR2_X1 U554 ( .A1(n152), .A2(n163), .ZN(n586) );
  INV_X2 U555 ( .A(n609), .ZN(n608) );
  INV_X1 U556 ( .A(n69), .ZN(n67) );
  NAND2_X1 U557 ( .A1(n586), .A2(n69), .ZN(n47) );
  INV_X1 U558 ( .A(n74), .ZN(n72) );
  NAND2_X1 U559 ( .A1(n73), .A2(n586), .ZN(n64) );
  INV_X1 U560 ( .A(n95), .ZN(n93) );
  AOI21_X1 U561 ( .B1(n80), .B2(n598), .A(n81), .ZN(n45) );
  NOR2_X1 U562 ( .A1(n578), .A2(n85), .ZN(n80) );
  INV_X1 U563 ( .A(n78), .ZN(n126) );
  NAND2_X1 U564 ( .A1(n587), .A2(n95), .ZN(n53) );
  OAI21_X1 U565 ( .B1(n75), .B2(n79), .A(n76), .ZN(n74) );
  NAND2_X1 U566 ( .A1(n530), .A2(n528), .ZN(n51) );
  NAND2_X1 U567 ( .A1(n125), .A2(n76), .ZN(n48) );
  INV_X1 U568 ( .A(n543), .ZN(n125) );
  XNOR2_X1 U569 ( .A(n84), .B(n50), .ZN(product[11]) );
  NAND2_X1 U570 ( .A1(n127), .A2(n83), .ZN(n50) );
  INV_X1 U571 ( .A(n578), .ZN(n127) );
  NAND2_X1 U572 ( .A1(n152), .A2(n163), .ZN(n69) );
  OAI21_X1 U573 ( .B1(n113), .B2(n115), .A(n114), .ZN(n112) );
  INV_X1 U574 ( .A(n113), .ZN(n135) );
  NAND2_X1 U575 ( .A1(n581), .A2(n106), .ZN(n56) );
  NAND2_X1 U576 ( .A1(n492), .A2(n98), .ZN(n54) );
  AOI21_X1 U577 ( .B1(n589), .B2(n112), .A(n493), .ZN(n107) );
  NOR2_X1 U578 ( .A1(n176), .A2(n185), .ZN(n78) );
  NOR2_X1 U579 ( .A1(n196), .A2(n203), .ZN(n85) );
  NAND2_X1 U580 ( .A1(n590), .A2(n103), .ZN(n55) );
  NAND2_X1 U581 ( .A1(n589), .A2(n111), .ZN(n57) );
  AOI21_X1 U582 ( .B1(n588), .B2(n120), .A(n117), .ZN(n115) );
  INV_X1 U583 ( .A(n119), .ZN(n117) );
  INV_X1 U584 ( .A(n122), .ZN(n120) );
  XNOR2_X1 U585 ( .A(n63), .B(n46), .ZN(product[15]) );
  NAND2_X1 U586 ( .A1(n591), .A2(n62), .ZN(n46) );
  AOI21_X1 U587 ( .B1(n74), .B2(n586), .A(n67), .ZN(n65) );
  XNOR2_X1 U588 ( .A(n59), .B(n120), .ZN(product[2]) );
  NAND2_X1 U589 ( .A1(n588), .A2(n119), .ZN(n59) );
  NAND2_X1 U590 ( .A1(n176), .A2(n185), .ZN(n79) );
  NAND2_X1 U591 ( .A1(n524), .A2(n203), .ZN(n86) );
  NAND2_X1 U592 ( .A1(n164), .A2(n175), .ZN(n76) );
  NAND2_X1 U593 ( .A1(n186), .A2(n195), .ZN(n83) );
  NAND2_X1 U594 ( .A1(n204), .A2(n211), .ZN(n90) );
  NAND2_X1 U595 ( .A1(n212), .A2(n217), .ZN(n95) );
  OR2_X1 U596 ( .A1(n212), .A2(n217), .ZN(n587) );
  NAND2_X1 U597 ( .A1(n328), .A2(n314), .ZN(n119) );
  OR2_X1 U598 ( .A1(n328), .A2(n314), .ZN(n588) );
  NOR2_X1 U599 ( .A1(n228), .A2(n231), .ZN(n105) );
  NOR2_X1 U600 ( .A1(n218), .A2(n223), .ZN(n97) );
  OR2_X1 U601 ( .A1(n232), .A2(n233), .ZN(n589) );
  NAND2_X1 U602 ( .A1(n218), .A2(n223), .ZN(n98) );
  NAND2_X1 U603 ( .A1(n228), .A2(n231), .ZN(n106) );
  NAND2_X1 U604 ( .A1(n232), .A2(n233), .ZN(n111) );
  OR2_X1 U605 ( .A1(n224), .A2(n227), .ZN(n590) );
  INV_X1 U606 ( .A(n41), .ZN(n235) );
  OR2_X1 U607 ( .A1(n151), .A2(n139), .ZN(n591) );
  AND2_X1 U608 ( .A1(n496), .A2(n122), .ZN(product[1]) );
  XNOR2_X1 U609 ( .A(n614), .B(a[14]), .ZN(n41) );
  OR2_X1 U610 ( .A1(n599), .A2(n604), .ZN(n392) );
  OAI22_X1 U611 ( .A1(n39), .A2(n336), .B1(n37), .B2(n335), .ZN(n263) );
  AND2_X1 U612 ( .A1(n600), .A2(n570), .ZN(n288) );
  XNOR2_X1 U613 ( .A(n606), .B(n599), .ZN(n376) );
  AND2_X1 U614 ( .A1(n600), .A2(n575), .ZN(n300) );
  XNOR2_X1 U615 ( .A(n500), .B(n599), .ZN(n352) );
  OAI22_X1 U616 ( .A1(n39), .A2(n615), .B1(n337), .B2(n37), .ZN(n252) );
  OR2_X1 U617 ( .A1(n599), .A2(n615), .ZN(n337) );
  OAI22_X1 U618 ( .A1(n42), .A2(n617), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U619 ( .A1(n599), .A2(n617), .ZN(n332) );
  XNOR2_X1 U620 ( .A(n612), .B(n599), .ZN(n343) );
  XNOR2_X1 U621 ( .A(n155), .B(n593), .ZN(n139) );
  XNOR2_X1 U622 ( .A(n153), .B(n141), .ZN(n593) );
  XNOR2_X1 U623 ( .A(n157), .B(n594), .ZN(n141) );
  XNOR2_X1 U624 ( .A(n145), .B(n143), .ZN(n594) );
  XNOR2_X1 U625 ( .A(n159), .B(n595), .ZN(n142) );
  XNOR2_X1 U626 ( .A(n315), .B(n261), .ZN(n595) );
  XNOR2_X1 U627 ( .A(n614), .B(n599), .ZN(n336) );
  AND2_X1 U628 ( .A1(n600), .A2(n247), .ZN(n314) );
  NAND2_X1 U629 ( .A1(n427), .A2(n37), .ZN(n39) );
  XOR2_X1 U630 ( .A(n614), .B(a[12]), .Z(n427) );
  AND2_X1 U631 ( .A1(n600), .A2(n522), .ZN(n264) );
  AND2_X1 U632 ( .A1(n600), .A2(n235), .ZN(n260) );
  OAI22_X1 U633 ( .A1(n39), .A2(n335), .B1(n37), .B2(n334), .ZN(n262) );
  AND2_X1 U634 ( .A1(n600), .A2(n564), .ZN(n270) );
  INV_X1 U635 ( .A(n25), .ZN(n611) );
  INV_X1 U636 ( .A(n19), .ZN(n609) );
  AND2_X1 U637 ( .A1(n600), .A2(n555), .ZN(n278) );
  INV_X1 U638 ( .A(n1), .ZN(n602) );
  NAND2_X1 U639 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U640 ( .A(n616), .B(a[14]), .Z(n426) );
  INV_X1 U641 ( .A(n7), .ZN(n604) );
  XNOR2_X1 U642 ( .A(n608), .B(n599), .ZN(n363) );
  AND2_X1 U643 ( .A1(n600), .A2(n249), .ZN(product[0]) );
  OR2_X1 U644 ( .A1(n599), .A2(n613), .ZN(n344) );
  OR2_X1 U645 ( .A1(n599), .A2(n609), .ZN(n364) );
  OR2_X1 U646 ( .A1(n599), .A2(n611), .ZN(n353) );
  OR2_X1 U647 ( .A1(n599), .A2(n607), .ZN(n377) );
  BUF_X2 U648 ( .A(n43), .Z(n599) );
  XNOR2_X1 U649 ( .A(n608), .B(b[9]), .ZN(n354) );
  OAI22_X1 U650 ( .A1(n39), .A2(n334), .B1(n37), .B2(n333), .ZN(n261) );
  XNOR2_X1 U651 ( .A(n614), .B(n422), .ZN(n333) );
  XNOR2_X1 U652 ( .A(n606), .B(b[11]), .ZN(n365) );
  XNOR2_X1 U653 ( .A(n614), .B(n424), .ZN(n335) );
  XNOR2_X1 U654 ( .A(n614), .B(n423), .ZN(n334) );
  OAI22_X1 U655 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U656 ( .A(n616), .B(n424), .ZN(n330) );
  XNOR2_X1 U657 ( .A(n616), .B(n599), .ZN(n331) );
  XNOR2_X1 U658 ( .A(n500), .B(n418), .ZN(n345) );
  XNOR2_X1 U659 ( .A(n265), .B(n596), .ZN(n145) );
  XNOR2_X1 U660 ( .A(n149), .B(n147), .ZN(n596) );
  XNOR2_X1 U661 ( .A(n603), .B(b[13]), .ZN(n378) );
  XNOR2_X1 U662 ( .A(n500), .B(n424), .ZN(n351) );
  XNOR2_X1 U663 ( .A(n612), .B(n424), .ZN(n342) );
  XNOR2_X1 U664 ( .A(n608), .B(n424), .ZN(n362) );
  XNOR2_X1 U665 ( .A(n612), .B(n422), .ZN(n340) );
  XNOR2_X1 U666 ( .A(n612), .B(n421), .ZN(n339) );
  XNOR2_X1 U667 ( .A(n612), .B(n423), .ZN(n341) );
  XNOR2_X1 U668 ( .A(n603), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U669 ( .A(n603), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U670 ( .A(n603), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U671 ( .A(n603), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U672 ( .A(n603), .B(n418), .ZN(n384) );
  XNOR2_X1 U673 ( .A(n603), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U674 ( .A(n603), .B(n419), .ZN(n385) );
  XNOR2_X1 U675 ( .A(n608), .B(n423), .ZN(n361) );
  XNOR2_X1 U676 ( .A(n500), .B(n423), .ZN(n350) );
  XNOR2_X1 U677 ( .A(n606), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U678 ( .A(n606), .B(n418), .ZN(n369) );
  XNOR2_X1 U679 ( .A(n606), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U680 ( .A(n606), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U681 ( .A(n608), .B(n422), .ZN(n360) );
  XNOR2_X1 U682 ( .A(n500), .B(n422), .ZN(n349) );
  XNOR2_X1 U683 ( .A(n500), .B(n420), .ZN(n347) );
  XNOR2_X1 U684 ( .A(n608), .B(n420), .ZN(n358) );
  XNOR2_X1 U685 ( .A(n507), .B(b[14]), .ZN(n394) );
  XNOR2_X1 U686 ( .A(n506), .B(b[13]), .ZN(n395) );
  XNOR2_X1 U687 ( .A(n506), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U688 ( .A(n506), .B(b[11]), .ZN(n397) );
  XNOR2_X1 U689 ( .A(n500), .B(n421), .ZN(n348) );
  XNOR2_X1 U690 ( .A(n608), .B(n421), .ZN(n359) );
  XNOR2_X1 U691 ( .A(n500), .B(n419), .ZN(n346) );
  XNOR2_X1 U692 ( .A(n608), .B(n419), .ZN(n357) );
  XNOR2_X1 U693 ( .A(n608), .B(n418), .ZN(n356) );
  XNOR2_X1 U694 ( .A(n608), .B(b[8]), .ZN(n355) );
  BUF_X1 U695 ( .A(n43), .Z(n600) );
  XNOR2_X1 U696 ( .A(n506), .B(b[15]), .ZN(n393) );
  OAI22_X1 U697 ( .A1(n34), .A2(n339), .B1(n338), .B2(n539), .ZN(n265) );
  OAI22_X1 U698 ( .A1(n34), .A2(n340), .B1(n339), .B2(n539), .ZN(n266) );
  OAI22_X1 U699 ( .A1(n34), .A2(n342), .B1(n341), .B2(n32), .ZN(n268) );
  OAI22_X1 U700 ( .A1(n34), .A2(n341), .B1(n340), .B2(n32), .ZN(n267) );
  OAI22_X1 U701 ( .A1(n34), .A2(n343), .B1(n342), .B2(n32), .ZN(n269) );
  OAI22_X1 U702 ( .A1(n34), .A2(n613), .B1(n344), .B2(n32), .ZN(n253) );
  OAI21_X1 U703 ( .B1(n562), .B2(n89), .A(n90), .ZN(n598) );
  XNOR2_X1 U704 ( .A(n88), .B(n51), .ZN(product[10]) );
  OAI21_X1 U705 ( .B1(n89), .B2(n91), .A(n90), .ZN(n88) );
  XNOR2_X1 U706 ( .A(n70), .B(n47), .ZN(product[14]) );
  NOR2_X1 U707 ( .A1(n204), .A2(n211), .ZN(n89) );
  OAI22_X1 U708 ( .A1(n29), .A2(n346), .B1(n345), .B2(n497), .ZN(n271) );
  OAI22_X1 U709 ( .A1(n29), .A2(n350), .B1(n349), .B2(n497), .ZN(n275) );
  OAI22_X1 U710 ( .A1(n29), .A2(n347), .B1(n346), .B2(n497), .ZN(n272) );
  OAI22_X1 U711 ( .A1(n29), .A2(n348), .B1(n347), .B2(n497), .ZN(n273) );
  OAI22_X1 U712 ( .A1(n29), .A2(n349), .B1(n348), .B2(n497), .ZN(n274) );
  OAI22_X1 U713 ( .A1(n29), .A2(n611), .B1(n353), .B2(n497), .ZN(n254) );
  OAI22_X1 U714 ( .A1(n29), .A2(n351), .B1(n350), .B2(n497), .ZN(n276) );
  OAI22_X1 U715 ( .A1(n29), .A2(n352), .B1(n351), .B2(n497), .ZN(n277) );
  NOR2_X1 U716 ( .A1(n234), .A2(n257), .ZN(n113) );
  NAND2_X1 U717 ( .A1(n135), .A2(n114), .ZN(n58) );
  OAI21_X1 U718 ( .B1(n503), .B2(n97), .A(n98), .ZN(n96) );
  OR2_X1 U719 ( .A1(n599), .A2(n535), .ZN(n409) );
  XNOR2_X1 U720 ( .A(n77), .B(n48), .ZN(product[13]) );
  OAI22_X1 U721 ( .A1(n540), .A2(n358), .B1(n357), .B2(n21), .ZN(n282) );
  OAI22_X1 U722 ( .A1(n540), .A2(n362), .B1(n361), .B2(n21), .ZN(n286) );
  OAI22_X1 U723 ( .A1(n23), .A2(n356), .B1(n355), .B2(n21), .ZN(n280) );
  OAI22_X1 U724 ( .A1(n23), .A2(n355), .B1(n354), .B2(n21), .ZN(n279) );
  OAI22_X1 U725 ( .A1(n23), .A2(n609), .B1(n364), .B2(n21), .ZN(n255) );
  OAI22_X1 U726 ( .A1(n23), .A2(n360), .B1(n359), .B2(n21), .ZN(n284) );
  OAI22_X1 U727 ( .A1(n540), .A2(n361), .B1(n360), .B2(n21), .ZN(n285) );
  OAI22_X1 U728 ( .A1(n540), .A2(n363), .B1(n362), .B2(n21), .ZN(n287) );
  OAI22_X1 U729 ( .A1(n540), .A2(n357), .B1(n356), .B2(n21), .ZN(n281) );
  XNOR2_X1 U730 ( .A(n605), .B(n424), .ZN(n375) );
  XNOR2_X1 U731 ( .A(n605), .B(n421), .ZN(n372) );
  XNOR2_X1 U732 ( .A(n605), .B(n423), .ZN(n374) );
  OAI22_X1 U733 ( .A1(n23), .A2(n359), .B1(n358), .B2(n21), .ZN(n283) );
  XNOR2_X1 U734 ( .A(n605), .B(n422), .ZN(n373) );
  XNOR2_X1 U735 ( .A(n605), .B(n419), .ZN(n370) );
  XNOR2_X1 U736 ( .A(n605), .B(n420), .ZN(n371) );
  XNOR2_X1 U737 ( .A(n55), .B(n527), .ZN(product[6]) );
  OAI21_X1 U738 ( .B1(n107), .B2(n105), .A(n106), .ZN(n104) );
  NAND2_X1 U739 ( .A1(n151), .A2(n139), .ZN(n62) );
  OAI22_X1 U740 ( .A1(n18), .A2(n370), .B1(n369), .B2(n16), .ZN(n293) );
  OAI22_X1 U741 ( .A1(n18), .A2(n375), .B1(n374), .B2(n16), .ZN(n298) );
  OAI22_X1 U742 ( .A1(n18), .A2(n367), .B1(n366), .B2(n16), .ZN(n290) );
  OAI22_X1 U743 ( .A1(n18), .A2(n372), .B1(n371), .B2(n16), .ZN(n295) );
  OAI22_X1 U744 ( .A1(n18), .A2(n607), .B1(n377), .B2(n16), .ZN(n256) );
  OAI22_X1 U745 ( .A1(n18), .A2(n368), .B1(n367), .B2(n16), .ZN(n291) );
  OAI22_X1 U746 ( .A1(n18), .A2(n376), .B1(n375), .B2(n16), .ZN(n299) );
  OAI22_X1 U747 ( .A1(n18), .A2(n374), .B1(n373), .B2(n16), .ZN(n297) );
  OAI22_X1 U748 ( .A1(n18), .A2(n369), .B1(n368), .B2(n16), .ZN(n292) );
  OAI22_X1 U749 ( .A1(n18), .A2(n373), .B1(n372), .B2(n16), .ZN(n296) );
  OAI22_X1 U750 ( .A1(n18), .A2(n371), .B1(n370), .B2(n16), .ZN(n294) );
  OAI22_X1 U751 ( .A1(n18), .A2(n366), .B1(n365), .B2(n16), .ZN(n289) );
  XNOR2_X1 U752 ( .A(n534), .B(n420), .ZN(n386) );
  XNOR2_X1 U753 ( .A(n534), .B(n422), .ZN(n388) );
  XNOR2_X1 U754 ( .A(n534), .B(n599), .ZN(n391) );
  XNOR2_X1 U755 ( .A(n534), .B(n421), .ZN(n387) );
  XNOR2_X1 U756 ( .A(n534), .B(n423), .ZN(n389) );
  XNOR2_X1 U757 ( .A(n534), .B(n424), .ZN(n390) );
  XNOR2_X1 U758 ( .A(n507), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U759 ( .A(n507), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U760 ( .A(n506), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U761 ( .A(n506), .B(n418), .ZN(n401) );
  XNOR2_X1 U762 ( .A(n507), .B(n420), .ZN(n403) );
  XNOR2_X1 U763 ( .A(n507), .B(n599), .ZN(n408) );
  XNOR2_X1 U764 ( .A(n507), .B(n419), .ZN(n402) );
  XNOR2_X1 U765 ( .A(n513), .B(n421), .ZN(n404) );
  XNOR2_X1 U766 ( .A(n513), .B(n422), .ZN(n405) );
  XNOR2_X1 U767 ( .A(n506), .B(n424), .ZN(n407) );
  XNOR2_X1 U768 ( .A(n507), .B(n423), .ZN(n406) );
  OAI21_X1 U769 ( .B1(n87), .B2(n514), .A(n490), .ZN(n84) );
  XOR2_X1 U770 ( .A(n56), .B(n579), .Z(product[5]) );
  OAI21_X1 U771 ( .B1(n64), .B2(n495), .A(n65), .ZN(n63) );
  OAI21_X1 U772 ( .B1(n584), .B2(n523), .A(n79), .ZN(n77) );
  OAI21_X1 U773 ( .B1(n584), .B2(n556), .A(n72), .ZN(n70) );
  INV_X1 U774 ( .A(n88), .ZN(n87) );
  XNOR2_X1 U775 ( .A(n57), .B(n112), .ZN(product[4]) );
  XNOR2_X1 U776 ( .A(n505), .B(n53), .ZN(product[8]) );
  XOR2_X1 U777 ( .A(n58), .B(n542), .Z(product[3]) );
  OAI22_X1 U778 ( .A1(n6), .A2(n395), .B1(n394), .B2(n549), .ZN(n316) );
  OAI22_X1 U779 ( .A1(n583), .A2(n394), .B1(n393), .B2(n549), .ZN(n315) );
  OAI22_X1 U780 ( .A1(n583), .A2(n396), .B1(n395), .B2(n549), .ZN(n317) );
  OAI22_X1 U781 ( .A1(n582), .A2(n397), .B1(n396), .B2(n549), .ZN(n318) );
  OAI22_X1 U782 ( .A1(n583), .A2(n398), .B1(n397), .B2(n549), .ZN(n319) );
  OAI22_X1 U783 ( .A1(n583), .A2(n400), .B1(n399), .B2(n549), .ZN(n321) );
  OAI22_X1 U784 ( .A1(n6), .A2(n399), .B1(n398), .B2(n549), .ZN(n320) );
  OAI22_X1 U785 ( .A1(n401), .A2(n582), .B1(n400), .B2(n549), .ZN(n322) );
  NAND2_X1 U786 ( .A1(n329), .A2(n258), .ZN(n122) );
  OAI22_X1 U787 ( .A1(n6), .A2(n404), .B1(n403), .B2(n549), .ZN(n325) );
  OAI22_X1 U788 ( .A1(n582), .A2(n403), .B1(n402), .B2(n549), .ZN(n324) );
  OAI22_X1 U789 ( .A1(n582), .A2(n406), .B1(n405), .B2(n549), .ZN(n327) );
  OAI22_X1 U790 ( .A1(n6), .A2(n405), .B1(n404), .B2(n549), .ZN(n326) );
  OAI22_X1 U791 ( .A1(n582), .A2(n407), .B1(n406), .B2(n549), .ZN(n328) );
  OAI22_X1 U792 ( .A1(n583), .A2(n408), .B1(n407), .B2(n549), .ZN(n329) );
  OAI22_X1 U793 ( .A1(n583), .A2(n535), .B1(n409), .B2(n549), .ZN(n258) );
  XOR2_X1 U794 ( .A(n541), .B(n54), .Z(product[7]) );
  OAI22_X1 U795 ( .A1(n577), .A2(n379), .B1(n378), .B2(n533), .ZN(n301) );
  OAI22_X1 U796 ( .A1(n577), .A2(n380), .B1(n379), .B2(n597), .ZN(n302) );
  OAI22_X1 U797 ( .A1(n577), .A2(n385), .B1(n384), .B2(n533), .ZN(n307) );
  OAI22_X1 U798 ( .A1(n577), .A2(n382), .B1(n381), .B2(n597), .ZN(n304) );
  OAI22_X1 U799 ( .A1(n577), .A2(n381), .B1(n380), .B2(n597), .ZN(n303) );
  NAND2_X1 U800 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U801 ( .A1(n576), .A2(n383), .B1(n597), .B2(n382), .ZN(n305) );
  OAI22_X1 U802 ( .A1(n576), .A2(n384), .B1(n597), .B2(n383), .ZN(n306) );
  OAI22_X1 U803 ( .A1(n577), .A2(n386), .B1(n385), .B2(n597), .ZN(n308) );
  OAI22_X1 U804 ( .A1(n577), .A2(n387), .B1(n386), .B2(n597), .ZN(n309) );
  OAI22_X1 U805 ( .A1(n577), .A2(n536), .B1(n392), .B2(n597), .ZN(n257) );
  OAI22_X1 U806 ( .A1(n577), .A2(n389), .B1(n388), .B2(n597), .ZN(n311) );
  OAI22_X1 U807 ( .A1(n577), .A2(n388), .B1(n387), .B2(n597), .ZN(n310) );
  OAI22_X1 U808 ( .A1(n576), .A2(n390), .B1(n597), .B2(n389), .ZN(n312) );
  INV_X1 U809 ( .A(n597), .ZN(n247) );
  OAI22_X1 U810 ( .A1(n577), .A2(n391), .B1(n390), .B2(n597), .ZN(n313) );
  INV_X1 U811 ( .A(n537), .ZN(n603) );
  INV_X1 U812 ( .A(n607), .ZN(n606) );
  INV_X1 U813 ( .A(n31), .ZN(n613) );
  INV_X1 U814 ( .A(n615), .ZN(n614) );
  INV_X1 U815 ( .A(n36), .ZN(n615) );
  INV_X1 U816 ( .A(n617), .ZN(n616) );
  INV_X1 U817 ( .A(n40), .ZN(n617) );
  XOR2_X1 U818 ( .A(n259), .B(n251), .Z(n148) );
  XOR2_X1 U819 ( .A(n289), .B(n279), .Z(n146) );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_0_DW01_add_2 ( A, B, CI, 
        SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n19, n20, n22, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n44, n45, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n65, n67, n68, n69, n70,
         n71, n73, n75, n76, n77, n78, n79, n81, n83, n84, n86, n88, n89, n91,
         n94, n95, n96, n98, n100, n157, n158, n159, n160, n161, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177;

  AOI21_X1 U122 ( .B1(n52), .B2(n60), .A(n53), .ZN(n51) );
  NOR2_X1 U123 ( .A1(A[11]), .A2(B[11]), .ZN(n157) );
  NOR2_X1 U124 ( .A1(A[11]), .A2(B[11]), .ZN(n35) );
  OR2_X2 U125 ( .A1(A[9]), .A2(B[9]), .ZN(n173) );
  AND2_X1 U126 ( .A1(A[9]), .A2(B[9]), .ZN(n158) );
  BUF_X1 U127 ( .A(n158), .Z(n159) );
  OR2_X1 U128 ( .A1(A[12]), .A2(B[12]), .ZN(n160) );
  OR2_X1 U129 ( .A1(A[15]), .A2(B[15]), .ZN(n161) );
  AND2_X1 U130 ( .A1(n171), .A2(n86), .ZN(SUM[0]) );
  NOR2_X1 U131 ( .A1(A[8]), .A2(B[8]), .ZN(n163) );
  NOR2_X1 U132 ( .A1(A[8]), .A2(B[8]), .ZN(n54) );
  AOI21_X1 U133 ( .B1(n158), .B2(n177), .A(n170), .ZN(n164) );
  NOR2_X1 U134 ( .A1(A[14]), .A2(B[14]), .ZN(n165) );
  NOR2_X1 U135 ( .A1(A[14]), .A2(B[14]), .ZN(n25) );
  OAI21_X1 U136 ( .B1(n51), .B2(n39), .A(n164), .ZN(n166) );
  AOI21_X1 U137 ( .B1(n166), .B2(n30), .A(n31), .ZN(n167) );
  AOI21_X1 U138 ( .B1(n166), .B2(n30), .A(n31), .ZN(n1) );
  OR2_X1 U139 ( .A1(A[10]), .A2(B[10]), .ZN(n168) );
  INV_X1 U140 ( .A(n170), .ZN(n44) );
  NOR2_X1 U141 ( .A1(A[12]), .A2(B[12]), .ZN(n169) );
  NOR2_X1 U142 ( .A1(A[12]), .A2(B[12]), .ZN(n32) );
  AND2_X1 U143 ( .A1(A[10]), .A2(B[10]), .ZN(n170) );
  OR2_X1 U144 ( .A1(A[0]), .A2(B[0]), .ZN(n171) );
  INV_X1 U145 ( .A(n60), .ZN(n59) );
  INV_X1 U146 ( .A(n51), .ZN(n50) );
  INV_X1 U147 ( .A(n67), .ZN(n65) );
  AOI21_X1 U148 ( .B1(n174), .B2(n84), .A(n81), .ZN(n79) );
  INV_X1 U149 ( .A(n83), .ZN(n81) );
  AOI21_X1 U150 ( .B1(n175), .B2(n76), .A(n73), .ZN(n71) );
  INV_X1 U151 ( .A(n75), .ZN(n73) );
  OR2_X1 U152 ( .A1(n25), .A2(n28), .ZN(n172) );
  OAI21_X1 U153 ( .B1(n79), .B2(n77), .A(n78), .ZN(n76) );
  AOI21_X1 U154 ( .B1(n50), .B2(n173), .A(n159), .ZN(n45) );
  NAND2_X1 U155 ( .A1(n94), .A2(n55), .ZN(n9) );
  INV_X1 U156 ( .A(n86), .ZN(n84) );
  OAI21_X1 U157 ( .B1(n59), .B2(n57), .A(n58), .ZN(n56) );
  NAND2_X1 U158 ( .A1(n100), .A2(n78), .ZN(n15) );
  INV_X1 U159 ( .A(n77), .ZN(n100) );
  INV_X1 U160 ( .A(n157), .ZN(n91) );
  INV_X1 U161 ( .A(n28), .ZN(n89) );
  NAND2_X1 U162 ( .A1(n173), .A2(n49), .ZN(n8) );
  NAND2_X1 U163 ( .A1(n95), .A2(n58), .ZN(n10) );
  INV_X1 U164 ( .A(n57), .ZN(n95) );
  NAND2_X1 U165 ( .A1(n176), .A2(n67), .ZN(n12) );
  NAND2_X1 U166 ( .A1(n175), .A2(n75), .ZN(n14) );
  NAND2_X1 U167 ( .A1(n174), .A2(n83), .ZN(n16) );
  NAND2_X1 U168 ( .A1(n96), .A2(n62), .ZN(n11) );
  INV_X1 U169 ( .A(n61), .ZN(n96) );
  NAND2_X1 U170 ( .A1(n98), .A2(n70), .ZN(n13) );
  INV_X1 U171 ( .A(n69), .ZN(n98) );
  XNOR2_X1 U172 ( .A(n34), .B(n5), .ZN(SUM[12]) );
  NAND2_X1 U173 ( .A1(n160), .A2(n33), .ZN(n5) );
  XOR2_X1 U174 ( .A(n59), .B(n10), .Z(SUM[7]) );
  XNOR2_X1 U175 ( .A(n12), .B(n68), .ZN(SUM[5]) );
  XNOR2_X1 U176 ( .A(n14), .B(n76), .ZN(SUM[3]) );
  XOR2_X1 U177 ( .A(n15), .B(n79), .Z(SUM[2]) );
  XNOR2_X1 U178 ( .A(n16), .B(n84), .ZN(SUM[1]) );
  NOR2_X1 U179 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  NOR2_X1 U180 ( .A1(A[7]), .A2(B[7]), .ZN(n57) );
  NAND2_X1 U181 ( .A1(n91), .A2(n36), .ZN(n6) );
  NAND2_X1 U182 ( .A1(n89), .A2(n29), .ZN(n4) );
  NOR2_X1 U183 ( .A1(A[2]), .A2(B[2]), .ZN(n77) );
  NAND2_X1 U184 ( .A1(n88), .A2(n26), .ZN(n3) );
  XOR2_X1 U185 ( .A(n45), .B(n7), .Z(SUM[10]) );
  NAND2_X1 U186 ( .A1(A[11]), .A2(B[11]), .ZN(n36) );
  OR2_X1 U187 ( .A1(A[1]), .A2(B[1]), .ZN(n174) );
  XNOR2_X1 U188 ( .A(n56), .B(n9), .ZN(SUM[8]) );
  XNOR2_X1 U189 ( .A(n50), .B(n8), .ZN(SUM[9]) );
  NOR2_X1 U190 ( .A1(A[6]), .A2(B[6]), .ZN(n61) );
  NOR2_X1 U191 ( .A1(A[4]), .A2(B[4]), .ZN(n69) );
  NAND2_X1 U192 ( .A1(A[7]), .A2(B[7]), .ZN(n58) );
  OR2_X1 U193 ( .A1(A[3]), .A2(B[3]), .ZN(n175) );
  NAND2_X1 U194 ( .A1(A[2]), .A2(B[2]), .ZN(n78) );
  NAND2_X1 U195 ( .A1(A[5]), .A2(B[5]), .ZN(n67) );
  NAND2_X1 U196 ( .A1(A[1]), .A2(B[1]), .ZN(n83) );
  NAND2_X1 U197 ( .A1(A[3]), .A2(B[3]), .ZN(n75) );
  NAND2_X1 U198 ( .A1(A[0]), .A2(B[0]), .ZN(n86) );
  OR2_X1 U199 ( .A1(A[5]), .A2(B[5]), .ZN(n176) );
  NAND2_X1 U200 ( .A1(A[6]), .A2(B[6]), .ZN(n62) );
  NAND2_X1 U201 ( .A1(A[4]), .A2(B[4]), .ZN(n70) );
  NAND2_X1 U202 ( .A1(A[14]), .A2(B[14]), .ZN(n26) );
  OR2_X1 U203 ( .A1(A[10]), .A2(B[10]), .ZN(n177) );
  NAND2_X1 U204 ( .A1(n161), .A2(n19), .ZN(n2) );
  INV_X1 U205 ( .A(n163), .ZN(n94) );
  NOR2_X1 U206 ( .A1(n163), .A2(n57), .ZN(n52) );
  OAI21_X1 U207 ( .B1(n54), .B2(n58), .A(n55), .ZN(n53) );
  NAND2_X1 U208 ( .A1(A[8]), .A2(B[8]), .ZN(n55) );
  INV_X1 U209 ( .A(n24), .ZN(n22) );
  NAND2_X1 U210 ( .A1(A[9]), .A2(B[9]), .ZN(n49) );
  AOI21_X1 U211 ( .B1(n176), .B2(n68), .A(n65), .ZN(n63) );
  OAI21_X1 U212 ( .B1(n71), .B2(n69), .A(n70), .ZN(n68) );
  INV_X1 U213 ( .A(n25), .ZN(n88) );
  NOR2_X1 U214 ( .A1(n169), .A2(n35), .ZN(n30) );
  OAI21_X1 U215 ( .B1(n32), .B2(n36), .A(n33), .ZN(n31) );
  NAND2_X1 U216 ( .A1(A[13]), .A2(B[13]), .ZN(n29) );
  XOR2_X1 U217 ( .A(n37), .B(n6), .Z(SUM[11]) );
  OAI21_X1 U218 ( .B1(n37), .B2(n157), .A(n36), .ZN(n34) );
  NAND2_X1 U219 ( .A1(A[12]), .A2(B[12]), .ZN(n33) );
  OAI21_X1 U220 ( .B1(n165), .B2(n29), .A(n26), .ZN(n24) );
  INV_X1 U221 ( .A(n38), .ZN(n37) );
  OAI21_X1 U222 ( .B1(n39), .B2(n51), .A(n40), .ZN(n38) );
  AOI21_X1 U223 ( .B1(n158), .B2(n177), .A(n170), .ZN(n40) );
  NAND2_X1 U224 ( .A1(A[15]), .A2(B[15]), .ZN(n19) );
  XOR2_X1 U225 ( .A(n11), .B(n63), .Z(SUM[6]) );
  XOR2_X1 U226 ( .A(n13), .B(n71), .Z(SUM[4]) );
  OAI21_X1 U227 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  XNOR2_X1 U228 ( .A(n20), .B(n2), .ZN(SUM[15]) );
  NAND2_X1 U229 ( .A1(n168), .A2(n44), .ZN(n7) );
  NAND2_X1 U230 ( .A1(n168), .A2(n173), .ZN(n39) );
  XNOR2_X1 U231 ( .A(n27), .B(n3), .ZN(SUM[14]) );
  XOR2_X1 U232 ( .A(n167), .B(n4), .Z(SUM[13]) );
  OAI21_X1 U233 ( .B1(n1), .B2(n28), .A(n29), .ZN(n27) );
  OAI21_X1 U234 ( .B1(n1), .B2(n172), .A(n22), .ZN(n20) );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_0 ( clk, clear_acc, 
        data_out_x, data_out, data_out_w, data_out_b, wr_en_y, m_valid, 
        m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [4:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
         N39, N40, N41, N42, N43, N44, n30, n31, n84, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n103, n104,
         n105, n106, n107, n108, n109, n110, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n85, n102,
         n111, n112;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(clear_acc), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n101), .CK(clk), .Q(n25) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n100), .CK(clk), .Q(n26) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n99), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n98), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n94), .CK(clk), .Q(n34) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n93), .CK(clk), .Q(n35) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n92), .CK(clk), .Q(n36) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n91), .CK(clk), .Q(n37) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n90), .CK(clk), .Q(n38) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n89), .CK(clk), .Q(n39) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n88), .CK(clk), .Q(n40) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n87), .CK(clk), .Q(n41) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n86), .CK(clk), .Q(n42) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_0_DW_mult_tc_1 mult_2021 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_0_DW01_add_2 add_2022 ( .A({n127, 
        n128, n129, n130, n131, n132, n118, n119, n120, n121, n122, n123, n124, 
        n125, n126, n133}), .B({f[15], n46, n47, n48, n49, n51, f[9:0]}), .CI(
        1'b0), .SUM(adder) );
  DFF_X1 delay_reg ( .D(n112), .CK(clk), .Q(n17), .QN(n84) );
  DFF_X1 \data_out_reg[15]  ( .D(n165), .CK(clk), .Q(data_out[15]), .QN(n134)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n164), .CK(clk), .Q(data_out[14]), .QN(n135)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n163), .CK(clk), .Q(data_out[13]), .QN(n136)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n162), .CK(clk), .Q(data_out[12]), .QN(n137)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n161), .CK(clk), .Q(data_out[11]), .QN(n138)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n160), .CK(clk), .Q(data_out[10]), .QN(n139)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n159), .CK(clk), .Q(data_out[9]), .QN(n140) );
  DFF_X1 \data_out_reg[8]  ( .D(n158), .CK(clk), .Q(data_out[8]), .QN(n141) );
  DFF_X1 \data_out_reg[7]  ( .D(n157), .CK(clk), .Q(data_out[7]), .QN(n142) );
  DFF_X1 \data_out_reg[6]  ( .D(n156), .CK(clk), .Q(data_out[6]), .QN(n143) );
  DFF_X1 \data_out_reg[5]  ( .D(n155), .CK(clk), .Q(data_out[5]), .QN(n144) );
  DFF_X1 \data_out_reg[4]  ( .D(n154), .CK(clk), .Q(data_out[4]), .QN(n145) );
  DFF_X1 \data_out_reg[3]  ( .D(n153), .CK(clk), .Q(data_out[3]), .QN(n146) );
  DFF_X1 \data_out_reg[2]  ( .D(n152), .CK(clk), .Q(data_out[2]), .QN(n147) );
  DFF_X1 \data_out_reg[1]  ( .D(n151), .CK(clk), .Q(data_out[1]), .QN(n148) );
  DFF_X1 \data_out_reg[0]  ( .D(n150), .CK(clk), .Q(data_out[0]), .QN(n149) );
  DFF_X1 \f_reg[0]  ( .D(n111), .CK(clk), .Q(f[0]), .QN(n117) );
  DFF_X1 \f_reg[1]  ( .D(n102), .CK(clk), .Q(f[1]), .QN(n116) );
  DFF_X1 \f_reg[2]  ( .D(n85), .CK(clk), .Q(f[2]), .QN(n115) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n96), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n95), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n97), .CK(clk), .Q(n29) );
  DFF_X1 \f_reg[3]  ( .D(n83), .CK(clk), .Q(f[3]), .QN(n64) );
  DFF_X1 \f_reg[4]  ( .D(n82), .CK(clk), .Q(f[4]), .QN(n65) );
  DFF_X1 \f_reg[5]  ( .D(n81), .CK(clk), .Q(f[5]), .QN(n66) );
  DFF_X1 \f_reg[6]  ( .D(n80), .CK(clk), .Q(f[6]), .QN(n67) );
  DFF_X1 \f_reg[7]  ( .D(n79), .CK(clk), .Q(f[7]), .QN(n110) );
  DFF_X1 \f_reg[8]  ( .D(n78), .CK(clk), .Q(f[8]), .QN(n109) );
  DFF_X1 \f_reg[9]  ( .D(n77), .CK(clk), .Q(f[9]), .QN(n108) );
  DFF_X1 \f_reg[10]  ( .D(n76), .CK(clk), .Q(n51), .QN(n107) );
  DFF_X1 \f_reg[11]  ( .D(n75), .CK(clk), .Q(n49), .QN(n106) );
  DFF_X1 \f_reg[14]  ( .D(n12), .CK(clk), .Q(n46), .QN(n103) );
  DFF_X1 \f_reg[13]  ( .D(n2), .CK(clk), .Q(n47), .QN(n104) );
  DFF_X1 \f_reg[12]  ( .D(n4), .CK(clk), .Q(n48), .QN(n105) );
  DFF_X1 \f_reg[15]  ( .D(n8), .CK(clk), .Q(f[15]), .QN(n72) );
  MUX2_X2 U3 ( .A(N38), .B(n33), .S(n17), .Z(n118) );
  AND2_X1 U4 ( .A1(clear_acc_delay), .A2(n84), .ZN(n1) );
  AND2_X1 U5 ( .A1(n45), .A2(n23), .ZN(n21) );
  NAND3_X1 U6 ( .A1(n10), .A2(n9), .A3(n11), .ZN(n2) );
  MUX2_X2 U8 ( .A(n32), .B(N39), .S(n84), .Z(n132) );
  NAND3_X1 U9 ( .A1(n6), .A2(n5), .A3(n7), .ZN(n4) );
  NAND2_X1 U10 ( .A1(data_out_b[12]), .A2(clear_acc), .ZN(n5) );
  NAND2_X1 U11 ( .A1(adder[12]), .A2(n21), .ZN(n6) );
  NAND2_X1 U12 ( .A1(n62), .A2(n48), .ZN(n7) );
  INV_X1 U13 ( .A(n45), .ZN(n62) );
  NAND3_X1 U14 ( .A1(n13), .A2(n14), .A3(n15), .ZN(n8) );
  MUX2_X2 U15 ( .A(n27), .B(N42), .S(n84), .Z(n129) );
  NAND2_X1 U16 ( .A1(data_out_b[13]), .A2(clear_acc), .ZN(n9) );
  NAND2_X1 U17 ( .A1(adder[13]), .A2(n21), .ZN(n10) );
  NAND2_X1 U18 ( .A1(n62), .A2(n47), .ZN(n11) );
  NAND3_X1 U19 ( .A1(n19), .A2(n18), .A3(n20), .ZN(n12) );
  NAND2_X1 U20 ( .A1(data_out_b[15]), .A2(clear_acc), .ZN(n13) );
  NAND2_X1 U21 ( .A1(adder[15]), .A2(n21), .ZN(n14) );
  NAND2_X1 U22 ( .A1(n62), .A2(f[15]), .ZN(n15) );
  MUX2_X2 U23 ( .A(n34), .B(N37), .S(n84), .Z(n119) );
  MUX2_X2 U24 ( .A(n29), .B(N40), .S(n84), .Z(n131) );
  CLKBUF_X1 U25 ( .A(N43), .Z(n16) );
  MUX2_X2 U26 ( .A(N43), .B(n26), .S(n17), .Z(n128) );
  MUX2_X2 U27 ( .A(n28), .B(N41), .S(n84), .Z(n130) );
  NAND2_X1 U28 ( .A1(data_out_b[14]), .A2(clear_acc), .ZN(n18) );
  NAND2_X1 U29 ( .A1(adder[14]), .A2(n21), .ZN(n19) );
  NAND2_X1 U30 ( .A1(n62), .A2(n46), .ZN(n20) );
  NAND2_X1 U31 ( .A1(n112), .A2(n22), .ZN(n30) );
  INV_X1 U32 ( .A(clear_acc), .ZN(n23) );
  NAND3_X1 U33 ( .A1(wr_en_y), .A2(n73), .A3(n72), .ZN(n31) );
  OAI22_X1 U34 ( .A1(n146), .A2(n30), .B1(n64), .B2(n31), .ZN(n153) );
  OAI22_X1 U35 ( .A1(n145), .A2(n30), .B1(n65), .B2(n31), .ZN(n154) );
  OAI22_X1 U36 ( .A1(n144), .A2(n30), .B1(n66), .B2(n31), .ZN(n155) );
  OAI22_X1 U37 ( .A1(n143), .A2(n30), .B1(n67), .B2(n31), .ZN(n156) );
  OAI22_X1 U38 ( .A1(n142), .A2(n30), .B1(n110), .B2(n31), .ZN(n157) );
  OAI22_X1 U39 ( .A1(n141), .A2(n30), .B1(n109), .B2(n31), .ZN(n158) );
  OAI22_X1 U40 ( .A1(n140), .A2(n30), .B1(n108), .B2(n31), .ZN(n159) );
  INV_X1 U41 ( .A(wr_en_y), .ZN(n22) );
  INV_X1 U42 ( .A(m_ready), .ZN(n24) );
  NAND2_X1 U43 ( .A1(m_valid), .A2(n24), .ZN(n43) );
  OAI21_X1 U44 ( .B1(sel[4]), .B2(n74), .A(n43), .ZN(n112) );
  MUX2_X1 U45 ( .A(n25), .B(N44), .S(n1), .Z(n101) );
  MUX2_X1 U46 ( .A(n25), .B(N44), .S(n84), .Z(n127) );
  MUX2_X1 U47 ( .A(n26), .B(n16), .S(n1), .Z(n100) );
  MUX2_X1 U48 ( .A(n27), .B(N42), .S(n1), .Z(n99) );
  MUX2_X1 U49 ( .A(n28), .B(N41), .S(n1), .Z(n98) );
  MUX2_X1 U50 ( .A(n29), .B(N40), .S(n1), .Z(n97) );
  MUX2_X1 U51 ( .A(n32), .B(N39), .S(n1), .Z(n96) );
  MUX2_X1 U52 ( .A(n33), .B(N38), .S(n1), .Z(n95) );
  MUX2_X1 U53 ( .A(n34), .B(N37), .S(n1), .Z(n94) );
  MUX2_X1 U54 ( .A(n35), .B(N36), .S(n1), .Z(n93) );
  MUX2_X1 U55 ( .A(n35), .B(N36), .S(n84), .Z(n120) );
  MUX2_X1 U56 ( .A(n36), .B(N35), .S(n1), .Z(n92) );
  MUX2_X1 U57 ( .A(n36), .B(N35), .S(n84), .Z(n121) );
  MUX2_X1 U58 ( .A(n37), .B(N34), .S(n1), .Z(n91) );
  MUX2_X1 U59 ( .A(n37), .B(N34), .S(n84), .Z(n122) );
  MUX2_X1 U60 ( .A(n38), .B(N33), .S(n1), .Z(n90) );
  MUX2_X1 U61 ( .A(n38), .B(N33), .S(n84), .Z(n123) );
  MUX2_X1 U62 ( .A(n39), .B(N32), .S(n1), .Z(n89) );
  MUX2_X1 U63 ( .A(n39), .B(N32), .S(n84), .Z(n124) );
  MUX2_X1 U64 ( .A(n40), .B(N31), .S(n1), .Z(n88) );
  MUX2_X1 U65 ( .A(n40), .B(N31), .S(n84), .Z(n125) );
  MUX2_X1 U66 ( .A(n41), .B(N30), .S(n1), .Z(n87) );
  MUX2_X1 U67 ( .A(n41), .B(N30), .S(n84), .Z(n126) );
  MUX2_X1 U68 ( .A(n42), .B(N29), .S(n1), .Z(n86) );
  MUX2_X1 U69 ( .A(n42), .B(N29), .S(n84), .Z(n133) );
  INV_X1 U70 ( .A(n43), .ZN(n44) );
  OAI21_X1 U71 ( .B1(n44), .B2(n17), .A(n23), .ZN(n45) );
  AOI222_X1 U72 ( .A1(data_out_b[11]), .A2(clear_acc), .B1(adder[11]), .B2(n21), .C1(n62), .C2(n49), .ZN(n50) );
  INV_X1 U73 ( .A(n50), .ZN(n75) );
  AOI222_X1 U74 ( .A1(data_out_b[10]), .A2(clear_acc), .B1(adder[10]), .B2(n21), .C1(n62), .C2(n51), .ZN(n52) );
  INV_X1 U75 ( .A(n52), .ZN(n76) );
  AOI222_X1 U76 ( .A1(data_out_b[8]), .A2(clear_acc), .B1(adder[8]), .B2(n21), 
        .C1(n62), .C2(f[8]), .ZN(n53) );
  INV_X1 U77 ( .A(n53), .ZN(n78) );
  AOI222_X1 U78 ( .A1(data_out_b[7]), .A2(clear_acc), .B1(adder[7]), .B2(n21), 
        .C1(n62), .C2(f[7]), .ZN(n54) );
  INV_X1 U79 ( .A(n54), .ZN(n79) );
  AOI222_X1 U80 ( .A1(data_out_b[6]), .A2(clear_acc), .B1(adder[6]), .B2(n21), 
        .C1(n62), .C2(f[6]), .ZN(n55) );
  INV_X1 U81 ( .A(n55), .ZN(n80) );
  AOI222_X1 U82 ( .A1(data_out_b[5]), .A2(clear_acc), .B1(adder[5]), .B2(n21), 
        .C1(n62), .C2(f[5]), .ZN(n56) );
  INV_X1 U83 ( .A(n56), .ZN(n81) );
  AOI222_X1 U84 ( .A1(data_out_b[4]), .A2(clear_acc), .B1(adder[4]), .B2(n21), 
        .C1(n62), .C2(f[4]), .ZN(n57) );
  INV_X1 U85 ( .A(n57), .ZN(n82) );
  AOI222_X1 U86 ( .A1(data_out_b[3]), .A2(clear_acc), .B1(adder[3]), .B2(n21), 
        .C1(n62), .C2(f[3]), .ZN(n58) );
  INV_X1 U87 ( .A(n58), .ZN(n83) );
  AOI222_X1 U88 ( .A1(data_out_b[2]), .A2(clear_acc), .B1(adder[2]), .B2(n21), 
        .C1(n62), .C2(f[2]), .ZN(n59) );
  INV_X1 U89 ( .A(n59), .ZN(n85) );
  AOI222_X1 U90 ( .A1(data_out_b[1]), .A2(clear_acc), .B1(adder[1]), .B2(n21), 
        .C1(n62), .C2(f[1]), .ZN(n60) );
  INV_X1 U91 ( .A(n60), .ZN(n102) );
  AOI222_X1 U92 ( .A1(data_out_b[0]), .A2(clear_acc), .B1(adder[0]), .B2(n21), 
        .C1(n62), .C2(f[0]), .ZN(n61) );
  INV_X1 U93 ( .A(n61), .ZN(n111) );
  AOI222_X1 U94 ( .A1(data_out_b[9]), .A2(clear_acc), .B1(adder[9]), .B2(n21), 
        .C1(n62), .C2(f[9]), .ZN(n63) );
  INV_X1 U95 ( .A(n63), .ZN(n77) );
  NOR4_X1 U96 ( .A1(n49), .A2(n48), .A3(n47), .A4(n46), .ZN(n71) );
  NOR4_X1 U97 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n51), .ZN(n70) );
  NAND4_X1 U98 ( .A1(n67), .A2(n66), .A3(n65), .A4(n64), .ZN(n68) );
  NOR4_X1 U99 ( .A1(n68), .A2(f[0]), .A3(f[1]), .A4(f[2]), .ZN(n69) );
  NAND3_X1 U100 ( .A1(n71), .A2(n70), .A3(n69), .ZN(n73) );
  OAI22_X1 U101 ( .A1(n149), .A2(n30), .B1(n117), .B2(n31), .ZN(n150) );
  OAI22_X1 U102 ( .A1(n148), .A2(n30), .B1(n116), .B2(n31), .ZN(n151) );
  OAI22_X1 U103 ( .A1(n147), .A2(n30), .B1(n115), .B2(n31), .ZN(n152) );
  OAI22_X1 U104 ( .A1(n139), .A2(n30), .B1(n107), .B2(n31), .ZN(n160) );
  OAI22_X1 U105 ( .A1(n138), .A2(n30), .B1(n106), .B2(n31), .ZN(n161) );
  OAI22_X1 U106 ( .A1(n137), .A2(n30), .B1(n105), .B2(n31), .ZN(n162) );
  OAI22_X1 U107 ( .A1(n136), .A2(n30), .B1(n104), .B2(n31), .ZN(n163) );
  OAI22_X1 U108 ( .A1(n135), .A2(n30), .B1(n103), .B2(n31), .ZN(n164) );
  OAI22_X1 U109 ( .A1(n134), .A2(n30), .B1(n72), .B2(n31), .ZN(n165) );
  AND4_X1 U110 ( .A1(sel[3]), .A2(sel[2]), .A3(sel[1]), .A4(sel[0]), .ZN(n74)
         );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_15_DW_mult_tc_1 ( a, b, 
        product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n7, n9, n12, n13, n16, n18, n19, n21, n23, n25, n27, n29, n31,
         n32, n34, n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n50,
         n51, n53, n54, n55, n56, n57, n58, n59, n62, n63, n64, n65, n67, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n93, n95, n96, n97, n98, n99,
         n103, n104, n105, n106, n107, n109, n111, n112, n113, n114, n115,
         n117, n119, n120, n122, n125, n127, n131, n133, n135, n139, n141,
         n142, n143, n144, n145, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n237, n247, n249, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n418, n419, n420, n421, n422, n423, n424, n426, n427,
         n428, n429, n433, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U148 ( .A(n265), .B(n144), .Z(n145) );
  XOR2_X1 U152 ( .A(n301), .B(n148), .Z(n149) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n263), .CI(n291), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n317), .B(n252), .CO(n173), .S(n174) );
  FA_X1 U167 ( .A(n180), .B(n187), .CI(n178), .CO(n175), .S(n176) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U169 ( .A(n193), .B(n282), .CI(n191), .CO(n179), .S(n180) );
  FA_X1 U170 ( .A(n268), .B(n292), .CI(n274), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U172 ( .A(n197), .B(n190), .CI(n188), .CO(n185), .S(n186) );
  FA_X1 U173 ( .A(n199), .B(n201), .CI(n192), .CO(n187), .S(n188) );
  FA_X1 U174 ( .A(n275), .B(n293), .CI(n194), .CO(n189), .S(n190) );
  FA_X1 U175 ( .A(n253), .B(n305), .CI(n283), .CO(n191), .S(n192) );
  HA_X1 U176 ( .A(n269), .B(n319), .CO(n193), .S(n194) );
  FA_X1 U177 ( .A(n205), .B(n200), .CI(n198), .CO(n195), .S(n196) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U179 ( .A(n294), .B(n284), .CI(n276), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n320), .B(n270), .CI(n306), .CO(n201), .S(n202) );
  FA_X1 U181 ( .A(n208), .B(n213), .CI(n206), .CO(n203), .S(n204) );
  FA_X1 U182 ( .A(n215), .B(n307), .CI(n210), .CO(n205), .S(n206) );
  FA_X1 U183 ( .A(n295), .B(n285), .CI(n254), .CO(n207), .S(n208) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U185 ( .A(n216), .B(n219), .CI(n214), .CO(n211), .S(n212) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n308), .B(n278), .CI(n322), .CO(n215), .S(n216) );
  FA_X1 U188 ( .A(n225), .B(n222), .CI(n220), .CO(n217), .S(n218) );
  FA_X1 U189 ( .A(n255), .B(n309), .CI(n297), .CO(n219), .S(n220) );
  HA_X1 U190 ( .A(n323), .B(n287), .CO(n221), .S(n222) );
  FA_X1 U191 ( .A(n229), .B(n298), .CI(n226), .CO(n223), .S(n224) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  HA_X1 U194 ( .A(n311), .B(n325), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n326), .B(n300), .CI(n312), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  OR2_X1 U414 ( .A1(n224), .A2(n227), .ZN(n490) );
  OR2_X1 U415 ( .A1(n224), .A2(n227), .ZN(n491) );
  AND2_X1 U416 ( .A1(n224), .A2(n227), .ZN(n492) );
  XNOR2_X1 U417 ( .A(n554), .B(n493), .ZN(product[9]) );
  AND2_X1 U418 ( .A1(n524), .A2(n90), .ZN(n493) );
  BUF_X1 U419 ( .A(n546), .Z(n554) );
  OR2_X1 U420 ( .A1(n196), .A2(n203), .ZN(n494) );
  BUF_X1 U421 ( .A(n37), .Z(n505) );
  NOR2_X1 U422 ( .A1(n164), .A2(n175), .ZN(n75) );
  OR2_X1 U423 ( .A1(n329), .A2(n258), .ZN(n495) );
  XNOR2_X1 U424 ( .A(n564), .B(n496), .ZN(product[12]) );
  AND2_X1 U425 ( .A1(n503), .A2(n79), .ZN(n496) );
  OR2_X1 U426 ( .A1(n526), .A2(n513), .ZN(n523) );
  OR2_X1 U427 ( .A1(n526), .A2(n513), .ZN(n18) );
  XNOR2_X1 U428 ( .A(n553), .B(a[8]), .ZN(n429) );
  INV_X1 U429 ( .A(n133), .ZN(n497) );
  CLKBUF_X1 U430 ( .A(n402), .Z(n507) );
  INV_X1 U431 ( .A(n589), .ZN(n498) );
  INV_X1 U432 ( .A(n561), .ZN(n499) );
  BUF_X1 U433 ( .A(n9), .Z(n576) );
  BUF_X1 U434 ( .A(n9), .Z(n518) );
  NOR2_X1 U435 ( .A1(n228), .A2(n231), .ZN(n105) );
  INV_X1 U436 ( .A(n494), .ZN(n500) );
  OAI21_X1 U437 ( .B1(n82), .B2(n86), .A(n83), .ZN(n501) );
  XOR2_X1 U438 ( .A(n590), .B(a[6]), .Z(n538) );
  NAND2_X2 U439 ( .A1(n433), .A2(n580), .ZN(n562) );
  INV_X1 U440 ( .A(n593), .ZN(n502) );
  INV_X1 U441 ( .A(n593), .ZN(n592) );
  OR2_X1 U442 ( .A1(n176), .A2(n185), .ZN(n503) );
  XNOR2_X1 U443 ( .A(n504), .B(n166), .ZN(n164) );
  XNOR2_X1 U444 ( .A(n177), .B(n168), .ZN(n504) );
  AOI21_X1 U445 ( .B1(n104), .B2(n569), .A(n492), .ZN(n506) );
  AOI21_X1 U446 ( .B1(n490), .B2(n104), .A(n492), .ZN(n99) );
  INV_X1 U447 ( .A(n544), .ZN(n508) );
  INV_X1 U448 ( .A(n544), .ZN(n509) );
  INV_X1 U449 ( .A(n544), .ZN(n27) );
  CLKBUF_X1 U450 ( .A(n564), .Z(n510) );
  XNOR2_X1 U451 ( .A(n588), .B(a[6]), .ZN(n511) );
  OR2_X2 U452 ( .A1(n538), .A2(n511), .ZN(n512) );
  OR2_X1 U453 ( .A1(n538), .A2(n511), .ZN(n23) );
  XNOR2_X1 U454 ( .A(n585), .B(a[4]), .ZN(n513) );
  INV_X2 U455 ( .A(n513), .ZN(n16) );
  XOR2_X1 U456 ( .A(n502), .B(a[10]), .Z(n514) );
  XNOR2_X1 U457 ( .A(n271), .B(n515), .ZN(n147) );
  XNOR2_X1 U458 ( .A(n289), .B(n279), .ZN(n515) );
  OAI22_X1 U459 ( .A1(n562), .A2(n403), .B1(n507), .B2(n542), .ZN(n516) );
  BUF_X2 U460 ( .A(n9), .Z(n517) );
  XOR2_X1 U461 ( .A(n588), .B(a[4]), .Z(n526) );
  INV_X1 U462 ( .A(n508), .ZN(n519) );
  NAND2_X1 U463 ( .A1(n566), .A2(n527), .ZN(n520) );
  NAND2_X1 U464 ( .A1(n566), .A2(n527), .ZN(n521) );
  NAND2_X1 U465 ( .A1(n566), .A2(n527), .ZN(n12) );
  INV_X1 U466 ( .A(n540), .ZN(n522) );
  OR2_X1 U467 ( .A1(n204), .A2(n211), .ZN(n524) );
  INV_X1 U468 ( .A(n586), .ZN(n525) );
  INV_X1 U469 ( .A(n540), .ZN(n32) );
  XOR2_X1 U470 ( .A(n583), .B(a[2]), .Z(n527) );
  INV_X1 U471 ( .A(n548), .ZN(n528) );
  INV_X1 U472 ( .A(n590), .ZN(n529) );
  INV_X1 U473 ( .A(n590), .ZN(n589) );
  XOR2_X1 U474 ( .A(n170), .B(n172), .Z(n530) );
  XOR2_X1 U475 ( .A(n530), .B(n179), .Z(n166) );
  NAND2_X1 U476 ( .A1(n170), .A2(n172), .ZN(n531) );
  NAND2_X1 U477 ( .A1(n170), .A2(n179), .ZN(n532) );
  NAND2_X1 U478 ( .A1(n172), .A2(n179), .ZN(n533) );
  NAND3_X1 U479 ( .A1(n531), .A2(n532), .A3(n533), .ZN(n165) );
  NAND2_X1 U480 ( .A1(n177), .A2(n168), .ZN(n534) );
  NAND2_X1 U481 ( .A1(n177), .A2(n166), .ZN(n535) );
  NAND2_X1 U482 ( .A1(n168), .A2(n166), .ZN(n536) );
  NAND3_X1 U483 ( .A1(n534), .A2(n535), .A3(n536), .ZN(n163) );
  OAI21_X1 U484 ( .B1(n99), .B2(n97), .A(n98), .ZN(n537) );
  INV_X2 U485 ( .A(n588), .ZN(n586) );
  XNOR2_X1 U486 ( .A(n585), .B(a[2]), .ZN(n566) );
  XNOR2_X1 U487 ( .A(n539), .B(n310), .ZN(n226) );
  XNOR2_X1 U488 ( .A(n324), .B(n288), .ZN(n539) );
  XNOR2_X1 U489 ( .A(n591), .B(a[10]), .ZN(n540) );
  INV_X1 U490 ( .A(n249), .ZN(n580) );
  INV_X1 U491 ( .A(n580), .ZN(n541) );
  INV_X1 U492 ( .A(n541), .ZN(n542) );
  INV_X1 U493 ( .A(n541), .ZN(n543) );
  XOR2_X1 U494 ( .A(n583), .B(a[2]), .Z(n9) );
  XNOR2_X1 U495 ( .A(n590), .B(a[8]), .ZN(n544) );
  CLKBUF_X1 U496 ( .A(n74), .Z(n545) );
  AOI21_X1 U497 ( .B1(n96), .B2(n568), .A(n93), .ZN(n546) );
  INV_X1 U498 ( .A(n585), .ZN(n547) );
  INV_X1 U499 ( .A(n585), .ZN(n548) );
  AOI21_X1 U500 ( .B1(n537), .B2(n568), .A(n93), .ZN(n91) );
  CLKBUF_X1 U501 ( .A(n521), .Z(n549) );
  NAND2_X1 U502 ( .A1(n514), .A2(n32), .ZN(n550) );
  INV_X1 U503 ( .A(n591), .ZN(n551) );
  INV_X1 U504 ( .A(n591), .ZN(n552) );
  XNOR2_X1 U505 ( .A(n88), .B(n51), .ZN(product[10]) );
  BUF_X1 U506 ( .A(n591), .Z(n553) );
  CLKBUF_X1 U507 ( .A(n506), .Z(n555) );
  OAI21_X1 U508 ( .B1(n91), .B2(n89), .A(n90), .ZN(n556) );
  AOI21_X1 U509 ( .B1(n571), .B2(n112), .A(n109), .ZN(n557) );
  NAND2_X2 U510 ( .A1(n429), .A2(n27), .ZN(n29) );
  INV_X2 U511 ( .A(n565), .ZN(n21) );
  NOR2_X2 U512 ( .A1(n186), .A2(n195), .ZN(n82) );
  NAND2_X1 U513 ( .A1(n310), .A2(n516), .ZN(n558) );
  NAND2_X1 U514 ( .A1(n310), .A2(n288), .ZN(n559) );
  NAND2_X1 U515 ( .A1(n516), .A2(n288), .ZN(n560) );
  NAND3_X1 U516 ( .A1(n558), .A2(n559), .A3(n560), .ZN(n225) );
  INV_X1 U517 ( .A(n582), .ZN(n561) );
  XNOR2_X1 U518 ( .A(n583), .B(n249), .ZN(n433) );
  NAND2_X1 U519 ( .A1(n433), .A2(n580), .ZN(n563) );
  AOI21_X1 U520 ( .B1(n556), .B2(n80), .A(n501), .ZN(n564) );
  XNOR2_X1 U521 ( .A(n588), .B(a[6]), .ZN(n565) );
  NAND2_X1 U522 ( .A1(n567), .A2(n69), .ZN(n47) );
  INV_X1 U523 ( .A(n73), .ZN(n71) );
  AOI21_X1 U524 ( .B1(n545), .B2(n567), .A(n67), .ZN(n65) );
  INV_X1 U525 ( .A(n69), .ZN(n67) );
  INV_X1 U526 ( .A(n74), .ZN(n72) );
  INV_X1 U527 ( .A(n95), .ZN(n93) );
  AOI21_X1 U528 ( .B1(n556), .B2(n80), .A(n81), .ZN(n45) );
  NOR2_X1 U529 ( .A1(n82), .A2(n85), .ZN(n80) );
  OAI21_X1 U530 ( .B1(n82), .B2(n86), .A(n83), .ZN(n81) );
  NAND2_X1 U531 ( .A1(n125), .A2(n76), .ZN(n48) );
  INV_X1 U532 ( .A(n75), .ZN(n125) );
  NAND2_X1 U533 ( .A1(n494), .A2(n86), .ZN(n51) );
  OR2_X1 U534 ( .A1(n152), .A2(n163), .ZN(n567) );
  OAI21_X1 U535 ( .B1(n546), .B2(n89), .A(n90), .ZN(n88) );
  NAND2_X1 U536 ( .A1(n568), .A2(n95), .ZN(n53) );
  OAI21_X1 U537 ( .B1(n75), .B2(n79), .A(n76), .ZN(n74) );
  NAND2_X1 U538 ( .A1(n127), .A2(n83), .ZN(n50) );
  INV_X1 U539 ( .A(n82), .ZN(n127) );
  NOR2_X1 U540 ( .A1(n75), .A2(n78), .ZN(n73) );
  NAND2_X1 U541 ( .A1(n152), .A2(n163), .ZN(n69) );
  OAI21_X1 U542 ( .B1(n113), .B2(n115), .A(n114), .ZN(n112) );
  AOI21_X1 U543 ( .B1(n571), .B2(n112), .A(n109), .ZN(n107) );
  INV_X1 U544 ( .A(n111), .ZN(n109) );
  NAND2_X1 U545 ( .A1(n133), .A2(n106), .ZN(n56) );
  INV_X1 U546 ( .A(n105), .ZN(n133) );
  NAND2_X1 U547 ( .A1(n131), .A2(n98), .ZN(n54) );
  INV_X1 U548 ( .A(n97), .ZN(n131) );
  NOR2_X1 U549 ( .A1(n176), .A2(n185), .ZN(n78) );
  NOR2_X1 U550 ( .A1(n196), .A2(n203), .ZN(n85) );
  XNOR2_X1 U551 ( .A(n594), .B(n578), .ZN(n336) );
  AOI21_X1 U552 ( .B1(n570), .B2(n120), .A(n117), .ZN(n115) );
  INV_X1 U553 ( .A(n119), .ZN(n117) );
  INV_X1 U554 ( .A(n122), .ZN(n120) );
  XNOR2_X1 U555 ( .A(n63), .B(n46), .ZN(product[15]) );
  NAND2_X1 U556 ( .A1(n572), .A2(n62), .ZN(n46) );
  NAND2_X1 U557 ( .A1(n73), .A2(n567), .ZN(n64) );
  XNOR2_X1 U558 ( .A(n57), .B(n112), .ZN(product[4]) );
  NAND2_X1 U559 ( .A1(n571), .A2(n111), .ZN(n57) );
  XNOR2_X1 U560 ( .A(n59), .B(n120), .ZN(product[2]) );
  NAND2_X1 U561 ( .A1(n570), .A2(n119), .ZN(n59) );
  NAND2_X1 U562 ( .A1(n176), .A2(n185), .ZN(n79) );
  NAND2_X1 U563 ( .A1(n196), .A2(n203), .ZN(n86) );
  NAND2_X1 U564 ( .A1(n164), .A2(n175), .ZN(n76) );
  NAND2_X1 U565 ( .A1(n186), .A2(n195), .ZN(n83) );
  NAND2_X1 U566 ( .A1(n212), .A2(n217), .ZN(n95) );
  NAND2_X1 U567 ( .A1(n204), .A2(n211), .ZN(n90) );
  OR2_X1 U568 ( .A1(n212), .A2(n217), .ZN(n568) );
  AND2_X1 U569 ( .A1(n579), .A2(n247), .ZN(n314) );
  OR2_X1 U570 ( .A1(n578), .A2(n528), .ZN(n392) );
  BUF_X1 U571 ( .A(n43), .Z(n578) );
  OAI22_X1 U572 ( .A1(n42), .A2(n597), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U573 ( .A1(n578), .A2(n597), .ZN(n332) );
  OR2_X1 U574 ( .A1(n224), .A2(n227), .ZN(n569) );
  OR2_X1 U575 ( .A1(n328), .A2(n314), .ZN(n570) );
  CLKBUF_X1 U576 ( .A(n43), .Z(n579) );
  NOR2_X1 U577 ( .A1(n218), .A2(n223), .ZN(n97) );
  NAND2_X1 U578 ( .A1(n228), .A2(n231), .ZN(n106) );
  OR2_X1 U579 ( .A1(n232), .A2(n233), .ZN(n571) );
  NAND2_X1 U580 ( .A1(n218), .A2(n223), .ZN(n98) );
  INV_X1 U581 ( .A(n37), .ZN(n237) );
  INV_X1 U582 ( .A(n41), .ZN(n235) );
  OR2_X1 U583 ( .A1(n151), .A2(n139), .ZN(n572) );
  OR2_X1 U584 ( .A1(n578), .A2(n593), .ZN(n344) );
  OR2_X1 U585 ( .A1(n578), .A2(n498), .ZN(n364) );
  OR2_X1 U586 ( .A1(n578), .A2(n553), .ZN(n353) );
  OR2_X1 U587 ( .A1(n578), .A2(n525), .ZN(n377) );
  AND2_X1 U588 ( .A1(n495), .A2(n122), .ZN(product[1]) );
  XNOR2_X1 U589 ( .A(n592), .B(a[12]), .ZN(n37) );
  XNOR2_X1 U590 ( .A(n594), .B(a[14]), .ZN(n41) );
  XNOR2_X1 U591 ( .A(n552), .B(n578), .ZN(n352) );
  OAI22_X1 U592 ( .A1(n39), .A2(n336), .B1(n505), .B2(n335), .ZN(n263) );
  XNOR2_X1 U593 ( .A(n587), .B(n578), .ZN(n376) );
  XOR2_X1 U594 ( .A(n592), .B(a[10]), .Z(n428) );
  XNOR2_X1 U595 ( .A(n31), .B(n578), .ZN(n343) );
  AND2_X1 U596 ( .A1(n579), .A2(n513), .ZN(n300) );
  XOR2_X1 U597 ( .A(n315), .B(n261), .Z(n150) );
  XNOR2_X1 U598 ( .A(n155), .B(n574), .ZN(n139) );
  XNOR2_X1 U599 ( .A(n153), .B(n141), .ZN(n574) );
  XNOR2_X1 U600 ( .A(n157), .B(n575), .ZN(n141) );
  XNOR2_X1 U601 ( .A(n145), .B(n143), .ZN(n575) );
  NAND2_X1 U602 ( .A1(n427), .A2(n37), .ZN(n39) );
  XOR2_X1 U603 ( .A(n594), .B(a[12]), .Z(n427) );
  AND2_X1 U604 ( .A1(n579), .A2(n237), .ZN(n264) );
  AND2_X1 U605 ( .A1(n579), .A2(n235), .ZN(n260) );
  OAI22_X1 U606 ( .A1(n39), .A2(n335), .B1(n505), .B2(n334), .ZN(n262) );
  AND2_X1 U607 ( .A1(n579), .A2(n511), .ZN(n288) );
  AND2_X1 U608 ( .A1(n579), .A2(n540), .ZN(n270) );
  INV_X1 U609 ( .A(n19), .ZN(n590) );
  INV_X1 U610 ( .A(n25), .ZN(n591) );
  AND2_X1 U611 ( .A1(n579), .A2(n519), .ZN(n278) );
  NAND2_X1 U612 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U613 ( .A(n596), .B(a[14]), .Z(n426) );
  INV_X1 U614 ( .A(n7), .ZN(n585) );
  XNOR2_X1 U615 ( .A(n589), .B(n578), .ZN(n363) );
  OAI22_X1 U616 ( .A1(n39), .A2(n595), .B1(n337), .B2(n505), .ZN(n252) );
  OR2_X1 U617 ( .A1(n578), .A2(n595), .ZN(n337) );
  AND2_X1 U618 ( .A1(n579), .A2(n249), .ZN(product[0]) );
  XNOR2_X1 U619 ( .A(n529), .B(b[9]), .ZN(n354) );
  OAI22_X1 U620 ( .A1(n39), .A2(n334), .B1(n505), .B2(n333), .ZN(n261) );
  XNOR2_X1 U621 ( .A(n594), .B(n422), .ZN(n333) );
  XNOR2_X1 U622 ( .A(n587), .B(b[11]), .ZN(n365) );
  XNOR2_X1 U623 ( .A(n594), .B(n424), .ZN(n335) );
  XNOR2_X1 U624 ( .A(n594), .B(n423), .ZN(n334) );
  OAI22_X1 U625 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U626 ( .A(n596), .B(n424), .ZN(n330) );
  XNOR2_X1 U627 ( .A(n596), .B(n578), .ZN(n331) );
  XNOR2_X1 U628 ( .A(n551), .B(n418), .ZN(n345) );
  XNOR2_X1 U629 ( .A(n502), .B(n420), .ZN(n338) );
  XNOR2_X1 U630 ( .A(n584), .B(b[13]), .ZN(n378) );
  XNOR2_X1 U631 ( .A(n551), .B(n424), .ZN(n351) );
  XNOR2_X1 U632 ( .A(n589), .B(n424), .ZN(n362) );
  XNOR2_X1 U633 ( .A(n31), .B(n424), .ZN(n342) );
  XNOR2_X1 U634 ( .A(n502), .B(n423), .ZN(n341) );
  XNOR2_X1 U635 ( .A(n502), .B(n422), .ZN(n340) );
  XNOR2_X1 U636 ( .A(n31), .B(n421), .ZN(n339) );
  XNOR2_X1 U637 ( .A(n584), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U638 ( .A(n548), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U639 ( .A(n547), .B(n418), .ZN(n384) );
  XNOR2_X1 U640 ( .A(n547), .B(n419), .ZN(n385) );
  XNOR2_X1 U641 ( .A(n548), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U642 ( .A(n547), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U643 ( .A(n584), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U644 ( .A(n529), .B(n422), .ZN(n360) );
  XNOR2_X1 U645 ( .A(n552), .B(n422), .ZN(n349) );
  XNOR2_X1 U646 ( .A(n587), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U647 ( .A(n587), .B(n418), .ZN(n369) );
  XNOR2_X1 U648 ( .A(n587), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U649 ( .A(n587), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U650 ( .A(n529), .B(n423), .ZN(n361) );
  XNOR2_X1 U651 ( .A(n552), .B(n423), .ZN(n350) );
  XNOR2_X1 U652 ( .A(n581), .B(b[11]), .ZN(n397) );
  XNOR2_X1 U653 ( .A(n581), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U654 ( .A(n581), .B(b[13]), .ZN(n395) );
  XNOR2_X1 U655 ( .A(n581), .B(b[14]), .ZN(n394) );
  XNOR2_X1 U656 ( .A(n589), .B(n421), .ZN(n359) );
  XNOR2_X1 U657 ( .A(n589), .B(n420), .ZN(n358) );
  XNOR2_X1 U658 ( .A(n551), .B(n421), .ZN(n348) );
  XNOR2_X1 U659 ( .A(n551), .B(n420), .ZN(n347) );
  XNOR2_X1 U660 ( .A(n529), .B(n418), .ZN(n356) );
  XNOR2_X1 U661 ( .A(n529), .B(n419), .ZN(n357) );
  XNOR2_X1 U662 ( .A(n552), .B(n419), .ZN(n346) );
  XNOR2_X1 U663 ( .A(n529), .B(b[8]), .ZN(n355) );
  XNOR2_X1 U664 ( .A(n499), .B(b[15]), .ZN(n393) );
  OAI22_X1 U665 ( .A1(n550), .A2(n339), .B1(n338), .B2(n522), .ZN(n265) );
  OAI22_X1 U666 ( .A1(n550), .A2(n340), .B1(n339), .B2(n522), .ZN(n266) );
  OAI22_X1 U667 ( .A1(n550), .A2(n341), .B1(n340), .B2(n522), .ZN(n267) );
  OAI22_X1 U668 ( .A1(n34), .A2(n342), .B1(n341), .B2(n522), .ZN(n268) );
  OAI22_X1 U669 ( .A1(n550), .A2(n343), .B1(n342), .B2(n522), .ZN(n269) );
  OAI22_X1 U670 ( .A1(n34), .A2(n593), .B1(n344), .B2(n522), .ZN(n253) );
  NAND2_X1 U671 ( .A1(n428), .A2(n32), .ZN(n34) );
  INV_X1 U672 ( .A(n13), .ZN(n588) );
  OAI21_X1 U673 ( .B1(n497), .B2(n557), .A(n106), .ZN(n577) );
  NAND2_X1 U674 ( .A1(n491), .A2(n103), .ZN(n55) );
  NAND2_X1 U675 ( .A1(n224), .A2(n227), .ZN(n103) );
  NAND2_X1 U676 ( .A1(n135), .A2(n114), .ZN(n58) );
  INV_X1 U677 ( .A(n113), .ZN(n135) );
  NOR2_X1 U678 ( .A1(n204), .A2(n211), .ZN(n89) );
  OAI22_X1 U679 ( .A1(n29), .A2(n350), .B1(n349), .B2(n508), .ZN(n275) );
  OAI22_X1 U680 ( .A1(n29), .A2(n346), .B1(n345), .B2(n508), .ZN(n271) );
  OAI22_X1 U681 ( .A1(n29), .A2(n347), .B1(n346), .B2(n509), .ZN(n272) );
  OAI22_X1 U682 ( .A1(n29), .A2(n348), .B1(n347), .B2(n508), .ZN(n273) );
  OAI22_X1 U683 ( .A1(n29), .A2(n349), .B1(n348), .B2(n509), .ZN(n274) );
  OAI22_X1 U684 ( .A1(n29), .A2(n351), .B1(n350), .B2(n509), .ZN(n276) );
  OAI22_X1 U685 ( .A1(n29), .A2(n553), .B1(n353), .B2(n509), .ZN(n254) );
  OAI22_X1 U686 ( .A1(n29), .A2(n352), .B1(n351), .B2(n508), .ZN(n277) );
  XNOR2_X1 U687 ( .A(n77), .B(n48), .ZN(product[13]) );
  INV_X1 U688 ( .A(n1), .ZN(n583) );
  INV_X1 U689 ( .A(n583), .ZN(n582) );
  OR2_X1 U690 ( .A1(n578), .A2(n561), .ZN(n409) );
  INV_X2 U691 ( .A(n583), .ZN(n581) );
  XNOR2_X1 U692 ( .A(n84), .B(n50), .ZN(product[11]) );
  NAND2_X1 U693 ( .A1(n232), .A2(n233), .ZN(n111) );
  XNOR2_X1 U694 ( .A(n70), .B(n47), .ZN(product[14]) );
  OAI22_X1 U695 ( .A1(n512), .A2(n358), .B1(n357), .B2(n21), .ZN(n282) );
  OAI22_X1 U696 ( .A1(n512), .A2(n356), .B1(n355), .B2(n21), .ZN(n280) );
  OAI22_X1 U697 ( .A1(n512), .A2(n355), .B1(n354), .B2(n21), .ZN(n279) );
  OAI22_X1 U698 ( .A1(n512), .A2(n362), .B1(n361), .B2(n21), .ZN(n286) );
  OAI22_X1 U699 ( .A1(n512), .A2(n360), .B1(n359), .B2(n21), .ZN(n284) );
  OAI22_X1 U700 ( .A1(n512), .A2(n357), .B1(n356), .B2(n21), .ZN(n281) );
  OAI22_X1 U701 ( .A1(n512), .A2(n498), .B1(n364), .B2(n21), .ZN(n255) );
  OAI22_X1 U702 ( .A1(n512), .A2(n361), .B1(n360), .B2(n21), .ZN(n285) );
  XNOR2_X1 U703 ( .A(n586), .B(n424), .ZN(n375) );
  OAI22_X1 U704 ( .A1(n23), .A2(n363), .B1(n362), .B2(n21), .ZN(n287) );
  OAI22_X1 U705 ( .A1(n359), .A2(n23), .B1(n358), .B2(n21), .ZN(n283) );
  XNOR2_X1 U706 ( .A(n586), .B(n421), .ZN(n372) );
  XNOR2_X1 U707 ( .A(n586), .B(n423), .ZN(n374) );
  XNOR2_X1 U708 ( .A(n586), .B(n422), .ZN(n373) );
  XNOR2_X1 U709 ( .A(n586), .B(n419), .ZN(n370) );
  XNOR2_X1 U710 ( .A(n586), .B(n420), .ZN(n371) );
  OAI21_X1 U711 ( .B1(n506), .B2(n97), .A(n98), .ZN(n96) );
  XNOR2_X1 U712 ( .A(n581), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U713 ( .A(n582), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U714 ( .A(n582), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U715 ( .A(n581), .B(n418), .ZN(n401) );
  XNOR2_X1 U716 ( .A(n581), .B(n423), .ZN(n406) );
  XNOR2_X1 U717 ( .A(n581), .B(n422), .ZN(n405) );
  XNOR2_X1 U718 ( .A(n581), .B(n578), .ZN(n408) );
  XNOR2_X1 U719 ( .A(n581), .B(n421), .ZN(n404) );
  XNOR2_X1 U720 ( .A(n582), .B(n420), .ZN(n403) );
  XNOR2_X1 U721 ( .A(n582), .B(n419), .ZN(n402) );
  XNOR2_X1 U722 ( .A(n581), .B(n424), .ZN(n407) );
  XNOR2_X1 U723 ( .A(n55), .B(n577), .ZN(product[6]) );
  INV_X1 U724 ( .A(n88), .ZN(n87) );
  OAI21_X1 U725 ( .B1(n87), .B2(n500), .A(n86), .ZN(n84) );
  OAI21_X1 U726 ( .B1(n105), .B2(n107), .A(n106), .ZN(n104) );
  NAND2_X1 U727 ( .A1(n151), .A2(n139), .ZN(n62) );
  OAI22_X1 U728 ( .A1(n18), .A2(n370), .B1(n369), .B2(n16), .ZN(n293) );
  OAI22_X1 U729 ( .A1(n523), .A2(n367), .B1(n366), .B2(n16), .ZN(n290) );
  OAI22_X1 U730 ( .A1(n523), .A2(n375), .B1(n374), .B2(n16), .ZN(n298) );
  OAI22_X1 U731 ( .A1(n523), .A2(n368), .B1(n367), .B2(n16), .ZN(n291) );
  OAI22_X1 U732 ( .A1(n523), .A2(n373), .B1(n372), .B2(n16), .ZN(n296) );
  OAI22_X1 U733 ( .A1(n523), .A2(n369), .B1(n368), .B2(n16), .ZN(n292) );
  OAI22_X1 U734 ( .A1(n523), .A2(n372), .B1(n371), .B2(n16), .ZN(n295) );
  OAI22_X1 U735 ( .A1(n18), .A2(n371), .B1(n370), .B2(n16), .ZN(n294) );
  OAI22_X1 U736 ( .A1(n18), .A2(n374), .B1(n373), .B2(n16), .ZN(n297) );
  OAI22_X1 U737 ( .A1(n523), .A2(n376), .B1(n375), .B2(n16), .ZN(n299) );
  OAI22_X1 U738 ( .A1(n18), .A2(n525), .B1(n377), .B2(n16), .ZN(n256) );
  OAI22_X1 U739 ( .A1(n18), .A2(n366), .B1(n365), .B2(n16), .ZN(n289) );
  XNOR2_X1 U740 ( .A(n584), .B(n420), .ZN(n386) );
  XNOR2_X1 U741 ( .A(n548), .B(n578), .ZN(n391) );
  XNOR2_X1 U742 ( .A(n547), .B(n422), .ZN(n388) );
  XNOR2_X1 U743 ( .A(n548), .B(n421), .ZN(n387) );
  XNOR2_X1 U744 ( .A(n584), .B(n424), .ZN(n390) );
  XNOR2_X1 U745 ( .A(n547), .B(n423), .ZN(n389) );
  XOR2_X1 U746 ( .A(n56), .B(n557), .Z(product[5]) );
  NAND2_X1 U747 ( .A1(n328), .A2(n314), .ZN(n119) );
  NOR2_X1 U748 ( .A1(n234), .A2(n257), .ZN(n113) );
  OAI21_X1 U749 ( .B1(n64), .B2(n510), .A(n65), .ZN(n63) );
  OAI21_X1 U750 ( .B1(n71), .B2(n45), .A(n72), .ZN(n70) );
  OAI21_X1 U751 ( .B1(n45), .B2(n78), .A(n79), .ZN(n77) );
  XNOR2_X1 U752 ( .A(n537), .B(n53), .ZN(product[8]) );
  XOR2_X1 U753 ( .A(n58), .B(n115), .Z(product[3]) );
  OAI22_X1 U754 ( .A1(n562), .A2(n395), .B1(n394), .B2(n543), .ZN(n316) );
  OAI22_X1 U755 ( .A1(n562), .A2(n394), .B1(n393), .B2(n542), .ZN(n315) );
  OAI22_X1 U756 ( .A1(n562), .A2(n396), .B1(n395), .B2(n543), .ZN(n317) );
  OAI22_X1 U757 ( .A1(n562), .A2(n397), .B1(n396), .B2(n543), .ZN(n318) );
  OAI22_X1 U758 ( .A1(n562), .A2(n398), .B1(n397), .B2(n542), .ZN(n319) );
  OAI22_X1 U759 ( .A1(n562), .A2(n400), .B1(n399), .B2(n543), .ZN(n321) );
  OAI22_X1 U760 ( .A1(n563), .A2(n399), .B1(n398), .B2(n542), .ZN(n320) );
  OAI22_X1 U761 ( .A1(n562), .A2(n401), .B1(n400), .B2(n542), .ZN(n322) );
  OAI22_X1 U762 ( .A1(n563), .A2(n402), .B1(n401), .B2(n543), .ZN(n323) );
  NAND2_X1 U763 ( .A1(n329), .A2(n258), .ZN(n122) );
  OAI22_X1 U764 ( .A1(n404), .A2(n563), .B1(n403), .B2(n543), .ZN(n325) );
  OAI22_X1 U765 ( .A1(n563), .A2(n403), .B1(n402), .B2(n542), .ZN(n324) );
  OAI22_X1 U766 ( .A1(n562), .A2(n406), .B1(n405), .B2(n542), .ZN(n327) );
  OAI22_X1 U767 ( .A1(n562), .A2(n405), .B1(n404), .B2(n543), .ZN(n326) );
  OAI22_X1 U768 ( .A1(n562), .A2(n407), .B1(n406), .B2(n542), .ZN(n328) );
  OAI22_X1 U769 ( .A1(n562), .A2(n408), .B1(n407), .B2(n543), .ZN(n329) );
  OAI22_X1 U770 ( .A1(n562), .A2(n561), .B1(n409), .B2(n542), .ZN(n258) );
  XOR2_X1 U771 ( .A(n555), .B(n54), .Z(product[7]) );
  OAI22_X1 U772 ( .A1(n549), .A2(n379), .B1(n378), .B2(n518), .ZN(n301) );
  OAI22_X1 U773 ( .A1(n549), .A2(n380), .B1(n379), .B2(n518), .ZN(n302) );
  OAI22_X1 U774 ( .A1(n549), .A2(n385), .B1(n384), .B2(n517), .ZN(n307) );
  OAI22_X1 U775 ( .A1(n520), .A2(n382), .B1(n381), .B2(n517), .ZN(n304) );
  OAI22_X1 U776 ( .A1(n520), .A2(n381), .B1(n380), .B2(n518), .ZN(n303) );
  NAND2_X1 U777 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U778 ( .A1(n12), .A2(n383), .B1(n382), .B2(n576), .ZN(n305) );
  OAI22_X1 U779 ( .A1(n520), .A2(n384), .B1(n383), .B2(n517), .ZN(n306) );
  OAI22_X1 U780 ( .A1(n521), .A2(n386), .B1(n385), .B2(n517), .ZN(n308) );
  OAI22_X1 U781 ( .A1(n521), .A2(n387), .B1(n386), .B2(n517), .ZN(n309) );
  OAI22_X1 U782 ( .A1(n521), .A2(n528), .B1(n392), .B2(n517), .ZN(n257) );
  OAI22_X1 U783 ( .A1(n12), .A2(n389), .B1(n388), .B2(n576), .ZN(n311) );
  OAI22_X1 U784 ( .A1(n520), .A2(n388), .B1(n518), .B2(n387), .ZN(n310) );
  OAI22_X1 U785 ( .A1(n521), .A2(n390), .B1(n389), .B2(n517), .ZN(n312) );
  INV_X1 U786 ( .A(n518), .ZN(n247) );
  OAI22_X1 U787 ( .A1(n521), .A2(n391), .B1(n390), .B2(n518), .ZN(n313) );
  INV_X1 U788 ( .A(n585), .ZN(n584) );
  INV_X1 U789 ( .A(n588), .ZN(n587) );
  INV_X1 U790 ( .A(n31), .ZN(n593) );
  INV_X1 U791 ( .A(n595), .ZN(n594) );
  INV_X1 U792 ( .A(n36), .ZN(n595) );
  INV_X1 U793 ( .A(n597), .ZN(n596) );
  INV_X1 U794 ( .A(n40), .ZN(n597) );
  XOR2_X1 U795 ( .A(n259), .B(n251), .Z(n148) );
  XOR2_X1 U796 ( .A(n149), .B(n147), .Z(n144) );
  XOR2_X1 U797 ( .A(n159), .B(n150), .Z(n142) );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_15_DW01_add_2 ( A, B, CI, 
        SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n19,
         n20, n22, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n44, n45, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n65, n67, n68, n69, n70, n71,
         n73, n75, n76, n77, n78, n79, n81, n83, n84, n86, n89, n90, n91, n94,
         n95, n96, n98, n100, n157, n158, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176;

  NOR2_X2 U122 ( .A1(A[8]), .A2(B[8]), .ZN(n54) );
  AOI21_X1 U123 ( .B1(n38), .B2(n30), .A(n31), .ZN(n157) );
  OR2_X1 U124 ( .A1(n25), .A2(n28), .ZN(n158) );
  AND2_X1 U125 ( .A1(n170), .A2(n86), .ZN(SUM[0]) );
  OR2_X1 U126 ( .A1(A[15]), .A2(B[15]), .ZN(n160) );
  XNOR2_X1 U127 ( .A(n161), .B(n37), .ZN(SUM[11]) );
  AND2_X1 U128 ( .A1(n91), .A2(n36), .ZN(n161) );
  NOR2_X1 U129 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  AND2_X1 U130 ( .A1(A[9]), .A2(B[9]), .ZN(n162) );
  CLKBUF_X1 U131 ( .A(n176), .Z(n163) );
  OR2_X1 U132 ( .A1(A[10]), .A2(B[10]), .ZN(n164) );
  OR2_X1 U133 ( .A1(A[10]), .A2(B[10]), .ZN(n175) );
  NOR2_X1 U134 ( .A1(A[14]), .A2(B[14]), .ZN(n165) );
  NOR2_X1 U135 ( .A1(A[14]), .A2(B[14]), .ZN(n25) );
  NOR2_X1 U136 ( .A1(A[12]), .A2(B[12]), .ZN(n166) );
  NOR2_X1 U137 ( .A1(A[12]), .A2(B[12]), .ZN(n32) );
  INV_X1 U138 ( .A(n91), .ZN(n167) );
  OR2_X1 U139 ( .A1(A[14]), .A2(B[14]), .ZN(n168) );
  AOI21_X1 U140 ( .B1(n38), .B2(n30), .A(n31), .ZN(n169) );
  OR2_X1 U141 ( .A1(A[0]), .A2(B[0]), .ZN(n170) );
  INV_X1 U142 ( .A(n60), .ZN(n59) );
  INV_X1 U143 ( .A(n38), .ZN(n37) );
  OAI21_X1 U144 ( .B1(n71), .B2(n69), .A(n70), .ZN(n68) );
  AOI21_X1 U145 ( .B1(n172), .B2(n84), .A(n81), .ZN(n79) );
  INV_X1 U146 ( .A(n83), .ZN(n81) );
  OAI21_X1 U147 ( .B1(n79), .B2(n77), .A(n78), .ZN(n76) );
  AOI21_X1 U148 ( .B1(n174), .B2(n68), .A(n65), .ZN(n63) );
  INV_X1 U149 ( .A(n67), .ZN(n65) );
  INV_X1 U150 ( .A(n24), .ZN(n22) );
  AOI21_X1 U151 ( .B1(n173), .B2(n76), .A(n73), .ZN(n71) );
  INV_X1 U152 ( .A(n75), .ZN(n73) );
  AOI21_X1 U153 ( .B1(n50), .B2(n171), .A(n162), .ZN(n45) );
  INV_X1 U154 ( .A(n86), .ZN(n84) );
  OAI21_X1 U155 ( .B1(n59), .B2(n57), .A(n58), .ZN(n56) );
  INV_X1 U156 ( .A(n35), .ZN(n91) );
  INV_X1 U157 ( .A(n28), .ZN(n89) );
  NAND2_X1 U158 ( .A1(n98), .A2(n70), .ZN(n13) );
  INV_X1 U159 ( .A(n69), .ZN(n98) );
  NAND2_X1 U160 ( .A1(n173), .A2(n75), .ZN(n14) );
  NAND2_X1 U161 ( .A1(n95), .A2(n58), .ZN(n10) );
  INV_X1 U162 ( .A(n57), .ZN(n95) );
  NAND2_X1 U163 ( .A1(n171), .A2(n49), .ZN(n8) );
  NAND2_X1 U164 ( .A1(n100), .A2(n78), .ZN(n15) );
  INV_X1 U165 ( .A(n77), .ZN(n100) );
  NAND2_X1 U166 ( .A1(n94), .A2(n55), .ZN(n9) );
  INV_X1 U167 ( .A(n54), .ZN(n94) );
  NAND2_X1 U168 ( .A1(n174), .A2(n67), .ZN(n12) );
  NAND2_X1 U169 ( .A1(n172), .A2(n83), .ZN(n16) );
  NAND2_X1 U170 ( .A1(n96), .A2(n62), .ZN(n11) );
  INV_X1 U171 ( .A(n61), .ZN(n96) );
  XNOR2_X1 U172 ( .A(n12), .B(n68), .ZN(SUM[5]) );
  XNOR2_X1 U173 ( .A(n14), .B(n76), .ZN(SUM[3]) );
  XOR2_X1 U174 ( .A(n15), .B(n79), .Z(SUM[2]) );
  XNOR2_X1 U175 ( .A(n16), .B(n84), .ZN(SUM[1]) );
  NAND2_X1 U176 ( .A1(n168), .A2(n26), .ZN(n3) );
  NAND2_X1 U177 ( .A1(n90), .A2(n33), .ZN(n5) );
  NAND2_X1 U178 ( .A1(n89), .A2(n29), .ZN(n4) );
  NOR2_X1 U179 ( .A1(A[11]), .A2(B[11]), .ZN(n35) );
  NOR2_X1 U180 ( .A1(A[7]), .A2(B[7]), .ZN(n57) );
  OR2_X1 U181 ( .A1(A[9]), .A2(B[9]), .ZN(n171) );
  NOR2_X1 U182 ( .A1(A[2]), .A2(B[2]), .ZN(n77) );
  NAND2_X1 U183 ( .A1(A[13]), .A2(B[13]), .ZN(n29) );
  NAND2_X1 U184 ( .A1(A[11]), .A2(B[11]), .ZN(n36) );
  OR2_X1 U185 ( .A1(A[1]), .A2(B[1]), .ZN(n172) );
  OR2_X1 U186 ( .A1(A[3]), .A2(B[3]), .ZN(n173) );
  NOR2_X1 U187 ( .A1(A[4]), .A2(B[4]), .ZN(n69) );
  NAND2_X1 U188 ( .A1(A[14]), .A2(B[14]), .ZN(n26) );
  NAND2_X1 U189 ( .A1(A[12]), .A2(B[12]), .ZN(n33) );
  XNOR2_X1 U190 ( .A(n50), .B(n8), .ZN(SUM[9]) );
  XNOR2_X1 U191 ( .A(n56), .B(n9), .ZN(SUM[8]) );
  NOR2_X1 U192 ( .A1(A[6]), .A2(B[6]), .ZN(n61) );
  NAND2_X1 U193 ( .A1(A[7]), .A2(B[7]), .ZN(n58) );
  OR2_X1 U194 ( .A1(A[5]), .A2(B[5]), .ZN(n174) );
  NAND2_X1 U195 ( .A1(A[2]), .A2(B[2]), .ZN(n78) );
  NAND2_X1 U196 ( .A1(A[9]), .A2(B[9]), .ZN(n49) );
  NAND2_X1 U197 ( .A1(A[5]), .A2(B[5]), .ZN(n67) );
  NAND2_X1 U198 ( .A1(A[1]), .A2(B[1]), .ZN(n83) );
  NAND2_X1 U199 ( .A1(A[0]), .A2(B[0]), .ZN(n86) );
  NAND2_X1 U200 ( .A1(A[4]), .A2(B[4]), .ZN(n70) );
  NAND2_X1 U201 ( .A1(A[6]), .A2(B[6]), .ZN(n62) );
  NAND2_X1 U202 ( .A1(A[8]), .A2(B[8]), .ZN(n55) );
  XOR2_X1 U203 ( .A(n7), .B(n45), .Z(SUM[10]) );
  XOR2_X1 U204 ( .A(n59), .B(n10), .Z(SUM[7]) );
  NAND2_X1 U205 ( .A1(n160), .A2(n19), .ZN(n2) );
  XOR2_X1 U206 ( .A(n11), .B(n63), .Z(SUM[6]) );
  OAI21_X1 U207 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  NOR2_X1 U208 ( .A1(n54), .A2(n57), .ZN(n52) );
  OAI21_X1 U209 ( .B1(n54), .B2(n58), .A(n55), .ZN(n53) );
  XOR2_X1 U210 ( .A(n13), .B(n71), .Z(SUM[4]) );
  NAND2_X1 U211 ( .A1(A[3]), .A2(B[3]), .ZN(n75) );
  INV_X1 U212 ( .A(n163), .ZN(n44) );
  AND2_X1 U213 ( .A1(A[10]), .A2(B[10]), .ZN(n176) );
  INV_X1 U214 ( .A(n51), .ZN(n50) );
  OAI21_X1 U215 ( .B1(n37), .B2(n167), .A(n36), .ZN(n34) );
  AOI21_X1 U216 ( .B1(n52), .B2(n60), .A(n53), .ZN(n51) );
  AOI21_X1 U217 ( .B1(n175), .B2(n162), .A(n176), .ZN(n40) );
  INV_X1 U218 ( .A(n166), .ZN(n90) );
  NOR2_X1 U219 ( .A1(n166), .A2(n35), .ZN(n30) );
  OAI21_X1 U220 ( .B1(n32), .B2(n36), .A(n33), .ZN(n31) );
  OAI21_X1 U221 ( .B1(n165), .B2(n29), .A(n26), .ZN(n24) );
  NAND2_X1 U222 ( .A1(A[15]), .A2(B[15]), .ZN(n19) );
  OAI21_X1 U223 ( .B1(n39), .B2(n51), .A(n40), .ZN(n38) );
  NAND2_X1 U224 ( .A1(n44), .A2(n164), .ZN(n7) );
  NAND2_X1 U225 ( .A1(n164), .A2(n171), .ZN(n39) );
  XNOR2_X1 U226 ( .A(n34), .B(n5), .ZN(SUM[12]) );
  XNOR2_X1 U227 ( .A(n20), .B(n2), .ZN(SUM[15]) );
  XNOR2_X1 U228 ( .A(n27), .B(n3), .ZN(SUM[14]) );
  XOR2_X1 U229 ( .A(n169), .B(n4), .Z(SUM[13]) );
  OAI21_X1 U230 ( .B1(n157), .B2(n28), .A(n29), .ZN(n27) );
  OAI21_X1 U231 ( .B1(n158), .B2(n157), .A(n22), .ZN(n20) );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_15 ( clk, clear_acc, 
        data_out_x, data_out, data_out_w, data_out_b, wr_en_y, m_valid, 
        m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [4:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
         N39, N40, N41, N42, N43, N44, n1, n2, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n85, n102, n111, n112, n113, n114, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n17), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n221), .CK(clk), .Q(n21) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n222), .CK(clk), .Q(n22) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n223), .CK(clk), .Q(n23) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n224), .CK(clk), .Q(n24) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n225), .CK(clk), .Q(n25) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n226), .CK(clk), .Q(n26) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n227), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n228), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n229), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n230), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n231), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n232), .CK(clk), .Q(n34) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n233), .CK(clk), .Q(n35) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n234), .CK(clk), .Q(n36) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n235), .CK(clk), .Q(n37) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n236), .CK(clk), .Q(n39) );
  DFF_X1 \f_reg[0]  ( .D(n111), .CK(clk), .Q(f[0]), .QN(n210) );
  DFF_X1 \f_reg[1]  ( .D(n102), .CK(clk), .Q(f[1]), .QN(n211) );
  DFF_X1 \f_reg[2]  ( .D(n85), .CK(clk), .Q(f[2]), .QN(n212) );
  DFF_X1 \f_reg[7]  ( .D(n79), .CK(clk), .Q(f[7]), .QN(n213) );
  DFF_X1 \f_reg[8]  ( .D(n78), .CK(clk), .Q(f[8]), .QN(n214) );
  DFF_X1 \f_reg[9]  ( .D(n77), .CK(clk), .Q(f[9]), .QN(n215) );
  DFF_X1 \f_reg[10]  ( .D(n76), .CK(clk), .Q(n49), .QN(n216) );
  DFF_X1 \f_reg[11]  ( .D(n75), .CK(clk), .Q(n47), .QN(n217) );
  DFF_X1 \f_reg[12]  ( .D(n1), .CK(clk), .Q(n46), .QN(n218) );
  DFF_X1 \f_reg[13]  ( .D(n74), .CK(clk), .Q(n44), .QN(n219) );
  DFF_X1 \f_reg[14]  ( .D(n2), .CK(clk), .Q(n43), .QN(n220) );
  DFF_X1 \f_reg[15]  ( .D(n73), .CK(clk), .Q(f[15]), .QN(n70) );
  DFF_X1 \data_out_reg[15]  ( .D(n113), .CK(clk), .Q(data_out[15]), .QN(n193)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n114), .CK(clk), .Q(data_out[14]), .QN(n192)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n164), .CK(clk), .Q(data_out[13]), .QN(n191)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n165), .CK(clk), .Q(data_out[12]), .QN(n190)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n166), .CK(clk), .Q(data_out[11]), .QN(n189)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n167), .CK(clk), .Q(data_out[10]), .QN(n188)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n168), .CK(clk), .Q(data_out[9]), .QN(n187) );
  DFF_X1 \data_out_reg[8]  ( .D(n169), .CK(clk), .Q(data_out[8]), .QN(n186) );
  DFF_X1 \data_out_reg[7]  ( .D(n170), .CK(clk), .Q(data_out[7]), .QN(n185) );
  DFF_X1 \data_out_reg[6]  ( .D(n171), .CK(clk), .Q(data_out[6]), .QN(n184) );
  DFF_X1 \data_out_reg[5]  ( .D(n172), .CK(clk), .Q(data_out[5]), .QN(n183) );
  DFF_X1 \data_out_reg[4]  ( .D(n173), .CK(clk), .Q(data_out[4]), .QN(n182) );
  DFF_X1 \data_out_reg[3]  ( .D(n174), .CK(clk), .Q(data_out[3]), .QN(n181) );
  DFF_X1 \data_out_reg[2]  ( .D(n175), .CK(clk), .Q(data_out[2]), .QN(n180) );
  DFF_X1 \data_out_reg[1]  ( .D(n176), .CK(clk), .Q(data_out[1]), .QN(n179) );
  DFF_X1 \data_out_reg[0]  ( .D(n177), .CK(clk), .Q(data_out[0]), .QN(n178) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_15_DW_mult_tc_1 mult_2021 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_15_DW01_add_2 add_2022 ( .A({
        n200, n199, n198, n197, n196, n195, n209, n208, n207, n206, n205, n204, 
        n203, n202, n201, n194}), .B({f[15], n43, n44, n46, n47, n49, f[9:0]}), 
        .CI(1'b0), .SUM(adder) );
  DFF_X1 \f_reg[3]  ( .D(n83), .CK(clk), .Q(f[3]), .QN(n62) );
  DFF_X1 \f_reg[4]  ( .D(n82), .CK(clk), .Q(f[4]), .QN(n63) );
  DFF_X1 \f_reg[5]  ( .D(n81), .CK(clk), .Q(f[5]), .QN(n64) );
  DFF_X1 \f_reg[6]  ( .D(n80), .CK(clk), .Q(f[6]), .QN(n65) );
  DFF_X2 delay_reg ( .D(n112), .CK(clk), .Q(n8), .QN(n237) );
  MUX2_X1 U3 ( .A(n27), .B(N38), .S(n237), .Z(n209) );
  INV_X1 U4 ( .A(n42), .ZN(n60) );
  AND2_X1 U5 ( .A1(n42), .A2(n18), .ZN(n15) );
  NAND3_X1 U6 ( .A1(n5), .A2(n4), .A3(n6), .ZN(n1) );
  NAND3_X1 U8 ( .A1(n13), .A2(n12), .A3(n14), .ZN(n2) );
  NAND2_X1 U9 ( .A1(data_out_b[12]), .A2(n17), .ZN(n4) );
  NAND2_X1 U10 ( .A1(adder[12]), .A2(n15), .ZN(n5) );
  NAND2_X1 U11 ( .A1(n60), .A2(n46), .ZN(n6) );
  AND2_X1 U12 ( .A1(n11), .A2(n9), .ZN(n7) );
  NAND2_X1 U13 ( .A1(n10), .A2(n7), .ZN(n73) );
  MUX2_X2 U14 ( .A(n25), .B(N40), .S(n237), .Z(n196) );
  MUX2_X2 U15 ( .A(N39), .B(n26), .S(n8), .Z(n195) );
  MUX2_X2 U16 ( .A(n23), .B(N42), .S(n237), .Z(n198) );
  MUX2_X2 U17 ( .A(n22), .B(N43), .S(n237), .Z(n199) );
  MUX2_X2 U18 ( .A(n24), .B(N41), .S(n237), .Z(n197) );
  NAND2_X1 U19 ( .A1(data_out_b[15]), .A2(n17), .ZN(n9) );
  NAND2_X1 U20 ( .A1(adder[15]), .A2(n15), .ZN(n10) );
  NAND2_X1 U21 ( .A1(n60), .A2(f[15]), .ZN(n11) );
  NAND2_X1 U22 ( .A1(data_out_b[14]), .A2(n17), .ZN(n12) );
  NAND2_X1 U23 ( .A1(adder[14]), .A2(n15), .ZN(n13) );
  NAND2_X1 U24 ( .A1(n60), .A2(n43), .ZN(n14) );
  INV_X1 U25 ( .A(n18), .ZN(n17) );
  NAND2_X1 U26 ( .A1(n112), .A2(n16), .ZN(n239) );
  INV_X1 U27 ( .A(clear_acc), .ZN(n18) );
  OAI22_X1 U28 ( .A1(n181), .A2(n239), .B1(n62), .B2(n238), .ZN(n174) );
  OAI22_X1 U29 ( .A1(n182), .A2(n239), .B1(n63), .B2(n238), .ZN(n173) );
  OAI22_X1 U30 ( .A1(n183), .A2(n239), .B1(n64), .B2(n238), .ZN(n172) );
  OAI22_X1 U31 ( .A1(n184), .A2(n239), .B1(n65), .B2(n238), .ZN(n171) );
  OAI22_X1 U32 ( .A1(n185), .A2(n239), .B1(n213), .B2(n238), .ZN(n170) );
  OAI22_X1 U33 ( .A1(n186), .A2(n239), .B1(n214), .B2(n238), .ZN(n169) );
  OAI22_X1 U34 ( .A1(n187), .A2(n239), .B1(n215), .B2(n238), .ZN(n168) );
  INV_X1 U35 ( .A(n20), .ZN(n38) );
  INV_X1 U36 ( .A(wr_en_y), .ZN(n16) );
  INV_X1 U37 ( .A(m_ready), .ZN(n19) );
  NAND2_X1 U38 ( .A1(m_valid), .A2(n19), .ZN(n40) );
  OAI21_X1 U39 ( .B1(sel[4]), .B2(n72), .A(n40), .ZN(n112) );
  NAND2_X1 U40 ( .A1(clear_acc_delay), .A2(n237), .ZN(n20) );
  MUX2_X1 U41 ( .A(n21), .B(N44), .S(n38), .Z(n221) );
  MUX2_X1 U42 ( .A(n21), .B(N44), .S(n237), .Z(n200) );
  MUX2_X1 U43 ( .A(n22), .B(N43), .S(n38), .Z(n222) );
  MUX2_X1 U44 ( .A(n23), .B(N42), .S(n38), .Z(n223) );
  MUX2_X1 U45 ( .A(n24), .B(N41), .S(n38), .Z(n224) );
  MUX2_X1 U46 ( .A(n25), .B(N40), .S(n38), .Z(n225) );
  MUX2_X1 U47 ( .A(n26), .B(N39), .S(n38), .Z(n226) );
  MUX2_X1 U48 ( .A(n27), .B(N38), .S(n38), .Z(n227) );
  MUX2_X1 U49 ( .A(n28), .B(N37), .S(n38), .Z(n228) );
  MUX2_X1 U50 ( .A(n28), .B(N37), .S(n237), .Z(n208) );
  MUX2_X1 U51 ( .A(n29), .B(N36), .S(n38), .Z(n229) );
  MUX2_X1 U52 ( .A(n29), .B(N36), .S(n237), .Z(n207) );
  MUX2_X1 U53 ( .A(n32), .B(N35), .S(n38), .Z(n230) );
  MUX2_X1 U54 ( .A(n32), .B(N35), .S(n237), .Z(n206) );
  MUX2_X1 U55 ( .A(n33), .B(N34), .S(n38), .Z(n231) );
  MUX2_X1 U56 ( .A(n33), .B(N34), .S(n237), .Z(n205) );
  MUX2_X1 U57 ( .A(n34), .B(N33), .S(n38), .Z(n232) );
  MUX2_X1 U58 ( .A(n34), .B(N33), .S(n237), .Z(n204) );
  MUX2_X1 U59 ( .A(n35), .B(N32), .S(n38), .Z(n233) );
  MUX2_X1 U60 ( .A(n35), .B(N32), .S(n237), .Z(n203) );
  MUX2_X1 U61 ( .A(n36), .B(N31), .S(n38), .Z(n234) );
  MUX2_X1 U62 ( .A(n36), .B(N31), .S(n237), .Z(n202) );
  MUX2_X1 U63 ( .A(n37), .B(N30), .S(n38), .Z(n235) );
  MUX2_X1 U64 ( .A(n37), .B(N30), .S(n237), .Z(n201) );
  MUX2_X1 U65 ( .A(n39), .B(N29), .S(n38), .Z(n236) );
  MUX2_X1 U66 ( .A(n39), .B(N29), .S(n237), .Z(n194) );
  INV_X1 U67 ( .A(n40), .ZN(n41) );
  OAI21_X1 U68 ( .B1(n41), .B2(n8), .A(n18), .ZN(n42) );
  AOI222_X1 U69 ( .A1(data_out_b[13]), .A2(n17), .B1(adder[13]), .B2(n15), 
        .C1(n60), .C2(n44), .ZN(n45) );
  INV_X1 U70 ( .A(n45), .ZN(n74) );
  AOI222_X1 U71 ( .A1(data_out_b[11]), .A2(n17), .B1(adder[11]), .B2(n15), 
        .C1(n60), .C2(n47), .ZN(n48) );
  INV_X1 U72 ( .A(n48), .ZN(n75) );
  AOI222_X1 U73 ( .A1(data_out_b[10]), .A2(n17), .B1(adder[10]), .B2(n15), 
        .C1(n60), .C2(n49), .ZN(n50) );
  INV_X1 U74 ( .A(n50), .ZN(n76) );
  AOI222_X1 U75 ( .A1(data_out_b[8]), .A2(n17), .B1(adder[8]), .B2(n15), .C1(
        n60), .C2(f[8]), .ZN(n51) );
  INV_X1 U76 ( .A(n51), .ZN(n78) );
  AOI222_X1 U77 ( .A1(data_out_b[7]), .A2(n17), .B1(adder[7]), .B2(n15), .C1(
        n60), .C2(f[7]), .ZN(n52) );
  INV_X1 U78 ( .A(n52), .ZN(n79) );
  AOI222_X1 U79 ( .A1(data_out_b[6]), .A2(n17), .B1(adder[6]), .B2(n15), .C1(
        n60), .C2(f[6]), .ZN(n53) );
  INV_X1 U80 ( .A(n53), .ZN(n80) );
  AOI222_X1 U81 ( .A1(data_out_b[5]), .A2(n17), .B1(adder[5]), .B2(n15), .C1(
        n60), .C2(f[5]), .ZN(n54) );
  INV_X1 U82 ( .A(n54), .ZN(n81) );
  AOI222_X1 U83 ( .A1(data_out_b[4]), .A2(n17), .B1(adder[4]), .B2(n15), .C1(
        n60), .C2(f[4]), .ZN(n55) );
  INV_X1 U84 ( .A(n55), .ZN(n82) );
  AOI222_X1 U85 ( .A1(data_out_b[3]), .A2(n17), .B1(adder[3]), .B2(n15), .C1(
        n60), .C2(f[3]), .ZN(n56) );
  INV_X1 U86 ( .A(n56), .ZN(n83) );
  AOI222_X1 U87 ( .A1(data_out_b[2]), .A2(n17), .B1(adder[2]), .B2(n15), .C1(
        n60), .C2(f[2]), .ZN(n57) );
  INV_X1 U88 ( .A(n57), .ZN(n85) );
  AOI222_X1 U89 ( .A1(data_out_b[1]), .A2(n17), .B1(adder[1]), .B2(n15), .C1(
        n60), .C2(f[1]), .ZN(n58) );
  INV_X1 U90 ( .A(n58), .ZN(n102) );
  AOI222_X1 U91 ( .A1(data_out_b[0]), .A2(n17), .B1(adder[0]), .B2(n15), .C1(
        n60), .C2(f[0]), .ZN(n59) );
  INV_X1 U92 ( .A(n59), .ZN(n111) );
  AOI222_X1 U93 ( .A1(data_out_b[9]), .A2(n17), .B1(adder[9]), .B2(n15), .C1(
        n60), .C2(f[9]), .ZN(n61) );
  INV_X1 U94 ( .A(n61), .ZN(n77) );
  NOR4_X1 U95 ( .A1(n47), .A2(n46), .A3(n44), .A4(n43), .ZN(n69) );
  NOR4_X1 U96 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n49), .ZN(n68) );
  NAND4_X1 U97 ( .A1(n65), .A2(n64), .A3(n63), .A4(n62), .ZN(n66) );
  NOR4_X1 U98 ( .A1(n66), .A2(f[0]), .A3(f[1]), .A4(f[2]), .ZN(n67) );
  NAND3_X1 U99 ( .A1(n69), .A2(n68), .A3(n67), .ZN(n71) );
  NAND3_X1 U100 ( .A1(wr_en_y), .A2(n71), .A3(n70), .ZN(n238) );
  OAI22_X1 U101 ( .A1(n178), .A2(n239), .B1(n210), .B2(n238), .ZN(n177) );
  OAI22_X1 U102 ( .A1(n179), .A2(n239), .B1(n211), .B2(n238), .ZN(n176) );
  OAI22_X1 U103 ( .A1(n180), .A2(n239), .B1(n212), .B2(n238), .ZN(n175) );
  OAI22_X1 U104 ( .A1(n188), .A2(n239), .B1(n216), .B2(n238), .ZN(n167) );
  OAI22_X1 U105 ( .A1(n189), .A2(n239), .B1(n217), .B2(n238), .ZN(n166) );
  OAI22_X1 U106 ( .A1(n190), .A2(n239), .B1(n218), .B2(n238), .ZN(n165) );
  OAI22_X1 U107 ( .A1(n191), .A2(n239), .B1(n219), .B2(n238), .ZN(n164) );
  OAI22_X1 U108 ( .A1(n192), .A2(n239), .B1(n220), .B2(n238), .ZN(n114) );
  OAI22_X1 U109 ( .A1(n193), .A2(n239), .B1(n70), .B2(n238), .ZN(n113) );
  AND4_X1 U110 ( .A1(sel[3]), .A2(sel[2]), .A3(sel[1]), .A4(sel[0]), .ZN(n72)
         );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_14_DW_mult_tc_1 ( a, b, 
        product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n9, n12, n13, n16, n18, n19, n23, n25, n27, n29, n31, n32,
         n34, n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n62, n63, n64, n65, n67, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n93, n95, n96, n97, n98, n99,
         n101, n103, n104, n105, n106, n107, n109, n111, n112, n113, n114,
         n115, n117, n119, n120, n122, n125, n127, n128, n131, n133, n135,
         n139, n141, n142, n143, n144, n145, n147, n148, n149, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n237, n247, n249, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n418, n419, n420, n421, n422, n423, n424, n426,
         n427, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U148 ( .A(n265), .B(n144), .Z(n145) );
  XOR2_X1 U152 ( .A(n301), .B(n148), .Z(n149) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n263), .CI(n291), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n317), .B(n252), .CO(n173), .S(n174) );
  FA_X1 U167 ( .A(n180), .B(n187), .CI(n178), .CO(n175), .S(n176) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U169 ( .A(n193), .B(n282), .CI(n191), .CO(n179), .S(n180) );
  FA_X1 U170 ( .A(n268), .B(n292), .CI(n274), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U172 ( .A(n197), .B(n190), .CI(n188), .CO(n185), .S(n186) );
  FA_X1 U173 ( .A(n199), .B(n201), .CI(n192), .CO(n187), .S(n188) );
  FA_X1 U175 ( .A(n253), .B(n305), .CI(n283), .CO(n191), .S(n192) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U179 ( .A(n294), .B(n284), .CI(n276), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n320), .B(n270), .CI(n306), .CO(n201), .S(n202) );
  FA_X1 U181 ( .A(n208), .B(n213), .CI(n206), .CO(n203), .S(n204) );
  FA_X1 U182 ( .A(n210), .B(n307), .CI(n215), .CO(n205), .S(n206) );
  FA_X1 U183 ( .A(n295), .B(n285), .CI(n254), .CO(n207), .S(n208) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U185 ( .A(n216), .B(n219), .CI(n214), .CO(n211), .S(n212) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n322), .B(n278), .CI(n308), .CO(n215), .S(n216) );
  FA_X1 U188 ( .A(n225), .B(n222), .CI(n220), .CO(n217), .S(n218) );
  FA_X1 U189 ( .A(n255), .B(n297), .CI(n309), .CO(n219), .S(n220) );
  HA_X1 U190 ( .A(n323), .B(n287), .CO(n221), .S(n222) );
  FA_X1 U192 ( .A(n310), .B(n288), .CI(n324), .CO(n225), .S(n226) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  HA_X1 U194 ( .A(n311), .B(n325), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n326), .B(n300), .CI(n312), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  BUF_X1 U414 ( .A(n96), .Z(n551) );
  BUF_X1 U415 ( .A(n73), .Z(n490) );
  NOR2_X1 U416 ( .A1(n553), .A2(n85), .ZN(n491) );
  XNOR2_X1 U417 ( .A(n13), .B(a[6]), .ZN(n493) );
  OR2_X4 U418 ( .A1(n520), .A2(n536), .ZN(n18) );
  NAND2_X2 U419 ( .A1(n492), .A2(n493), .ZN(n23) );
  XNOR2_X1 U420 ( .A(n593), .B(a[6]), .ZN(n492) );
  INV_X1 U421 ( .A(n563), .ZN(n27) );
  OR2_X1 U422 ( .A1(n329), .A2(n258), .ZN(n494) );
  BUF_X2 U423 ( .A(n9), .Z(n495) );
  CLKBUF_X1 U424 ( .A(n9), .Z(n580) );
  INV_X1 U425 ( .A(n595), .ZN(n544) );
  CLKBUF_X1 U426 ( .A(n95), .Z(n496) );
  XNOR2_X1 U427 ( .A(n271), .B(n497), .ZN(n147) );
  XNOR2_X1 U428 ( .A(n289), .B(n279), .ZN(n497) );
  XNOR2_X1 U429 ( .A(n509), .B(n498), .ZN(product[12]) );
  AND2_X1 U430 ( .A1(n547), .A2(n79), .ZN(n498) );
  XOR2_X1 U431 ( .A(n591), .B(a[6]), .Z(n499) );
  XNOR2_X1 U432 ( .A(n589), .B(a[2]), .ZN(n500) );
  CLKBUF_X1 U433 ( .A(n585), .Z(n501) );
  CLKBUF_X3 U434 ( .A(n585), .Z(n502) );
  CLKBUF_X3 U435 ( .A(n585), .Z(n503) );
  INV_X1 U436 ( .A(n586), .ZN(n585) );
  XNOR2_X1 U437 ( .A(n226), .B(n504), .ZN(n224) );
  XNOR2_X1 U438 ( .A(n229), .B(n298), .ZN(n504) );
  AOI21_X1 U439 ( .B1(n573), .B2(n120), .A(n117), .ZN(n505) );
  INV_X1 U440 ( .A(n542), .ZN(n506) );
  NAND2_X1 U441 ( .A1(n500), .A2(n539), .ZN(n507) );
  NOR2_X1 U442 ( .A1(n228), .A2(n231), .ZN(n508) );
  NOR2_X1 U443 ( .A1(n228), .A2(n231), .ZN(n105) );
  AOI21_X1 U444 ( .B1(n522), .B2(n491), .A(n81), .ZN(n509) );
  CLKBUF_X1 U445 ( .A(n565), .Z(n510) );
  XOR2_X1 U446 ( .A(n275), .B(n293), .Z(n511) );
  XOR2_X1 U447 ( .A(n194), .B(n511), .Z(n190) );
  NAND2_X1 U448 ( .A1(n194), .A2(n275), .ZN(n512) );
  NAND2_X1 U449 ( .A1(n194), .A2(n293), .ZN(n513) );
  NAND2_X1 U450 ( .A1(n275), .A2(n293), .ZN(n514) );
  NAND3_X1 U451 ( .A1(n512), .A2(n513), .A3(n514), .ZN(n189) );
  XOR2_X1 U452 ( .A(n205), .B(n200), .Z(n515) );
  XOR2_X1 U453 ( .A(n198), .B(n515), .Z(n196) );
  NAND2_X1 U454 ( .A1(n198), .A2(n205), .ZN(n516) );
  NAND2_X1 U455 ( .A1(n198), .A2(n200), .ZN(n517) );
  NAND2_X1 U456 ( .A1(n205), .A2(n200), .ZN(n518) );
  NAND3_X1 U457 ( .A1(n516), .A2(n517), .A3(n518), .ZN(n195) );
  XNOR2_X1 U458 ( .A(n589), .B(a[4]), .ZN(n519) );
  INV_X2 U459 ( .A(n519), .ZN(n16) );
  XNOR2_X1 U460 ( .A(n589), .B(a[4]), .ZN(n520) );
  OR2_X2 U461 ( .A1(n521), .A2(n563), .ZN(n29) );
  XNOR2_X1 U462 ( .A(n594), .B(a[8]), .ZN(n521) );
  OAI21_X1 U463 ( .B1(n89), .B2(n533), .A(n90), .ZN(n522) );
  OR2_X2 U464 ( .A1(n562), .A2(n249), .ZN(n541) );
  INV_X1 U465 ( .A(n544), .ZN(n523) );
  AND2_X1 U466 ( .A1(n269), .A2(n319), .ZN(n193) );
  XOR2_X1 U467 ( .A(n170), .B(n172), .Z(n524) );
  XOR2_X1 U468 ( .A(n524), .B(n179), .Z(n166) );
  XOR2_X1 U469 ( .A(n177), .B(n168), .Z(n525) );
  XOR2_X1 U470 ( .A(n525), .B(n166), .Z(n164) );
  NAND2_X1 U471 ( .A1(n170), .A2(n172), .ZN(n526) );
  NAND2_X1 U472 ( .A1(n170), .A2(n179), .ZN(n527) );
  NAND2_X1 U473 ( .A1(n172), .A2(n179), .ZN(n528) );
  NAND3_X1 U474 ( .A1(n526), .A2(n527), .A3(n528), .ZN(n165) );
  NAND2_X1 U475 ( .A1(n177), .A2(n168), .ZN(n529) );
  NAND2_X1 U476 ( .A1(n177), .A2(n166), .ZN(n530) );
  NAND2_X1 U477 ( .A1(n168), .A2(n166), .ZN(n531) );
  NAND3_X1 U478 ( .A1(n529), .A2(n530), .A3(n531), .ZN(n163) );
  CLKBUF_X1 U479 ( .A(n78), .Z(n532) );
  XOR2_X1 U480 ( .A(n319), .B(n269), .Z(n194) );
  AOI21_X1 U481 ( .B1(n96), .B2(n570), .A(n93), .ZN(n533) );
  AOI21_X1 U482 ( .B1(n571), .B2(n112), .A(n109), .ZN(n534) );
  OAI21_X2 U483 ( .B1(n113), .B2(n115), .A(n114), .ZN(n112) );
  XNOR2_X1 U484 ( .A(n589), .B(a[4]), .ZN(n535) );
  XNOR2_X1 U485 ( .A(n13), .B(a[4]), .ZN(n536) );
  INV_X1 U486 ( .A(n589), .ZN(n537) );
  INV_X1 U487 ( .A(n589), .ZN(n538) );
  INV_X2 U488 ( .A(n7), .ZN(n589) );
  XNOR2_X1 U489 ( .A(n584), .B(a[2]), .ZN(n539) );
  OR2_X2 U490 ( .A1(n562), .A2(n249), .ZN(n540) );
  OR2_X1 U491 ( .A1(n562), .A2(n249), .ZN(n6) );
  NAND2_X1 U492 ( .A1(n196), .A2(n203), .ZN(n86) );
  CLKBUF_X1 U493 ( .A(n499), .Z(n542) );
  BUF_X2 U494 ( .A(n499), .Z(n543) );
  INV_X1 U495 ( .A(n595), .ZN(n594) );
  INV_X1 U496 ( .A(n592), .ZN(n545) );
  INV_X1 U497 ( .A(n128), .ZN(n546) );
  OR2_X1 U498 ( .A1(n176), .A2(n185), .ZN(n547) );
  OR2_X1 U499 ( .A1(n204), .A2(n211), .ZN(n548) );
  INV_X1 U500 ( .A(n597), .ZN(n549) );
  INV_X1 U501 ( .A(n597), .ZN(n550) );
  OAI21_X1 U502 ( .B1(n508), .B2(n534), .A(n106), .ZN(n552) );
  NOR2_X1 U503 ( .A1(n186), .A2(n195), .ZN(n553) );
  CLKBUF_X1 U504 ( .A(n568), .Z(n554) );
  NOR2_X1 U505 ( .A1(n186), .A2(n195), .ZN(n82) );
  OR2_X2 U506 ( .A1(n555), .A2(n564), .ZN(n34) );
  XNOR2_X1 U507 ( .A(n596), .B(a[10]), .ZN(n555) );
  NAND2_X1 U508 ( .A1(n226), .A2(n229), .ZN(n556) );
  NAND2_X1 U509 ( .A1(n226), .A2(n298), .ZN(n557) );
  NAND2_X1 U510 ( .A1(n229), .A2(n298), .ZN(n558) );
  NAND3_X1 U511 ( .A1(n556), .A2(n557), .A3(n558), .ZN(n223) );
  AOI21_X1 U512 ( .B1(n574), .B2(n552), .A(n101), .ZN(n559) );
  INV_X2 U513 ( .A(n591), .ZN(n590) );
  OAI21_X1 U514 ( .B1(n91), .B2(n89), .A(n90), .ZN(n560) );
  OAI21_X1 U515 ( .B1(n91), .B2(n89), .A(n90), .ZN(n88) );
  NOR2_X1 U516 ( .A1(n164), .A2(n175), .ZN(n561) );
  NOR2_X1 U517 ( .A1(n164), .A2(n175), .ZN(n75) );
  BUF_X2 U518 ( .A(n9), .Z(n579) );
  XNOR2_X1 U519 ( .A(n584), .B(n249), .ZN(n562) );
  XNOR2_X1 U520 ( .A(n593), .B(a[8]), .ZN(n563) );
  INV_X1 U521 ( .A(n564), .ZN(n32) );
  XNOR2_X1 U522 ( .A(n595), .B(a[10]), .ZN(n564) );
  XNOR2_X1 U523 ( .A(n560), .B(n51), .ZN(product[10]) );
  INV_X1 U524 ( .A(n589), .ZN(n587) );
  XNOR2_X1 U525 ( .A(n589), .B(a[2]), .ZN(n567) );
  INV_X2 U526 ( .A(n593), .ZN(n592) );
  NAND2_X1 U527 ( .A1(n539), .A2(n567), .ZN(n565) );
  INV_X1 U528 ( .A(n249), .ZN(n566) );
  NAND2_X1 U529 ( .A1(n567), .A2(n539), .ZN(n12) );
  BUF_X1 U530 ( .A(n43), .Z(n582) );
  AOI21_X1 U531 ( .B1(n560), .B2(n491), .A(n81), .ZN(n568) );
  NAND2_X1 U532 ( .A1(n569), .A2(n69), .ZN(n47) );
  INV_X1 U533 ( .A(n73), .ZN(n71) );
  AOI21_X1 U534 ( .B1(n569), .B2(n74), .A(n67), .ZN(n65) );
  INV_X1 U535 ( .A(n69), .ZN(n67) );
  INV_X1 U536 ( .A(n74), .ZN(n72) );
  INV_X1 U537 ( .A(n95), .ZN(n93) );
  AOI21_X1 U538 ( .B1(n522), .B2(n80), .A(n81), .ZN(n45) );
  NOR2_X1 U539 ( .A1(n553), .A2(n85), .ZN(n80) );
  OAI21_X1 U540 ( .B1(n82), .B2(n86), .A(n83), .ZN(n81) );
  NAND2_X1 U541 ( .A1(n128), .A2(n86), .ZN(n51) );
  INV_X1 U542 ( .A(n85), .ZN(n128) );
  NAND2_X1 U543 ( .A1(n548), .A2(n90), .ZN(n52) );
  OR2_X1 U544 ( .A1(n152), .A2(n163), .ZN(n569) );
  NAND2_X1 U545 ( .A1(n496), .A2(n570), .ZN(n53) );
  OAI21_X1 U546 ( .B1(n561), .B2(n79), .A(n76), .ZN(n74) );
  NAND2_X1 U547 ( .A1(n125), .A2(n76), .ZN(n48) );
  INV_X1 U548 ( .A(n75), .ZN(n125) );
  NOR2_X1 U549 ( .A1(n75), .A2(n78), .ZN(n73) );
  XNOR2_X1 U550 ( .A(n84), .B(n50), .ZN(product[11]) );
  NAND2_X1 U551 ( .A1(n127), .A2(n83), .ZN(n50) );
  INV_X1 U552 ( .A(n553), .ZN(n127) );
  NAND2_X1 U553 ( .A1(n152), .A2(n163), .ZN(n69) );
  INV_X1 U554 ( .A(n119), .ZN(n117) );
  AOI21_X1 U555 ( .B1(n571), .B2(n112), .A(n109), .ZN(n107) );
  INV_X1 U556 ( .A(n103), .ZN(n101) );
  NAND2_X1 U557 ( .A1(n131), .A2(n98), .ZN(n54) );
  INV_X1 U558 ( .A(n97), .ZN(n131) );
  OR2_X1 U559 ( .A1(n212), .A2(n217), .ZN(n570) );
  NOR2_X1 U560 ( .A1(n176), .A2(n185), .ZN(n78) );
  NOR2_X1 U561 ( .A1(n196), .A2(n203), .ZN(n85) );
  NAND2_X1 U562 ( .A1(n573), .A2(n119), .ZN(n59) );
  XOR2_X1 U563 ( .A(n56), .B(n534), .Z(product[5]) );
  NAND2_X1 U564 ( .A1(n133), .A2(n106), .ZN(n56) );
  INV_X1 U565 ( .A(n508), .ZN(n133) );
  OAI21_X1 U566 ( .B1(n105), .B2(n107), .A(n106), .ZN(n104) );
  NAND2_X1 U567 ( .A1(n176), .A2(n185), .ZN(n79) );
  NAND2_X1 U568 ( .A1(n164), .A2(n175), .ZN(n76) );
  NAND2_X1 U569 ( .A1(n186), .A2(n195), .ZN(n83) );
  NAND2_X1 U570 ( .A1(n204), .A2(n211), .ZN(n90) );
  INV_X1 U571 ( .A(n113), .ZN(n135) );
  XNOR2_X1 U572 ( .A(n63), .B(n46), .ZN(product[15]) );
  NAND2_X1 U573 ( .A1(n572), .A2(n62), .ZN(n46) );
  NAND2_X1 U574 ( .A1(n490), .A2(n569), .ZN(n64) );
  XNOR2_X1 U575 ( .A(n57), .B(n112), .ZN(product[4]) );
  NAND2_X1 U576 ( .A1(n571), .A2(n111), .ZN(n57) );
  XNOR2_X1 U577 ( .A(n55), .B(n552), .ZN(product[6]) );
  NAND2_X1 U578 ( .A1(n574), .A2(n103), .ZN(n55) );
  OR2_X1 U579 ( .A1(n232), .A2(n233), .ZN(n571) );
  OR2_X1 U580 ( .A1(n139), .A2(n151), .ZN(n572) );
  NAND2_X1 U581 ( .A1(n228), .A2(n231), .ZN(n106) );
  INV_X1 U582 ( .A(n37), .ZN(n237) );
  NAND2_X1 U583 ( .A1(n224), .A2(n227), .ZN(n103) );
  OR2_X1 U584 ( .A1(n328), .A2(n314), .ZN(n573) );
  OR2_X1 U585 ( .A1(n224), .A2(n227), .ZN(n574) );
  NAND2_X1 U586 ( .A1(n218), .A2(n223), .ZN(n98) );
  INV_X1 U587 ( .A(n41), .ZN(n235) );
  AND2_X1 U588 ( .A1(n494), .A2(n122), .ZN(product[1]) );
  XNOR2_X1 U589 ( .A(n596), .B(a[12]), .ZN(n37) );
  XNOR2_X1 U590 ( .A(n598), .B(a[14]), .ZN(n41) );
  OR2_X1 U591 ( .A1(n582), .A2(n589), .ZN(n392) );
  AND2_X1 U592 ( .A1(n506), .A2(n583), .ZN(n288) );
  OAI22_X1 U593 ( .A1(n39), .A2(n336), .B1(n37), .B2(n335), .ZN(n263) );
  XNOR2_X1 U594 ( .A(n544), .B(n582), .ZN(n352) );
  XNOR2_X1 U595 ( .A(n155), .B(n576), .ZN(n139) );
  XNOR2_X1 U596 ( .A(n153), .B(n141), .ZN(n576) );
  XNOR2_X1 U597 ( .A(n157), .B(n577), .ZN(n141) );
  XNOR2_X1 U598 ( .A(n145), .B(n143), .ZN(n577) );
  OAI22_X1 U599 ( .A1(n42), .A2(n601), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U600 ( .A1(n582), .A2(n601), .ZN(n332) );
  XNOR2_X1 U601 ( .A(n590), .B(n582), .ZN(n376) );
  XNOR2_X1 U602 ( .A(n549), .B(n582), .ZN(n343) );
  XNOR2_X1 U603 ( .A(n159), .B(n578), .ZN(n142) );
  XNOR2_X1 U604 ( .A(n315), .B(n261), .ZN(n578) );
  XNOR2_X1 U605 ( .A(n598), .B(n582), .ZN(n336) );
  NAND2_X1 U606 ( .A1(n427), .A2(n37), .ZN(n39) );
  XOR2_X1 U607 ( .A(n598), .B(a[12]), .Z(n427) );
  AND2_X1 U608 ( .A1(n583), .A2(n535), .ZN(n300) );
  AND2_X1 U609 ( .A1(n583), .A2(n237), .ZN(n264) );
  AND2_X1 U610 ( .A1(n583), .A2(n564), .ZN(n270) );
  AND2_X1 U611 ( .A1(n583), .A2(n235), .ZN(n260) );
  OAI22_X1 U612 ( .A1(n39), .A2(n335), .B1(n37), .B2(n334), .ZN(n262) );
  INV_X1 U613 ( .A(n19), .ZN(n593) );
  INV_X1 U614 ( .A(n25), .ZN(n595) );
  AND2_X1 U615 ( .A1(n583), .A2(n563), .ZN(n278) );
  NAND2_X1 U616 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U617 ( .A(n600), .B(a[14]), .Z(n426) );
  OAI22_X1 U618 ( .A1(n39), .A2(n599), .B1(n337), .B2(n37), .ZN(n252) );
  OR2_X1 U619 ( .A1(n582), .A2(n599), .ZN(n337) );
  XNOR2_X1 U620 ( .A(n592), .B(n582), .ZN(n363) );
  AND2_X1 U621 ( .A1(n583), .A2(n247), .ZN(n314) );
  AND2_X1 U622 ( .A1(n583), .A2(n249), .ZN(product[0]) );
  OR2_X1 U623 ( .A1(n582), .A2(n597), .ZN(n344) );
  OR2_X1 U624 ( .A1(n582), .A2(n523), .ZN(n353) );
  OR2_X1 U625 ( .A1(n582), .A2(n545), .ZN(n364) );
  OR2_X1 U626 ( .A1(n582), .A2(n591), .ZN(n377) );
  XNOR2_X1 U627 ( .A(n592), .B(b[9]), .ZN(n354) );
  OAI22_X1 U628 ( .A1(n39), .A2(n334), .B1(n37), .B2(n333), .ZN(n261) );
  XNOR2_X1 U629 ( .A(n598), .B(n422), .ZN(n333) );
  XNOR2_X1 U630 ( .A(n590), .B(b[11]), .ZN(n365) );
  XNOR2_X1 U631 ( .A(n598), .B(n424), .ZN(n335) );
  XNOR2_X1 U632 ( .A(n598), .B(n423), .ZN(n334) );
  OAI22_X1 U633 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U634 ( .A(n600), .B(n424), .ZN(n330) );
  XNOR2_X1 U635 ( .A(n600), .B(n582), .ZN(n331) );
  XNOR2_X1 U636 ( .A(n544), .B(n418), .ZN(n345) );
  XNOR2_X1 U637 ( .A(n549), .B(n420), .ZN(n338) );
  XNOR2_X1 U638 ( .A(n587), .B(b[13]), .ZN(n378) );
  XNOR2_X1 U639 ( .A(n594), .B(n424), .ZN(n351) );
  XNOR2_X1 U640 ( .A(n550), .B(n424), .ZN(n342) );
  XNOR2_X1 U641 ( .A(n592), .B(n424), .ZN(n362) );
  XNOR2_X1 U642 ( .A(n550), .B(n423), .ZN(n341) );
  XNOR2_X1 U643 ( .A(n549), .B(n422), .ZN(n340) );
  XNOR2_X1 U644 ( .A(n550), .B(n421), .ZN(n339) );
  XNOR2_X1 U645 ( .A(n588), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U646 ( .A(n588), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U647 ( .A(n538), .B(n418), .ZN(n384) );
  XNOR2_X1 U648 ( .A(n537), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U649 ( .A(n537), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U650 ( .A(n538), .B(n419), .ZN(n385) );
  XNOR2_X1 U651 ( .A(n537), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U652 ( .A(n592), .B(n422), .ZN(n360) );
  XNOR2_X1 U653 ( .A(n544), .B(n422), .ZN(n349) );
  XNOR2_X1 U654 ( .A(n590), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U655 ( .A(n590), .B(n418), .ZN(n369) );
  XNOR2_X1 U656 ( .A(n590), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U657 ( .A(n590), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U658 ( .A(n592), .B(n423), .ZN(n361) );
  XNOR2_X1 U659 ( .A(n544), .B(n423), .ZN(n350) );
  XNOR2_X1 U660 ( .A(n592), .B(n420), .ZN(n358) );
  XNOR2_X1 U661 ( .A(n544), .B(n420), .ZN(n347) );
  XNOR2_X1 U662 ( .A(n592), .B(n421), .ZN(n359) );
  XNOR2_X1 U663 ( .A(n594), .B(n421), .ZN(n348) );
  XNOR2_X1 U664 ( .A(n592), .B(n419), .ZN(n357) );
  XNOR2_X1 U665 ( .A(n544), .B(n419), .ZN(n346) );
  XNOR2_X1 U666 ( .A(n592), .B(n418), .ZN(n356) );
  XNOR2_X1 U667 ( .A(n592), .B(b[8]), .ZN(n355) );
  XNOR2_X1 U668 ( .A(n503), .B(b[11]), .ZN(n397) );
  XNOR2_X1 U669 ( .A(n503), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U670 ( .A(n502), .B(b[13]), .ZN(n395) );
  XNOR2_X1 U671 ( .A(n503), .B(b[14]), .ZN(n394) );
  BUF_X1 U672 ( .A(n43), .Z(n583) );
  XNOR2_X1 U673 ( .A(n502), .B(b[15]), .ZN(n393) );
  XNOR2_X1 U674 ( .A(n584), .B(a[2]), .ZN(n9) );
  NAND2_X1 U675 ( .A1(n212), .A2(n217), .ZN(n95) );
  INV_X1 U676 ( .A(n13), .ZN(n591) );
  NOR2_X1 U677 ( .A1(n218), .A2(n223), .ZN(n97) );
  OAI22_X1 U678 ( .A1(n34), .A2(n339), .B1(n338), .B2(n32), .ZN(n265) );
  OAI22_X1 U679 ( .A1(n34), .A2(n340), .B1(n339), .B2(n32), .ZN(n266) );
  OAI22_X1 U680 ( .A1(n34), .A2(n342), .B1(n341), .B2(n32), .ZN(n268) );
  OAI22_X1 U681 ( .A1(n34), .A2(n341), .B1(n340), .B2(n32), .ZN(n267) );
  OAI22_X1 U682 ( .A1(n34), .A2(n343), .B1(n342), .B2(n32), .ZN(n269) );
  OAI22_X1 U683 ( .A1(n34), .A2(n597), .B1(n344), .B2(n32), .ZN(n253) );
  INV_X1 U684 ( .A(n503), .ZN(n581) );
  XOR2_X1 U685 ( .A(n58), .B(n505), .Z(product[3]) );
  OAI22_X1 U686 ( .A1(n541), .A2(n395), .B1(n394), .B2(n566), .ZN(n316) );
  OAI22_X1 U687 ( .A1(n540), .A2(n394), .B1(n393), .B2(n566), .ZN(n315) );
  NAND2_X1 U688 ( .A1(n328), .A2(n314), .ZN(n119) );
  OAI22_X1 U689 ( .A1(n541), .A2(n400), .B1(n399), .B2(n566), .ZN(n321) );
  OAI22_X1 U690 ( .A1(n541), .A2(n401), .B1(n400), .B2(n566), .ZN(n322) );
  OAI22_X1 U691 ( .A1(n540), .A2(n397), .B1(n396), .B2(n566), .ZN(n318) );
  OAI22_X1 U692 ( .A1(n540), .A2(n396), .B1(n395), .B2(n566), .ZN(n317) );
  OAI22_X1 U693 ( .A1(n540), .A2(n398), .B1(n397), .B2(n566), .ZN(n319) );
  OAI22_X1 U694 ( .A1(n541), .A2(n406), .B1(n405), .B2(n566), .ZN(n327) );
  OAI22_X1 U695 ( .A1(n6), .A2(n399), .B1(n398), .B2(n566), .ZN(n320) );
  OAI22_X1 U696 ( .A1(n541), .A2(n402), .B1(n401), .B2(n566), .ZN(n323) );
  OAI22_X1 U697 ( .A1(n6), .A2(n404), .B1(n403), .B2(n566), .ZN(n325) );
  OAI22_X1 U698 ( .A1(n541), .A2(n408), .B1(n407), .B2(n566), .ZN(n329) );
  OAI22_X1 U699 ( .A1(n540), .A2(n403), .B1(n402), .B2(n566), .ZN(n324) );
  OAI22_X1 U700 ( .A1(n6), .A2(n405), .B1(n404), .B2(n566), .ZN(n326) );
  OAI22_X1 U701 ( .A1(n540), .A2(n407), .B1(n406), .B2(n566), .ZN(n328) );
  NOR2_X1 U702 ( .A1(n204), .A2(n211), .ZN(n89) );
  OAI22_X1 U703 ( .A1(n29), .A2(n346), .B1(n345), .B2(n27), .ZN(n271) );
  OAI22_X1 U704 ( .A1(n29), .A2(n350), .B1(n349), .B2(n27), .ZN(n275) );
  OAI22_X1 U705 ( .A1(n29), .A2(n347), .B1(n346), .B2(n27), .ZN(n272) );
  OAI22_X1 U706 ( .A1(n29), .A2(n348), .B1(n347), .B2(n27), .ZN(n273) );
  OAI22_X1 U707 ( .A1(n29), .A2(n351), .B1(n350), .B2(n27), .ZN(n276) );
  OAI22_X1 U708 ( .A1(n29), .A2(n349), .B1(n348), .B2(n27), .ZN(n274) );
  OAI22_X1 U709 ( .A1(n29), .A2(n523), .B1(n353), .B2(n27), .ZN(n254) );
  OAI22_X1 U710 ( .A1(n29), .A2(n352), .B1(n351), .B2(n27), .ZN(n277) );
  INV_X1 U711 ( .A(n586), .ZN(n584) );
  XNOR2_X1 U712 ( .A(n590), .B(n424), .ZN(n375) );
  XNOR2_X1 U713 ( .A(n590), .B(n419), .ZN(n370) );
  XNOR2_X1 U714 ( .A(n590), .B(n420), .ZN(n371) );
  XNOR2_X1 U715 ( .A(n590), .B(n423), .ZN(n374) );
  XNOR2_X1 U716 ( .A(n590), .B(n422), .ZN(n373) );
  XNOR2_X1 U717 ( .A(n590), .B(n421), .ZN(n372) );
  INV_X1 U718 ( .A(n1), .ZN(n586) );
  OR2_X1 U719 ( .A1(n582), .A2(n581), .ZN(n409) );
  XNOR2_X1 U720 ( .A(n70), .B(n47), .ZN(product[14]) );
  OAI21_X1 U721 ( .B1(n87), .B2(n546), .A(n86), .ZN(n84) );
  NOR2_X1 U722 ( .A1(n234), .A2(n257), .ZN(n113) );
  INV_X1 U723 ( .A(n111), .ZN(n109) );
  OAI22_X1 U724 ( .A1(n23), .A2(n356), .B1(n355), .B2(n543), .ZN(n280) );
  OAI22_X1 U725 ( .A1(n23), .A2(n358), .B1(n357), .B2(n543), .ZN(n282) );
  OAI22_X1 U726 ( .A1(n23), .A2(n355), .B1(n354), .B2(n543), .ZN(n279) );
  OAI22_X1 U727 ( .A1(n23), .A2(n362), .B1(n361), .B2(n543), .ZN(n286) );
  OAI22_X1 U728 ( .A1(n23), .A2(n360), .B1(n359), .B2(n543), .ZN(n284) );
  OAI22_X1 U729 ( .A1(n23), .A2(n361), .B1(n360), .B2(n543), .ZN(n285) );
  OAI22_X1 U730 ( .A1(n23), .A2(n545), .B1(n364), .B2(n543), .ZN(n255) );
  OAI22_X1 U731 ( .A1(n23), .A2(n357), .B1(n356), .B2(n543), .ZN(n281) );
  OAI22_X1 U732 ( .A1(n23), .A2(n363), .B1(n362), .B2(n543), .ZN(n287) );
  OAI22_X1 U733 ( .A1(n359), .A2(n23), .B1(n358), .B2(n542), .ZN(n283) );
  NAND2_X1 U734 ( .A1(n151), .A2(n139), .ZN(n62) );
  INV_X1 U735 ( .A(n88), .ZN(n87) );
  XNOR2_X1 U736 ( .A(n77), .B(n48), .ZN(product[13]) );
  NAND2_X1 U737 ( .A1(n232), .A2(n233), .ZN(n111) );
  XNOR2_X1 U738 ( .A(n502), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U739 ( .A(n502), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U740 ( .A(n503), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U741 ( .A(n501), .B(n418), .ZN(n401) );
  XNOR2_X1 U742 ( .A(n503), .B(n582), .ZN(n408) );
  XNOR2_X1 U743 ( .A(n502), .B(n419), .ZN(n402) );
  XNOR2_X1 U744 ( .A(n501), .B(n420), .ZN(n403) );
  XNOR2_X1 U745 ( .A(n502), .B(n423), .ZN(n406) );
  XNOR2_X1 U746 ( .A(n502), .B(n424), .ZN(n407) );
  XNOR2_X1 U747 ( .A(n503), .B(n422), .ZN(n405) );
  XNOR2_X1 U748 ( .A(n501), .B(n421), .ZN(n404) );
  OAI22_X1 U749 ( .A1(n18), .A2(n370), .B1(n369), .B2(n16), .ZN(n293) );
  OAI22_X1 U750 ( .A1(n18), .A2(n367), .B1(n366), .B2(n16), .ZN(n290) );
  OAI22_X1 U751 ( .A1(n18), .A2(n375), .B1(n374), .B2(n16), .ZN(n298) );
  OAI22_X1 U752 ( .A1(n18), .A2(n368), .B1(n367), .B2(n16), .ZN(n291) );
  OAI22_X1 U753 ( .A1(n18), .A2(n372), .B1(n371), .B2(n16), .ZN(n295) );
  OAI22_X1 U754 ( .A1(n18), .A2(n373), .B1(n372), .B2(n16), .ZN(n296) );
  OAI22_X1 U755 ( .A1(n18), .A2(n374), .B1(n373), .B2(n16), .ZN(n297) );
  OAI22_X1 U756 ( .A1(n18), .A2(n369), .B1(n368), .B2(n16), .ZN(n292) );
  OAI22_X1 U757 ( .A1(n18), .A2(n376), .B1(n375), .B2(n16), .ZN(n299) );
  OAI22_X1 U758 ( .A1(n18), .A2(n591), .B1(n377), .B2(n16), .ZN(n256) );
  OAI22_X1 U759 ( .A1(n18), .A2(n371), .B1(n370), .B2(n16), .ZN(n294) );
  OAI22_X1 U760 ( .A1(n18), .A2(n366), .B1(n365), .B2(n16), .ZN(n289) );
  XNOR2_X1 U761 ( .A(n538), .B(n420), .ZN(n386) );
  XNOR2_X1 U762 ( .A(n587), .B(n421), .ZN(n387) );
  XNOR2_X1 U763 ( .A(n587), .B(n582), .ZN(n391) );
  XNOR2_X1 U764 ( .A(n588), .B(n422), .ZN(n388) );
  XNOR2_X1 U765 ( .A(n587), .B(n424), .ZN(n390) );
  XNOR2_X1 U766 ( .A(n537), .B(n423), .ZN(n389) );
  NAND2_X1 U767 ( .A1(n135), .A2(n114), .ZN(n58) );
  OAI21_X1 U768 ( .B1(n568), .B2(n71), .A(n72), .ZN(n70) );
  OAI21_X1 U769 ( .B1(n45), .B2(n532), .A(n79), .ZN(n77) );
  OAI21_X1 U770 ( .B1(n64), .B2(n554), .A(n65), .ZN(n63) );
  XOR2_X1 U771 ( .A(n533), .B(n52), .Z(product[9]) );
  XNOR2_X1 U772 ( .A(n551), .B(n53), .ZN(product[8]) );
  AOI21_X1 U773 ( .B1(n96), .B2(n570), .A(n93), .ZN(n91) );
  XNOR2_X1 U774 ( .A(n59), .B(n120), .ZN(product[2]) );
  AOI21_X1 U775 ( .B1(n573), .B2(n120), .A(n117), .ZN(n115) );
  INV_X1 U776 ( .A(n122), .ZN(n120) );
  NAND2_X1 U777 ( .A1(n329), .A2(n258), .ZN(n122) );
  OAI21_X1 U778 ( .B1(n99), .B2(n97), .A(n98), .ZN(n96) );
  AOI21_X1 U779 ( .B1(n104), .B2(n574), .A(n101), .ZN(n99) );
  OAI22_X1 U780 ( .A1(n540), .A2(n581), .B1(n409), .B2(n566), .ZN(n258) );
  XOR2_X1 U781 ( .A(n559), .B(n54), .Z(product[7]) );
  OAI22_X1 U782 ( .A1(n507), .A2(n379), .B1(n378), .B2(n495), .ZN(n301) );
  OAI22_X1 U783 ( .A1(n507), .A2(n380), .B1(n379), .B2(n579), .ZN(n302) );
  OAI22_X1 U784 ( .A1(n510), .A2(n385), .B1(n495), .B2(n384), .ZN(n307) );
  OAI22_X1 U785 ( .A1(n507), .A2(n382), .B1(n381), .B2(n495), .ZN(n304) );
  OAI22_X1 U786 ( .A1(n507), .A2(n381), .B1(n380), .B2(n495), .ZN(n303) );
  NAND2_X1 U787 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U788 ( .A1(n565), .A2(n383), .B1(n382), .B2(n580), .ZN(n305) );
  OAI22_X1 U789 ( .A1(n12), .A2(n384), .B1(n383), .B2(n495), .ZN(n306) );
  OAI22_X1 U790 ( .A1(n510), .A2(n386), .B1(n385), .B2(n579), .ZN(n308) );
  OAI22_X1 U791 ( .A1(n507), .A2(n387), .B1(n386), .B2(n495), .ZN(n309) );
  OAI22_X1 U792 ( .A1(n507), .A2(n589), .B1(n392), .B2(n579), .ZN(n257) );
  OAI22_X1 U793 ( .A1(n565), .A2(n389), .B1(n388), .B2(n580), .ZN(n311) );
  OAI22_X1 U794 ( .A1(n12), .A2(n388), .B1(n387), .B2(n579), .ZN(n310) );
  OAI22_X1 U795 ( .A1(n12), .A2(n390), .B1(n389), .B2(n579), .ZN(n312) );
  INV_X1 U796 ( .A(n579), .ZN(n247) );
  OAI22_X1 U797 ( .A1(n12), .A2(n391), .B1(n390), .B2(n495), .ZN(n313) );
  INV_X1 U798 ( .A(n589), .ZN(n588) );
  INV_X1 U799 ( .A(n597), .ZN(n596) );
  INV_X1 U800 ( .A(n31), .ZN(n597) );
  INV_X1 U801 ( .A(n599), .ZN(n598) );
  INV_X1 U802 ( .A(n36), .ZN(n599) );
  INV_X1 U803 ( .A(n601), .ZN(n600) );
  INV_X1 U804 ( .A(n40), .ZN(n601) );
  XOR2_X1 U805 ( .A(n259), .B(n251), .Z(n148) );
  XOR2_X1 U806 ( .A(n149), .B(n147), .Z(n144) );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_14_DW01_add_2 ( A, B, CI, 
        SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n5, n9, n10, n11, n12, n13, n14, n15, n16, n19, n20, n22, n24,
         n25, n26, n27, n28, n29, n30, n32, n33, n34, n35, n36, n37, n39, n40,
         n44, n45, n47, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n65, n67, n68, n69, n70, n71, n73, n75, n76, n77,
         n78, n79, n81, n83, n84, n86, n89, n90, n91, n94, n95, n96, n98, n100,
         n157, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182;

  INV_X1 U122 ( .A(n89), .ZN(n157) );
  NOR2_X2 U123 ( .A1(A[11]), .A2(B[11]), .ZN(n35) );
  NOR2_X1 U124 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  AND2_X1 U125 ( .A1(n176), .A2(n86), .ZN(SUM[0]) );
  XNOR2_X1 U126 ( .A(n51), .B(n159), .ZN(SUM[9]) );
  AND2_X1 U127 ( .A1(n177), .A2(n49), .ZN(n159) );
  XNOR2_X1 U128 ( .A(n45), .B(n160), .ZN(SUM[10]) );
  AND2_X1 U129 ( .A1(n180), .A2(n44), .ZN(n160) );
  OR2_X1 U130 ( .A1(A[15]), .A2(B[15]), .ZN(n161) );
  XNOR2_X1 U131 ( .A(n37), .B(n162), .ZN(SUM[11]) );
  AND2_X1 U132 ( .A1(n91), .A2(n36), .ZN(n162) );
  OAI21_X1 U133 ( .B1(n32), .B2(n36), .A(n33), .ZN(n163) );
  BUF_X1 U134 ( .A(n26), .Z(n164) );
  OR2_X1 U135 ( .A1(n25), .A2(n28), .ZN(n165) );
  AOI21_X1 U136 ( .B1(n180), .B2(n47), .A(n182), .ZN(n166) );
  NOR2_X1 U137 ( .A1(A[8]), .A2(B[8]), .ZN(n167) );
  OAI21_X1 U138 ( .B1(n39), .B2(n51), .A(n40), .ZN(n168) );
  AOI21_X2 U139 ( .B1(n52), .B2(n60), .A(n53), .ZN(n51) );
  NOR2_X1 U140 ( .A1(A[14]), .A2(B[14]), .ZN(n169) );
  XNOR2_X1 U141 ( .A(n175), .B(n170), .ZN(SUM[13]) );
  AND2_X1 U142 ( .A1(n89), .A2(n29), .ZN(n170) );
  OAI21_X1 U143 ( .B1(n39), .B2(n51), .A(n166), .ZN(n171) );
  OR2_X1 U144 ( .A1(A[14]), .A2(B[14]), .ZN(n172) );
  NOR2_X1 U145 ( .A1(A[14]), .A2(B[14]), .ZN(n25) );
  OR2_X2 U146 ( .A1(A[10]), .A2(B[10]), .ZN(n180) );
  NOR2_X1 U147 ( .A1(A[12]), .A2(B[12]), .ZN(n173) );
  NOR2_X1 U148 ( .A1(A[12]), .A2(B[12]), .ZN(n32) );
  AOI21_X1 U149 ( .B1(n171), .B2(n30), .A(n163), .ZN(n174) );
  AOI21_X1 U150 ( .B1(n168), .B2(n30), .A(n163), .ZN(n175) );
  OR2_X1 U151 ( .A1(A[0]), .A2(B[0]), .ZN(n176) );
  INV_X1 U152 ( .A(n60), .ZN(n59) );
  INV_X1 U153 ( .A(n51), .ZN(n50) );
  INV_X1 U154 ( .A(n168), .ZN(n37) );
  OAI21_X1 U155 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  AOI21_X1 U156 ( .B1(n181), .B2(n68), .A(n65), .ZN(n63) );
  INV_X1 U157 ( .A(n67), .ZN(n65) );
  AOI21_X1 U158 ( .B1(n178), .B2(n76), .A(n73), .ZN(n71) );
  INV_X1 U159 ( .A(n75), .ZN(n73) );
  OAI21_X1 U160 ( .B1(n79), .B2(n77), .A(n78), .ZN(n76) );
  INV_X1 U161 ( .A(n24), .ZN(n22) );
  OAI21_X1 U162 ( .B1(n71), .B2(n69), .A(n70), .ZN(n68) );
  AOI21_X1 U163 ( .B1(n50), .B2(n177), .A(n47), .ZN(n45) );
  NAND2_X1 U164 ( .A1(n94), .A2(n55), .ZN(n9) );
  INV_X1 U165 ( .A(n86), .ZN(n84) );
  OAI21_X1 U166 ( .B1(n59), .B2(n57), .A(n58), .ZN(n56) );
  INV_X1 U167 ( .A(n49), .ZN(n47) );
  AOI21_X1 U168 ( .B1(n179), .B2(n84), .A(n81), .ZN(n79) );
  INV_X1 U169 ( .A(n83), .ZN(n81) );
  NAND2_X1 U170 ( .A1(n95), .A2(n58), .ZN(n10) );
  INV_X1 U171 ( .A(n57), .ZN(n95) );
  NAND2_X1 U172 ( .A1(n98), .A2(n70), .ZN(n13) );
  INV_X1 U173 ( .A(n69), .ZN(n98) );
  NAND2_X1 U174 ( .A1(n96), .A2(n62), .ZN(n11) );
  INV_X1 U175 ( .A(n61), .ZN(n96) );
  INV_X1 U176 ( .A(n173), .ZN(n90) );
  INV_X1 U177 ( .A(n28), .ZN(n89) );
  NAND2_X1 U178 ( .A1(n100), .A2(n78), .ZN(n15) );
  INV_X1 U179 ( .A(n77), .ZN(n100) );
  NAND2_X1 U180 ( .A1(n181), .A2(n67), .ZN(n12) );
  NAND2_X1 U181 ( .A1(n178), .A2(n75), .ZN(n14) );
  NAND2_X1 U182 ( .A1(n179), .A2(n83), .ZN(n16) );
  INV_X1 U183 ( .A(n182), .ZN(n44) );
  XNOR2_X1 U184 ( .A(n34), .B(n5), .ZN(SUM[12]) );
  NAND2_X1 U185 ( .A1(n33), .A2(n90), .ZN(n5) );
  XOR2_X1 U186 ( .A(n59), .B(n10), .Z(SUM[7]) );
  XNOR2_X1 U187 ( .A(n12), .B(n68), .ZN(SUM[5]) );
  XOR2_X1 U188 ( .A(n13), .B(n71), .Z(SUM[4]) );
  NOR2_X1 U189 ( .A1(A[7]), .A2(B[7]), .ZN(n57) );
  OR2_X1 U190 ( .A1(A[9]), .A2(B[9]), .ZN(n177) );
  NOR2_X1 U191 ( .A1(A[4]), .A2(B[4]), .ZN(n69) );
  NOR2_X1 U192 ( .A1(A[2]), .A2(B[2]), .ZN(n77) );
  NAND2_X1 U193 ( .A1(n172), .A2(n164), .ZN(n3) );
  OR2_X1 U194 ( .A1(A[3]), .A2(B[3]), .ZN(n178) );
  OR2_X1 U195 ( .A1(A[1]), .A2(B[1]), .ZN(n179) );
  NAND2_X1 U196 ( .A1(n161), .A2(n19), .ZN(n2) );
  NOR2_X1 U197 ( .A1(A[6]), .A2(B[6]), .ZN(n61) );
  NOR2_X1 U198 ( .A1(A[8]), .A2(B[8]), .ZN(n54) );
  XNOR2_X1 U199 ( .A(n56), .B(n9), .ZN(SUM[8]) );
  XNOR2_X1 U200 ( .A(n14), .B(n76), .ZN(SUM[3]) );
  XNOR2_X1 U201 ( .A(n16), .B(n84), .ZN(SUM[1]) );
  NAND2_X1 U202 ( .A1(A[7]), .A2(B[7]), .ZN(n58) );
  OR2_X1 U203 ( .A1(A[5]), .A2(B[5]), .ZN(n181) );
  NAND2_X1 U204 ( .A1(A[4]), .A2(B[4]), .ZN(n70) );
  NAND2_X1 U205 ( .A1(A[2]), .A2(B[2]), .ZN(n78) );
  NAND2_X1 U206 ( .A1(A[9]), .A2(B[9]), .ZN(n49) );
  NAND2_X1 U207 ( .A1(A[5]), .A2(B[5]), .ZN(n67) );
  NAND2_X1 U208 ( .A1(A[1]), .A2(B[1]), .ZN(n83) );
  NAND2_X1 U209 ( .A1(A[3]), .A2(B[3]), .ZN(n75) );
  NAND2_X1 U210 ( .A1(A[0]), .A2(B[0]), .ZN(n86) );
  NAND2_X1 U211 ( .A1(A[6]), .A2(B[6]), .ZN(n62) );
  NAND2_X1 U212 ( .A1(A[8]), .A2(B[8]), .ZN(n55) );
  NAND2_X1 U213 ( .A1(A[14]), .A2(B[14]), .ZN(n26) );
  XOR2_X1 U214 ( .A(n11), .B(n63), .Z(SUM[6]) );
  XOR2_X1 U215 ( .A(n15), .B(n79), .Z(SUM[2]) );
  AND2_X1 U216 ( .A1(A[10]), .A2(B[10]), .ZN(n182) );
  NAND2_X1 U217 ( .A1(A[13]), .A2(B[13]), .ZN(n29) );
  NAND2_X1 U218 ( .A1(A[12]), .A2(B[12]), .ZN(n33) );
  INV_X1 U219 ( .A(n167), .ZN(n94) );
  NOR2_X1 U220 ( .A1(n167), .A2(n57), .ZN(n52) );
  OAI21_X1 U221 ( .B1(n54), .B2(n58), .A(n55), .ZN(n53) );
  AOI21_X1 U222 ( .B1(n180), .B2(n47), .A(n182), .ZN(n40) );
  NAND2_X1 U223 ( .A1(A[11]), .A2(B[11]), .ZN(n36) );
  OAI21_X1 U224 ( .B1(n37), .B2(n35), .A(n36), .ZN(n34) );
  INV_X1 U225 ( .A(n35), .ZN(n91) );
  NOR2_X1 U226 ( .A1(n173), .A2(n35), .ZN(n30) );
  NAND2_X1 U227 ( .A1(A[15]), .A2(B[15]), .ZN(n19) );
  OAI21_X1 U228 ( .B1(n169), .B2(n29), .A(n26), .ZN(n24) );
  NAND2_X1 U229 ( .A1(n180), .A2(n177), .ZN(n39) );
  XNOR2_X1 U230 ( .A(n20), .B(n2), .ZN(SUM[15]) );
  XNOR2_X1 U231 ( .A(n27), .B(n3), .ZN(SUM[14]) );
  OAI21_X1 U232 ( .B1(n175), .B2(n157), .A(n29), .ZN(n27) );
  OAI21_X1 U233 ( .B1(n174), .B2(n165), .A(n22), .ZN(n20) );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_14 ( clk, clear_acc, 
        data_out_x, data_out, data_out_w, data_out_b, wr_en_y, m_valid, 
        m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [4:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
         N39, N40, N41, N42, N43, N44, n1, n2, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n85, n102, n111, n112, n113, n114, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n22), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n223), .CK(clk), .Q(n25) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n224), .CK(clk), .Q(n26) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n225), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n226), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n227), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n228), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n229), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n230), .CK(clk), .Q(n34) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n231), .CK(clk), .Q(n35) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n232), .CK(clk), .Q(n36) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n233), .CK(clk), .Q(n37) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n234), .CK(clk), .Q(n38) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n235), .CK(clk), .Q(n39) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n236), .CK(clk), .Q(n40) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n237), .CK(clk), .Q(n41) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n238), .CK(clk), .Q(n42) );
  DFF_X1 \f_reg[0]  ( .D(n112), .CK(clk), .Q(f[0]), .QN(n212) );
  DFF_X1 \f_reg[1]  ( .D(n111), .CK(clk), .Q(f[1]), .QN(n213) );
  DFF_X1 \f_reg[2]  ( .D(n102), .CK(clk), .Q(f[2]), .QN(n214) );
  DFF_X1 \f_reg[7]  ( .D(n80), .CK(clk), .Q(f[7]), .QN(n215) );
  DFF_X1 \f_reg[8]  ( .D(n79), .CK(clk), .Q(f[8]), .QN(n216) );
  DFF_X1 \f_reg[9]  ( .D(n78), .CK(clk), .Q(f[9]), .QN(n217) );
  DFF_X1 \f_reg[10]  ( .D(n77), .CK(clk), .Q(n51), .QN(n218) );
  DFF_X1 \f_reg[11]  ( .D(n76), .CK(clk), .Q(n49), .QN(n219) );
  DFF_X1 \f_reg[12]  ( .D(n8), .CK(clk), .Q(n48), .QN(n220) );
  DFF_X1 \f_reg[13]  ( .D(n1), .CK(clk), .Q(n47), .QN(n221) );
  DFF_X1 \f_reg[14]  ( .D(n75), .CK(clk), .Q(n46), .QN(n222) );
  DFF_X1 \f_reg[15]  ( .D(n9), .CK(clk), .Q(f[15]), .QN(n72) );
  DFF_X1 \data_out_reg[15]  ( .D(n114), .CK(clk), .Q(data_out[15]), .QN(n195)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n165), .CK(clk), .Q(data_out[14]), .QN(n194)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n166), .CK(clk), .Q(data_out[13]), .QN(n193)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n167), .CK(clk), .Q(data_out[12]), .QN(n192)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n168), .CK(clk), .Q(data_out[11]), .QN(n191)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n169), .CK(clk), .Q(data_out[10]), .QN(n190)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n170), .CK(clk), .Q(data_out[9]), .QN(n189) );
  DFF_X1 \data_out_reg[8]  ( .D(n171), .CK(clk), .Q(data_out[8]), .QN(n188) );
  DFF_X1 \data_out_reg[7]  ( .D(n172), .CK(clk), .Q(data_out[7]), .QN(n187) );
  DFF_X1 \data_out_reg[6]  ( .D(n173), .CK(clk), .Q(data_out[6]), .QN(n186) );
  DFF_X1 \data_out_reg[5]  ( .D(n174), .CK(clk), .Q(data_out[5]), .QN(n185) );
  DFF_X1 \data_out_reg[4]  ( .D(n175), .CK(clk), .Q(data_out[4]), .QN(n184) );
  DFF_X1 \data_out_reg[3]  ( .D(n176), .CK(clk), .Q(data_out[3]), .QN(n183) );
  DFF_X1 \data_out_reg[2]  ( .D(n177), .CK(clk), .Q(data_out[2]), .QN(n182) );
  DFF_X1 \data_out_reg[1]  ( .D(n178), .CK(clk), .Q(data_out[1]), .QN(n181) );
  DFF_X1 \data_out_reg[0]  ( .D(n179), .CK(clk), .Q(data_out[0]), .QN(n180) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_14_DW_mult_tc_1 mult_2021 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_14_DW01_add_2 add_2022 ( .A({
        n202, n201, n200, n199, n198, n197, n211, n210, n209, n208, n207, n206, 
        n205, n204, n203, n196}), .B({f[15], n46, n47, n48, n49, n51, f[9:0]}), 
        .CI(1'b0), .SUM(adder) );
  DFF_X1 \f_reg[3]  ( .D(n85), .CK(clk), .Q(f[3]), .QN(n64) );
  DFF_X1 \f_reg[4]  ( .D(n83), .CK(clk), .Q(f[4]), .QN(n65) );
  DFF_X1 \f_reg[5]  ( .D(n82), .CK(clk), .Q(f[5]), .QN(n66) );
  DFF_X1 \f_reg[6]  ( .D(n81), .CK(clk), .Q(f[6]), .QN(n67) );
  DFF_X2 delay_reg ( .D(n113), .CK(clk), .Q(n7), .QN(n239) );
  MUX2_X1 U3 ( .A(N42), .B(n27), .S(n7), .Z(n200) );
  NAND3_X1 U4 ( .A1(n4), .A2(n2), .A3(n5), .ZN(n1) );
  NAND2_X1 U5 ( .A1(data_out_b[13]), .A2(n22), .ZN(n2) );
  NAND2_X1 U6 ( .A1(adder[13]), .A2(n20), .ZN(n4) );
  NAND2_X1 U8 ( .A1(n62), .A2(n47), .ZN(n5) );
  AND2_X4 U9 ( .A1(n45), .A2(n23), .ZN(n20) );
  AND2_X1 U10 ( .A1(clear_acc_delay), .A2(n239), .ZN(n6) );
  NAND3_X1 U11 ( .A1(n11), .A2(n10), .A3(n12), .ZN(n8) );
  NAND3_X1 U12 ( .A1(n15), .A2(n14), .A3(n16), .ZN(n9) );
  MUX2_X2 U13 ( .A(n34), .B(N37), .S(n239), .Z(n210) );
  MUX2_X2 U14 ( .A(n26), .B(N43), .S(n239), .Z(n201) );
  NAND2_X1 U15 ( .A1(data_out_b[12]), .A2(n22), .ZN(n10) );
  NAND2_X1 U16 ( .A1(adder[12]), .A2(n20), .ZN(n11) );
  NAND2_X1 U17 ( .A1(n62), .A2(n48), .ZN(n12) );
  AND2_X1 U18 ( .A1(n19), .A2(n17), .ZN(n13) );
  NAND2_X1 U19 ( .A1(n18), .A2(n13), .ZN(n75) );
  MUX2_X1 U20 ( .A(n29), .B(N40), .S(n239), .Z(n198) );
  MUX2_X2 U21 ( .A(n28), .B(N41), .S(n239), .Z(n199) );
  NAND2_X1 U22 ( .A1(data_out_b[15]), .A2(n22), .ZN(n14) );
  NAND2_X1 U23 ( .A1(adder[15]), .A2(n20), .ZN(n15) );
  NAND2_X1 U24 ( .A1(n62), .A2(f[15]), .ZN(n16) );
  NAND2_X1 U25 ( .A1(data_out_b[14]), .A2(n22), .ZN(n17) );
  NAND2_X1 U26 ( .A1(adder[14]), .A2(n20), .ZN(n18) );
  NAND2_X1 U27 ( .A1(n62), .A2(n46), .ZN(n19) );
  INV_X1 U28 ( .A(n23), .ZN(n22) );
  NAND2_X1 U29 ( .A1(n113), .A2(n21), .ZN(n241) );
  INV_X1 U30 ( .A(n45), .ZN(n62) );
  INV_X1 U31 ( .A(clear_acc), .ZN(n23) );
  OAI22_X1 U32 ( .A1(n183), .A2(n241), .B1(n64), .B2(n240), .ZN(n176) );
  OAI22_X1 U33 ( .A1(n184), .A2(n241), .B1(n65), .B2(n240), .ZN(n175) );
  OAI22_X1 U34 ( .A1(n185), .A2(n241), .B1(n66), .B2(n240), .ZN(n174) );
  OAI22_X1 U35 ( .A1(n186), .A2(n241), .B1(n67), .B2(n240), .ZN(n173) );
  OAI22_X1 U36 ( .A1(n187), .A2(n241), .B1(n215), .B2(n240), .ZN(n172) );
  OAI22_X1 U37 ( .A1(n188), .A2(n241), .B1(n216), .B2(n240), .ZN(n171) );
  OAI22_X1 U38 ( .A1(n189), .A2(n241), .B1(n217), .B2(n240), .ZN(n170) );
  INV_X1 U39 ( .A(wr_en_y), .ZN(n21) );
  INV_X1 U40 ( .A(m_ready), .ZN(n24) );
  NAND2_X1 U41 ( .A1(m_valid), .A2(n24), .ZN(n43) );
  OAI21_X1 U42 ( .B1(sel[4]), .B2(n74), .A(n43), .ZN(n113) );
  MUX2_X1 U43 ( .A(n25), .B(N44), .S(n6), .Z(n223) );
  MUX2_X1 U44 ( .A(n25), .B(N44), .S(n239), .Z(n202) );
  MUX2_X1 U45 ( .A(n26), .B(N43), .S(n6), .Z(n224) );
  MUX2_X1 U46 ( .A(n27), .B(N42), .S(n6), .Z(n225) );
  MUX2_X1 U47 ( .A(n28), .B(N41), .S(n6), .Z(n226) );
  MUX2_X1 U48 ( .A(n29), .B(N40), .S(n6), .Z(n227) );
  MUX2_X1 U49 ( .A(n32), .B(N39), .S(n6), .Z(n228) );
  MUX2_X1 U50 ( .A(n32), .B(N39), .S(n239), .Z(n197) );
  MUX2_X1 U51 ( .A(n33), .B(N38), .S(n6), .Z(n229) );
  MUX2_X1 U52 ( .A(n33), .B(N38), .S(n239), .Z(n211) );
  MUX2_X1 U53 ( .A(n34), .B(N37), .S(n6), .Z(n230) );
  MUX2_X1 U54 ( .A(n35), .B(N36), .S(n6), .Z(n231) );
  MUX2_X1 U55 ( .A(n35), .B(N36), .S(n239), .Z(n209) );
  MUX2_X1 U56 ( .A(n36), .B(N35), .S(n6), .Z(n232) );
  MUX2_X1 U57 ( .A(n36), .B(N35), .S(n239), .Z(n208) );
  MUX2_X1 U58 ( .A(n37), .B(N34), .S(n6), .Z(n233) );
  MUX2_X1 U59 ( .A(n37), .B(N34), .S(n239), .Z(n207) );
  MUX2_X1 U60 ( .A(n38), .B(N33), .S(n6), .Z(n234) );
  MUX2_X1 U61 ( .A(n38), .B(N33), .S(n239), .Z(n206) );
  MUX2_X1 U62 ( .A(n39), .B(N32), .S(n6), .Z(n235) );
  MUX2_X1 U63 ( .A(n39), .B(N32), .S(n239), .Z(n205) );
  MUX2_X1 U64 ( .A(n40), .B(N31), .S(n6), .Z(n236) );
  MUX2_X1 U65 ( .A(n40), .B(N31), .S(n239), .Z(n204) );
  MUX2_X1 U66 ( .A(n41), .B(N30), .S(n6), .Z(n237) );
  MUX2_X1 U67 ( .A(n41), .B(N30), .S(n239), .Z(n203) );
  MUX2_X1 U68 ( .A(n42), .B(N29), .S(n6), .Z(n238) );
  MUX2_X1 U69 ( .A(n42), .B(N29), .S(n239), .Z(n196) );
  INV_X1 U70 ( .A(n43), .ZN(n44) );
  OAI21_X1 U71 ( .B1(n44), .B2(n7), .A(n23), .ZN(n45) );
  AOI222_X1 U72 ( .A1(data_out_b[11]), .A2(n22), .B1(adder[11]), .B2(n20), 
        .C1(n62), .C2(n49), .ZN(n50) );
  INV_X1 U73 ( .A(n50), .ZN(n76) );
  AOI222_X1 U74 ( .A1(data_out_b[10]), .A2(n22), .B1(adder[10]), .B2(n20), 
        .C1(n62), .C2(n51), .ZN(n52) );
  INV_X1 U75 ( .A(n52), .ZN(n77) );
  AOI222_X1 U76 ( .A1(data_out_b[8]), .A2(n22), .B1(adder[8]), .B2(n20), .C1(
        n62), .C2(f[8]), .ZN(n53) );
  INV_X1 U77 ( .A(n53), .ZN(n79) );
  AOI222_X1 U78 ( .A1(data_out_b[7]), .A2(n22), .B1(adder[7]), .B2(n20), .C1(
        n62), .C2(f[7]), .ZN(n54) );
  INV_X1 U79 ( .A(n54), .ZN(n80) );
  AOI222_X1 U80 ( .A1(data_out_b[6]), .A2(n22), .B1(adder[6]), .B2(n20), .C1(
        n62), .C2(f[6]), .ZN(n55) );
  INV_X1 U81 ( .A(n55), .ZN(n81) );
  AOI222_X1 U82 ( .A1(data_out_b[5]), .A2(n22), .B1(adder[5]), .B2(n20), .C1(
        n62), .C2(f[5]), .ZN(n56) );
  INV_X1 U83 ( .A(n56), .ZN(n82) );
  AOI222_X1 U84 ( .A1(data_out_b[4]), .A2(n22), .B1(adder[4]), .B2(n20), .C1(
        n62), .C2(f[4]), .ZN(n57) );
  INV_X1 U85 ( .A(n57), .ZN(n83) );
  AOI222_X1 U86 ( .A1(data_out_b[3]), .A2(n22), .B1(adder[3]), .B2(n20), .C1(
        n62), .C2(f[3]), .ZN(n58) );
  INV_X1 U87 ( .A(n58), .ZN(n85) );
  AOI222_X1 U88 ( .A1(data_out_b[2]), .A2(n22), .B1(adder[2]), .B2(n20), .C1(
        n62), .C2(f[2]), .ZN(n59) );
  INV_X1 U89 ( .A(n59), .ZN(n102) );
  AOI222_X1 U90 ( .A1(data_out_b[1]), .A2(n22), .B1(adder[1]), .B2(n20), .C1(
        n62), .C2(f[1]), .ZN(n60) );
  INV_X1 U91 ( .A(n60), .ZN(n111) );
  AOI222_X1 U92 ( .A1(data_out_b[0]), .A2(n22), .B1(adder[0]), .B2(n20), .C1(
        n62), .C2(f[0]), .ZN(n61) );
  INV_X1 U93 ( .A(n61), .ZN(n112) );
  AOI222_X1 U94 ( .A1(data_out_b[9]), .A2(n22), .B1(adder[9]), .B2(n20), .C1(
        n62), .C2(f[9]), .ZN(n63) );
  INV_X1 U95 ( .A(n63), .ZN(n78) );
  NOR4_X1 U96 ( .A1(n49), .A2(n48), .A3(n47), .A4(n46), .ZN(n71) );
  NOR4_X1 U97 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n51), .ZN(n70) );
  NAND4_X1 U98 ( .A1(n67), .A2(n66), .A3(n65), .A4(n64), .ZN(n68) );
  NOR4_X1 U99 ( .A1(n68), .A2(f[0]), .A3(f[1]), .A4(f[2]), .ZN(n69) );
  NAND3_X1 U100 ( .A1(n71), .A2(n70), .A3(n69), .ZN(n73) );
  NAND3_X1 U101 ( .A1(wr_en_y), .A2(n73), .A3(n72), .ZN(n240) );
  OAI22_X1 U102 ( .A1(n180), .A2(n241), .B1(n212), .B2(n240), .ZN(n179) );
  OAI22_X1 U103 ( .A1(n181), .A2(n241), .B1(n213), .B2(n240), .ZN(n178) );
  OAI22_X1 U104 ( .A1(n182), .A2(n241), .B1(n214), .B2(n240), .ZN(n177) );
  OAI22_X1 U105 ( .A1(n190), .A2(n241), .B1(n218), .B2(n240), .ZN(n169) );
  OAI22_X1 U106 ( .A1(n191), .A2(n241), .B1(n219), .B2(n240), .ZN(n168) );
  OAI22_X1 U107 ( .A1(n192), .A2(n241), .B1(n220), .B2(n240), .ZN(n167) );
  OAI22_X1 U108 ( .A1(n193), .A2(n241), .B1(n221), .B2(n240), .ZN(n166) );
  OAI22_X1 U109 ( .A1(n194), .A2(n241), .B1(n222), .B2(n240), .ZN(n165) );
  OAI22_X1 U110 ( .A1(n195), .A2(n241), .B1(n72), .B2(n240), .ZN(n114) );
  AND4_X1 U111 ( .A1(sel[3]), .A2(sel[2]), .A3(sel[1]), .A4(sel[0]), .ZN(n74)
         );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_13_DW_mult_tc_1 ( a, b, 
        product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n9, n12, n13, n16, n18, n19, n21, n23, n25, n27, n29, n31,
         n32, n34, n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n50,
         n52, n53, n55, n56, n57, n58, n59, n62, n63, n64, n65, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n93, n95, n96, n97, n98, n99, n103,
         n104, n105, n106, n107, n111, n112, n113, n114, n115, n117, n119,
         n120, n122, n125, n127, n133, n135, n139, n141, n142, n143, n144,
         n145, n146, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n237, n239, n245, n247, n249, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n418, n419, n420, n421, n422, n423, n424, n426, n427, n428,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U148 ( .A(n265), .B(n144), .Z(n145) );
  XOR2_X1 U152 ( .A(n301), .B(n148), .Z(n149) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U161 ( .A(n177), .B(n168), .CI(n166), .CO(n163), .S(n164) );
  FA_X1 U162 ( .A(n170), .B(n172), .CI(n179), .CO(n165), .S(n166) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n263), .CI(n291), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n317), .B(n252), .CO(n173), .S(n174) );
  FA_X1 U167 ( .A(n180), .B(n187), .CI(n178), .CO(n175), .S(n176) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U169 ( .A(n193), .B(n282), .CI(n191), .CO(n179), .S(n180) );
  FA_X1 U170 ( .A(n268), .B(n292), .CI(n274), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U172 ( .A(n197), .B(n190), .CI(n188), .CO(n185), .S(n186) );
  FA_X1 U173 ( .A(n199), .B(n201), .CI(n192), .CO(n187), .S(n188) );
  FA_X1 U174 ( .A(n275), .B(n293), .CI(n194), .CO(n189), .S(n190) );
  FA_X1 U175 ( .A(n253), .B(n283), .CI(n305), .CO(n191), .S(n192) );
  HA_X1 U176 ( .A(n269), .B(n319), .CO(n193), .S(n194) );
  FA_X1 U177 ( .A(n205), .B(n200), .CI(n198), .CO(n195), .S(n196) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U179 ( .A(n284), .B(n294), .CI(n276), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n320), .B(n270), .CI(n306), .CO(n201), .S(n202) );
  FA_X1 U181 ( .A(n208), .B(n213), .CI(n206), .CO(n203), .S(n204) );
  FA_X1 U182 ( .A(n215), .B(n307), .CI(n210), .CO(n205), .S(n206) );
  FA_X1 U183 ( .A(n295), .B(n285), .CI(n254), .CO(n207), .S(n208) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U185 ( .A(n216), .B(n219), .CI(n214), .CO(n211), .S(n212) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n322), .B(n278), .CI(n308), .CO(n215), .S(n216) );
  FA_X1 U188 ( .A(n225), .B(n222), .CI(n220), .CO(n217), .S(n218) );
  FA_X1 U189 ( .A(n255), .B(n309), .CI(n297), .CO(n219), .S(n220) );
  HA_X1 U190 ( .A(n287), .B(n323), .CO(n221), .S(n222) );
  FA_X1 U191 ( .A(n229), .B(n298), .CI(n226), .CO(n223), .S(n224) );
  FA_X1 U192 ( .A(n324), .B(n288), .CI(n310), .CO(n225), .S(n226) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  HA_X1 U194 ( .A(n311), .B(n325), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n326), .B(n300), .CI(n312), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  XNOR2_X1 U414 ( .A(n550), .B(n490), .ZN(product[7]) );
  AND2_X1 U415 ( .A1(n526), .A2(n98), .ZN(n490) );
  OR2_X2 U416 ( .A1(n152), .A2(n163), .ZN(n557) );
  OR2_X1 U417 ( .A1(n224), .A2(n227), .ZN(n491) );
  OR2_X1 U418 ( .A1(n224), .A2(n227), .ZN(n563) );
  BUF_X2 U419 ( .A(n9), .Z(n562) );
  AND2_X1 U420 ( .A1(n232), .A2(n233), .ZN(n539) );
  BUF_X2 U421 ( .A(n570), .Z(n532) );
  INV_X1 U422 ( .A(n539), .ZN(n111) );
  OR2_X1 U423 ( .A1(n328), .A2(n314), .ZN(n492) );
  OR2_X1 U424 ( .A1(n329), .A2(n258), .ZN(n493) );
  CLKBUF_X3 U425 ( .A(n570), .Z(n522) );
  OR2_X2 U426 ( .A1(n217), .A2(n212), .ZN(n494) );
  OR2_X1 U427 ( .A1(n232), .A2(n233), .ZN(n495) );
  AND2_X1 U428 ( .A1(n224), .A2(n227), .ZN(n496) );
  CLKBUF_X1 U429 ( .A(n553), .Z(n497) );
  CLKBUF_X1 U430 ( .A(n86), .Z(n498) );
  INV_X1 U431 ( .A(n529), .ZN(n499) );
  INV_X1 U432 ( .A(n575), .ZN(n500) );
  NAND2_X1 U433 ( .A1(n555), .A2(n535), .ZN(n501) );
  NAND2_X1 U434 ( .A1(n555), .A2(n535), .ZN(n502) );
  NAND2_X1 U435 ( .A1(n555), .A2(n535), .ZN(n544) );
  BUF_X2 U436 ( .A(n9), .Z(n535) );
  INV_X1 U437 ( .A(n568), .ZN(n552) );
  INV_X1 U438 ( .A(n552), .ZN(n503) );
  INV_X1 U439 ( .A(n554), .ZN(n504) );
  XNOR2_X1 U440 ( .A(n574), .B(a[4]), .ZN(n556) );
  BUF_X2 U441 ( .A(n566), .Z(n505) );
  INV_X1 U442 ( .A(n576), .ZN(n506) );
  XOR2_X1 U443 ( .A(n568), .B(n249), .Z(n541) );
  INV_X1 U444 ( .A(n531), .ZN(n507) );
  BUF_X1 U445 ( .A(n570), .Z(n531) );
  BUF_X1 U446 ( .A(n534), .Z(n508) );
  AOI21_X1 U447 ( .B1(n96), .B2(n494), .A(n93), .ZN(n509) );
  XOR2_X1 U448 ( .A(n576), .B(a[6]), .Z(n540) );
  INV_X1 U449 ( .A(n239), .ZN(n510) );
  OR2_X2 U450 ( .A1(n511), .A2(n548), .ZN(n29) );
  XNOR2_X1 U451 ( .A(n577), .B(a[8]), .ZN(n511) );
  INV_X1 U452 ( .A(n548), .ZN(n27) );
  AOI21_X1 U453 ( .B1(n563), .B2(n104), .A(n496), .ZN(n512) );
  NOR2_X1 U454 ( .A1(n186), .A2(n195), .ZN(n513) );
  NOR2_X1 U455 ( .A1(n186), .A2(n195), .ZN(n82) );
  OR2_X2 U456 ( .A1(n541), .A2(n547), .ZN(n542) );
  XNOR2_X1 U457 ( .A(n149), .B(n514), .ZN(n144) );
  XNOR2_X1 U458 ( .A(n271), .B(n146), .ZN(n514) );
  OR2_X1 U459 ( .A1(n196), .A2(n203), .ZN(n515) );
  XNOR2_X1 U460 ( .A(n45), .B(n516), .ZN(product[12]) );
  AND2_X1 U461 ( .A1(n524), .A2(n79), .ZN(n516) );
  OAI21_X1 U462 ( .B1(n513), .B2(n86), .A(n83), .ZN(n517) );
  BUF_X2 U463 ( .A(n577), .Z(n518) );
  BUF_X2 U464 ( .A(n577), .Z(n519) );
  INV_X1 U465 ( .A(n578), .ZN(n577) );
  OAI21_X1 U466 ( .B1(n99), .B2(n97), .A(n98), .ZN(n520) );
  OAI21_X1 U467 ( .B1(n512), .B2(n97), .A(n98), .ZN(n96) );
  XNOR2_X2 U468 ( .A(n569), .B(a[4]), .ZN(n521) );
  INV_X1 U469 ( .A(n536), .ZN(n523) );
  OR2_X1 U470 ( .A1(n176), .A2(n185), .ZN(n524) );
  CLKBUF_X1 U471 ( .A(n18), .Z(n525) );
  OR2_X1 U472 ( .A1(n218), .A2(n223), .ZN(n526) );
  OR2_X2 U473 ( .A1(n540), .A2(n554), .ZN(n527) );
  OR2_X1 U474 ( .A1(n540), .A2(n554), .ZN(n23) );
  NOR2_X1 U475 ( .A1(n196), .A2(n203), .ZN(n85) );
  XNOR2_X1 U476 ( .A(n571), .B(a[2]), .ZN(n555) );
  INV_X1 U477 ( .A(n580), .ZN(n528) );
  INV_X1 U478 ( .A(n580), .ZN(n529) );
  OR2_X1 U479 ( .A1(n204), .A2(n211), .ZN(n530) );
  INV_X1 U480 ( .A(n571), .ZN(n570) );
  INV_X1 U481 ( .A(n576), .ZN(n575) );
  CLKBUF_X1 U482 ( .A(n104), .Z(n533) );
  OAI21_X1 U483 ( .B1(n546), .B2(n89), .A(n90), .ZN(n88) );
  NOR2_X1 U484 ( .A1(n164), .A2(n175), .ZN(n534) );
  INV_X1 U485 ( .A(n574), .ZN(n536) );
  CLKBUF_X1 U486 ( .A(n532), .Z(n537) );
  INV_X1 U487 ( .A(n239), .ZN(n538) );
  XOR2_X1 U488 ( .A(n578), .B(a[10]), .Z(n32) );
  INV_X1 U489 ( .A(n554), .ZN(n21) );
  OR2_X1 U490 ( .A1(n541), .A2(n547), .ZN(n6) );
  OR2_X2 U491 ( .A1(n541), .A2(n547), .ZN(n543) );
  NAND2_X1 U492 ( .A1(n555), .A2(n535), .ZN(n12) );
  XNOR2_X1 U493 ( .A(n1), .B(a[2]), .ZN(n9) );
  INV_X1 U494 ( .A(n249), .ZN(n566) );
  OAI21_X1 U495 ( .B1(n91), .B2(n89), .A(n90), .ZN(n545) );
  AOI21_X1 U496 ( .B1(n520), .B2(n494), .A(n93), .ZN(n546) );
  INV_X1 U497 ( .A(n566), .ZN(n547) );
  XNOR2_X1 U498 ( .A(n576), .B(a[8]), .ZN(n548) );
  XNOR2_X1 U499 ( .A(n88), .B(n549), .ZN(product[10]) );
  NAND2_X1 U500 ( .A1(n515), .A2(n86), .ZN(n549) );
  INV_X1 U501 ( .A(n571), .ZN(n569) );
  CLKBUF_X1 U502 ( .A(n512), .Z(n550) );
  INV_X1 U503 ( .A(n568), .ZN(n551) );
  AOI21_X1 U504 ( .B1(n545), .B2(n80), .A(n517), .ZN(n553) );
  XNOR2_X1 U505 ( .A(n574), .B(a[6]), .ZN(n554) );
  OAI21_X1 U506 ( .B1(n113), .B2(n115), .A(n114), .ZN(n112) );
  NOR2_X1 U507 ( .A1(n164), .A2(n175), .ZN(n75) );
  NAND2_X2 U508 ( .A1(n556), .A2(n16), .ZN(n18) );
  NAND2_X1 U509 ( .A1(n557), .A2(n69), .ZN(n47) );
  INV_X1 U510 ( .A(n73), .ZN(n71) );
  AOI21_X1 U511 ( .B1(n74), .B2(n557), .A(n67), .ZN(n65) );
  INV_X1 U512 ( .A(n69), .ZN(n67) );
  INV_X1 U513 ( .A(n74), .ZN(n72) );
  INV_X1 U514 ( .A(n95), .ZN(n93) );
  NAND2_X1 U515 ( .A1(n530), .A2(n90), .ZN(n52) );
  NAND2_X1 U516 ( .A1(n125), .A2(n76), .ZN(n48) );
  INV_X1 U517 ( .A(n508), .ZN(n125) );
  NAND2_X1 U518 ( .A1(n127), .A2(n83), .ZN(n50) );
  OAI21_X1 U519 ( .B1(n75), .B2(n79), .A(n76), .ZN(n74) );
  NOR2_X1 U520 ( .A1(n534), .A2(n78), .ZN(n73) );
  NAND2_X1 U521 ( .A1(n152), .A2(n163), .ZN(n69) );
  NAND2_X1 U522 ( .A1(n494), .A2(n95), .ZN(n53) );
  AOI21_X1 U523 ( .B1(n491), .B2(n104), .A(n496), .ZN(n99) );
  INV_X1 U524 ( .A(n113), .ZN(n135) );
  NAND2_X1 U525 ( .A1(n133), .A2(n106), .ZN(n56) );
  INV_X1 U526 ( .A(n105), .ZN(n133) );
  NOR2_X1 U527 ( .A1(n176), .A2(n185), .ZN(n78) );
  AOI21_X1 U528 ( .B1(n492), .B2(n120), .A(n117), .ZN(n115) );
  INV_X1 U529 ( .A(n119), .ZN(n117) );
  INV_X1 U530 ( .A(n122), .ZN(n120) );
  XNOR2_X1 U531 ( .A(n59), .B(n120), .ZN(product[2]) );
  NAND2_X1 U532 ( .A1(n492), .A2(n119), .ZN(n59) );
  NAND2_X1 U533 ( .A1(n176), .A2(n185), .ZN(n79) );
  NAND2_X1 U534 ( .A1(n164), .A2(n175), .ZN(n76) );
  NAND2_X1 U535 ( .A1(n196), .A2(n203), .ZN(n86) );
  NAND2_X1 U536 ( .A1(n212), .A2(n217), .ZN(n95) );
  NAND2_X1 U537 ( .A1(n204), .A2(n211), .ZN(n90) );
  XNOR2_X1 U538 ( .A(n57), .B(n112), .ZN(product[4]) );
  NAND2_X1 U539 ( .A1(n495), .A2(n111), .ZN(n57) );
  XNOR2_X1 U540 ( .A(n63), .B(n46), .ZN(product[15]) );
  NAND2_X1 U541 ( .A1(n558), .A2(n62), .ZN(n46) );
  NAND2_X1 U542 ( .A1(n73), .A2(n557), .ZN(n64) );
  NOR2_X1 U543 ( .A1(n234), .A2(n257), .ZN(n113) );
  OR2_X1 U544 ( .A1(n151), .A2(n139), .ZN(n558) );
  NOR2_X1 U545 ( .A1(n218), .A2(n223), .ZN(n97) );
  NAND2_X1 U546 ( .A1(n218), .A2(n223), .ZN(n98) );
  INV_X1 U547 ( .A(n37), .ZN(n237) );
  INV_X1 U548 ( .A(n41), .ZN(n235) );
  AND2_X1 U549 ( .A1(n493), .A2(n122), .ZN(product[1]) );
  XNOR2_X1 U550 ( .A(n528), .B(a[12]), .ZN(n37) );
  XNOR2_X1 U551 ( .A(n581), .B(a[14]), .ZN(n41) );
  OR2_X1 U552 ( .A1(n564), .A2(n507), .ZN(n392) );
  OAI22_X1 U553 ( .A1(n39), .A2(n336), .B1(n37), .B2(n335), .ZN(n263) );
  XOR2_X1 U554 ( .A(n579), .B(a[10]), .Z(n428) );
  OAI22_X1 U555 ( .A1(n543), .A2(n400), .B1(n399), .B2(n505), .ZN(n321) );
  XNOR2_X1 U556 ( .A(n518), .B(n564), .ZN(n352) );
  XNOR2_X1 U557 ( .A(n155), .B(n560), .ZN(n139) );
  XNOR2_X1 U558 ( .A(n153), .B(n141), .ZN(n560) );
  XNOR2_X1 U559 ( .A(n157), .B(n561), .ZN(n141) );
  XNOR2_X1 U560 ( .A(n145), .B(n143), .ZN(n561) );
  OAI22_X1 U561 ( .A1(n543), .A2(n408), .B1(n407), .B2(n505), .ZN(n329) );
  OAI22_X1 U562 ( .A1(n542), .A2(n406), .B1(n405), .B2(n505), .ZN(n327) );
  OAI22_X1 U563 ( .A1(n543), .A2(n402), .B1(n401), .B2(n505), .ZN(n323) );
  OAI22_X1 U564 ( .A1(n6), .A2(n404), .B1(n403), .B2(n505), .ZN(n325) );
  OAI22_X1 U565 ( .A1(n542), .A2(n398), .B1(n397), .B2(n505), .ZN(n319) );
  XNOR2_X1 U566 ( .A(n528), .B(n564), .ZN(n343) );
  AND2_X1 U567 ( .A1(n565), .A2(n235), .ZN(n260) );
  OAI22_X1 U568 ( .A1(n39), .A2(n335), .B1(n37), .B2(n334), .ZN(n262) );
  OAI22_X1 U569 ( .A1(n542), .A2(n395), .B1(n394), .B2(n505), .ZN(n316) );
  OAI22_X1 U570 ( .A1(n42), .A2(n583), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U571 ( .A1(n564), .A2(n583), .ZN(n332) );
  AND2_X1 U572 ( .A1(n565), .A2(n245), .ZN(n300) );
  OAI22_X1 U573 ( .A1(n543), .A2(n405), .B1(n404), .B2(n505), .ZN(n326) );
  XOR2_X1 U574 ( .A(n315), .B(n261), .Z(n150) );
  OAI22_X1 U575 ( .A1(n543), .A2(n394), .B1(n393), .B2(n505), .ZN(n315) );
  XNOR2_X1 U576 ( .A(n581), .B(n564), .ZN(n336) );
  NAND2_X1 U577 ( .A1(n427), .A2(n37), .ZN(n39) );
  XOR2_X1 U578 ( .A(n581), .B(a[12]), .Z(n427) );
  XNOR2_X1 U579 ( .A(n573), .B(n564), .ZN(n376) );
  AND2_X1 U580 ( .A1(n565), .A2(n237), .ZN(n264) );
  OAI22_X1 U581 ( .A1(n543), .A2(n397), .B1(n396), .B2(n505), .ZN(n318) );
  AND2_X1 U582 ( .A1(n565), .A2(n554), .ZN(n288) );
  OAI22_X1 U583 ( .A1(n6), .A2(n403), .B1(n402), .B2(n505), .ZN(n324) );
  AND2_X1 U584 ( .A1(n565), .A2(n239), .ZN(n270) );
  OAI22_X1 U585 ( .A1(n542), .A2(n399), .B1(n398), .B2(n505), .ZN(n320) );
  INV_X1 U586 ( .A(n19), .ZN(n576) );
  INV_X1 U587 ( .A(n25), .ZN(n578) );
  AND2_X1 U588 ( .A1(n565), .A2(n548), .ZN(n278) );
  OAI22_X1 U589 ( .A1(n542), .A2(n401), .B1(n400), .B2(n505), .ZN(n322) );
  NAND2_X1 U590 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U591 ( .A(n40), .B(a[14]), .Z(n426) );
  INV_X1 U592 ( .A(n7), .ZN(n571) );
  OAI22_X1 U593 ( .A1(n39), .A2(n582), .B1(n337), .B2(n37), .ZN(n252) );
  OAI22_X1 U594 ( .A1(n542), .A2(n396), .B1(n395), .B2(n505), .ZN(n317) );
  OR2_X1 U595 ( .A1(n564), .A2(n582), .ZN(n337) );
  AND2_X1 U596 ( .A1(n565), .A2(n247), .ZN(n314) );
  AND2_X1 U597 ( .A1(n565), .A2(n249), .ZN(product[0]) );
  OR2_X1 U598 ( .A1(n564), .A2(n523), .ZN(n377) );
  OR2_X1 U599 ( .A1(n564), .A2(n500), .ZN(n364) );
  OR2_X1 U600 ( .A1(n564), .A2(n578), .ZN(n353) );
  OR2_X1 U601 ( .A1(n564), .A2(n499), .ZN(n344) );
  OAI22_X1 U602 ( .A1(n39), .A2(n334), .B1(n37), .B2(n333), .ZN(n261) );
  XNOR2_X1 U603 ( .A(n581), .B(n422), .ZN(n333) );
  XNOR2_X1 U604 ( .A(n573), .B(b[11]), .ZN(n365) );
  XNOR2_X1 U605 ( .A(n581), .B(n424), .ZN(n335) );
  XNOR2_X1 U606 ( .A(n581), .B(n423), .ZN(n334) );
  OAI22_X1 U607 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U608 ( .A(n40), .B(n424), .ZN(n330) );
  XNOR2_X1 U609 ( .A(n40), .B(n564), .ZN(n331) );
  XNOR2_X1 U610 ( .A(n551), .B(b[11]), .ZN(n397) );
  XNOR2_X1 U611 ( .A(n552), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U612 ( .A(n551), .B(b[13]), .ZN(n395) );
  XNOR2_X1 U613 ( .A(n567), .B(b[14]), .ZN(n394) );
  XNOR2_X1 U614 ( .A(n518), .B(n418), .ZN(n345) );
  XNOR2_X1 U615 ( .A(n528), .B(n420), .ZN(n338) );
  XNOR2_X1 U616 ( .A(n537), .B(b[13]), .ZN(n378) );
  XNOR2_X1 U617 ( .A(n579), .B(n423), .ZN(n341) );
  XNOR2_X1 U618 ( .A(n529), .B(n424), .ZN(n342) );
  XNOR2_X1 U619 ( .A(n529), .B(n422), .ZN(n340) );
  XNOR2_X1 U620 ( .A(n579), .B(n421), .ZN(n339) );
  XNOR2_X1 U621 ( .A(n519), .B(n424), .ZN(n351) );
  XNOR2_X1 U622 ( .A(n522), .B(n418), .ZN(n384) );
  XNOR2_X1 U623 ( .A(n532), .B(n419), .ZN(n385) );
  XNOR2_X1 U624 ( .A(n522), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U625 ( .A(n532), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U626 ( .A(n532), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U627 ( .A(n522), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U628 ( .A(n537), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U629 ( .A(n573), .B(n418), .ZN(n369) );
  XNOR2_X1 U630 ( .A(n573), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U631 ( .A(n573), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U632 ( .A(n573), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U633 ( .A(n519), .B(n422), .ZN(n349) );
  XNOR2_X1 U634 ( .A(n518), .B(n423), .ZN(n350) );
  XNOR2_X1 U635 ( .A(n518), .B(n420), .ZN(n347) );
  XNOR2_X1 U636 ( .A(n519), .B(n421), .ZN(n348) );
  XNOR2_X1 U637 ( .A(n519), .B(n419), .ZN(n346) );
  XNOR2_X1 U638 ( .A(n551), .B(b[15]), .ZN(n393) );
  BUF_X1 U639 ( .A(n43), .Z(n565) );
  OAI22_X1 U640 ( .A1(n34), .A2(n339), .B1(n338), .B2(n510), .ZN(n265) );
  OAI22_X1 U641 ( .A1(n34), .A2(n340), .B1(n339), .B2(n510), .ZN(n266) );
  OAI22_X1 U642 ( .A1(n34), .A2(n341), .B1(n340), .B2(n510), .ZN(n267) );
  OAI22_X1 U643 ( .A1(n34), .A2(n342), .B1(n341), .B2(n510), .ZN(n268) );
  OAI22_X1 U644 ( .A1(n34), .A2(n343), .B1(n342), .B2(n538), .ZN(n269) );
  OAI22_X1 U645 ( .A1(n34), .A2(n499), .B1(n344), .B2(n538), .ZN(n253) );
  INV_X1 U646 ( .A(n32), .ZN(n239) );
  NAND2_X1 U647 ( .A1(n428), .A2(n32), .ZN(n34) );
  XNOR2_X1 U648 ( .A(n569), .B(a[4]), .ZN(n16) );
  AOI21_X1 U649 ( .B1(n495), .B2(n112), .A(n539), .ZN(n107) );
  XNOR2_X1 U650 ( .A(n84), .B(n50), .ZN(product[11]) );
  NAND2_X1 U651 ( .A1(n135), .A2(n114), .ZN(n58) );
  NAND2_X1 U652 ( .A1(n228), .A2(n231), .ZN(n106) );
  NOR2_X1 U653 ( .A1(n228), .A2(n231), .ZN(n105) );
  INV_X1 U654 ( .A(n13), .ZN(n574) );
  INV_X1 U655 ( .A(n513), .ZN(n127) );
  NOR2_X1 U656 ( .A1(n85), .A2(n82), .ZN(n80) );
  OAI21_X1 U657 ( .B1(n82), .B2(n86), .A(n83), .ZN(n81) );
  NAND2_X1 U658 ( .A1(n186), .A2(n195), .ZN(n83) );
  NAND2_X1 U659 ( .A1(n328), .A2(n314), .ZN(n119) );
  OAI22_X1 U660 ( .A1(n542), .A2(n407), .B1(n406), .B2(n505), .ZN(n328) );
  NAND2_X1 U661 ( .A1(n224), .A2(n227), .ZN(n103) );
  XNOR2_X1 U662 ( .A(n77), .B(n48), .ZN(product[13]) );
  NOR2_X1 U663 ( .A1(n204), .A2(n211), .ZN(n89) );
  OAI22_X1 U664 ( .A1(n29), .A2(n350), .B1(n349), .B2(n27), .ZN(n275) );
  OAI22_X1 U665 ( .A1(n29), .A2(n346), .B1(n345), .B2(n27), .ZN(n271) );
  OAI22_X1 U666 ( .A1(n29), .A2(n347), .B1(n346), .B2(n27), .ZN(n272) );
  OAI22_X1 U667 ( .A1(n29), .A2(n348), .B1(n347), .B2(n27), .ZN(n273) );
  OAI22_X1 U668 ( .A1(n29), .A2(n349), .B1(n348), .B2(n27), .ZN(n274) );
  OAI22_X1 U669 ( .A1(n29), .A2(n578), .B1(n353), .B2(n27), .ZN(n254) );
  OAI22_X1 U670 ( .A1(n29), .A2(n351), .B1(n350), .B2(n27), .ZN(n276) );
  XNOR2_X1 U671 ( .A(n506), .B(n419), .ZN(n357) );
  OAI22_X1 U672 ( .A1(n29), .A2(n352), .B1(n351), .B2(n27), .ZN(n277) );
  XNOR2_X1 U673 ( .A(n506), .B(n418), .ZN(n356) );
  XNOR2_X1 U674 ( .A(n506), .B(n422), .ZN(n360) );
  XNOR2_X1 U675 ( .A(n506), .B(b[9]), .ZN(n354) );
  XNOR2_X1 U676 ( .A(n506), .B(b[8]), .ZN(n355) );
  XNOR2_X1 U677 ( .A(n506), .B(n423), .ZN(n361) );
  XNOR2_X1 U678 ( .A(n575), .B(n421), .ZN(n359) );
  XNOR2_X1 U679 ( .A(n575), .B(n420), .ZN(n358) );
  XNOR2_X1 U680 ( .A(n506), .B(n564), .ZN(n363) );
  XNOR2_X1 U681 ( .A(n575), .B(n424), .ZN(n362) );
  XNOR2_X1 U682 ( .A(n55), .B(n533), .ZN(product[6]) );
  INV_X1 U683 ( .A(n1), .ZN(n568) );
  NAND2_X1 U684 ( .A1(n151), .A2(n139), .ZN(n62) );
  OAI21_X1 U685 ( .B1(n87), .B2(n85), .A(n498), .ZN(n84) );
  NAND2_X1 U686 ( .A1(n491), .A2(n103), .ZN(n55) );
  OAI22_X1 U687 ( .A1(n543), .A2(n503), .B1(n409), .B2(n505), .ZN(n258) );
  OR2_X1 U688 ( .A1(n564), .A2(n503), .ZN(n409) );
  INV_X1 U689 ( .A(n568), .ZN(n567) );
  INV_X1 U690 ( .A(n545), .ZN(n87) );
  AOI21_X1 U691 ( .B1(n88), .B2(n80), .A(n81), .ZN(n45) );
  XNOR2_X1 U692 ( .A(n70), .B(n47), .ZN(product[14]) );
  OAI22_X1 U693 ( .A1(n527), .A2(n358), .B1(n357), .B2(n504), .ZN(n282) );
  OAI22_X1 U694 ( .A1(n527), .A2(n356), .B1(n355), .B2(n504), .ZN(n280) );
  OAI22_X1 U695 ( .A1(n527), .A2(n362), .B1(n361), .B2(n504), .ZN(n286) );
  OAI22_X1 U696 ( .A1(n527), .A2(n500), .B1(n364), .B2(n504), .ZN(n255) );
  OAI22_X1 U697 ( .A1(n527), .A2(n360), .B1(n359), .B2(n504), .ZN(n284) );
  OAI22_X1 U698 ( .A1(n527), .A2(n361), .B1(n360), .B2(n504), .ZN(n285) );
  OAI22_X1 U699 ( .A1(n527), .A2(n357), .B1(n356), .B2(n504), .ZN(n281) );
  OAI22_X1 U700 ( .A1(n23), .A2(n363), .B1(n362), .B2(n21), .ZN(n287) );
  OAI22_X1 U701 ( .A1(n527), .A2(n355), .B1(n354), .B2(n21), .ZN(n279) );
  XNOR2_X1 U702 ( .A(n536), .B(n421), .ZN(n372) );
  XNOR2_X1 U703 ( .A(n536), .B(n423), .ZN(n374) );
  XNOR2_X1 U704 ( .A(n536), .B(n424), .ZN(n375) );
  OAI22_X1 U705 ( .A1(n23), .A2(n359), .B1(n358), .B2(n21), .ZN(n283) );
  XNOR2_X1 U706 ( .A(n572), .B(n422), .ZN(n373) );
  XNOR2_X1 U707 ( .A(n572), .B(n419), .ZN(n370) );
  XNOR2_X1 U708 ( .A(n572), .B(n420), .ZN(n371) );
  XOR2_X1 U709 ( .A(n509), .B(n52), .Z(product[9]) );
  OAI22_X1 U710 ( .A1(n525), .A2(n370), .B1(n369), .B2(n521), .ZN(n293) );
  OAI22_X1 U711 ( .A1(n525), .A2(n367), .B1(n366), .B2(n521), .ZN(n290) );
  OAI22_X1 U712 ( .A1(n18), .A2(n372), .B1(n371), .B2(n521), .ZN(n295) );
  OAI22_X1 U713 ( .A1(n18), .A2(n368), .B1(n367), .B2(n521), .ZN(n291) );
  OAI22_X1 U714 ( .A1(n525), .A2(n375), .B1(n374), .B2(n521), .ZN(n298) );
  OAI22_X1 U715 ( .A1(n18), .A2(n369), .B1(n368), .B2(n521), .ZN(n292) );
  OAI22_X1 U716 ( .A1(n18), .A2(n371), .B1(n370), .B2(n521), .ZN(n294) );
  OAI22_X1 U717 ( .A1(n18), .A2(n373), .B1(n372), .B2(n521), .ZN(n296) );
  OAI22_X1 U718 ( .A1(n18), .A2(n523), .B1(n377), .B2(n521), .ZN(n256) );
  OAI22_X1 U719 ( .A1(n18), .A2(n376), .B1(n375), .B2(n521), .ZN(n299) );
  OAI22_X1 U720 ( .A1(n18), .A2(n374), .B1(n373), .B2(n521), .ZN(n297) );
  OAI22_X1 U721 ( .A1(n18), .A2(n366), .B1(n365), .B2(n521), .ZN(n289) );
  XNOR2_X1 U722 ( .A(n522), .B(n420), .ZN(n386) );
  INV_X1 U723 ( .A(n16), .ZN(n245) );
  XNOR2_X1 U724 ( .A(n522), .B(n564), .ZN(n391) );
  XNOR2_X1 U725 ( .A(n532), .B(n424), .ZN(n390) );
  XNOR2_X1 U726 ( .A(n532), .B(n423), .ZN(n389) );
  XNOR2_X1 U727 ( .A(n531), .B(n422), .ZN(n388) );
  XNOR2_X1 U728 ( .A(n531), .B(n421), .ZN(n387) );
  XNOR2_X1 U729 ( .A(n520), .B(n53), .ZN(product[8]) );
  AOI21_X1 U730 ( .B1(n96), .B2(n494), .A(n93), .ZN(n91) );
  OAI21_X1 U731 ( .B1(n64), .B2(n497), .A(n65), .ZN(n63) );
  OAI21_X1 U732 ( .B1(n45), .B2(n78), .A(n79), .ZN(n77) );
  OAI21_X1 U733 ( .B1(n553), .B2(n71), .A(n72), .ZN(n70) );
  XNOR2_X1 U734 ( .A(n552), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U735 ( .A(n567), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U736 ( .A(n552), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U737 ( .A(n551), .B(n418), .ZN(n401) );
  XNOR2_X1 U738 ( .A(n567), .B(n564), .ZN(n408) );
  XNOR2_X1 U739 ( .A(n552), .B(n422), .ZN(n405) );
  XNOR2_X1 U740 ( .A(n551), .B(n421), .ZN(n404) );
  XNOR2_X1 U741 ( .A(n567), .B(n419), .ZN(n402) );
  XNOR2_X1 U742 ( .A(n552), .B(n420), .ZN(n403) );
  XNOR2_X1 U743 ( .A(n567), .B(n424), .ZN(n407) );
  XNOR2_X1 U744 ( .A(n551), .B(n423), .ZN(n406) );
  OAI21_X1 U745 ( .B1(n105), .B2(n107), .A(n106), .ZN(n104) );
  XOR2_X1 U746 ( .A(n56), .B(n107), .Z(product[5]) );
  XOR2_X1 U747 ( .A(n58), .B(n115), .Z(product[3]) );
  NAND2_X1 U748 ( .A1(n329), .A2(n258), .ZN(n122) );
  OAI22_X1 U749 ( .A1(n501), .A2(n379), .B1(n378), .B2(n562), .ZN(n301) );
  OAI22_X1 U750 ( .A1(n544), .A2(n380), .B1(n379), .B2(n562), .ZN(n302) );
  OAI22_X1 U751 ( .A1(n544), .A2(n385), .B1(n384), .B2(n562), .ZN(n307) );
  OAI22_X1 U752 ( .A1(n501), .A2(n382), .B1(n381), .B2(n562), .ZN(n304) );
  OAI22_X1 U753 ( .A1(n502), .A2(n381), .B1(n380), .B2(n562), .ZN(n303) );
  NAND2_X1 U754 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U755 ( .A1(n383), .A2(n502), .B1(n382), .B2(n562), .ZN(n305) );
  OAI22_X1 U756 ( .A1(n544), .A2(n384), .B1(n383), .B2(n562), .ZN(n306) );
  OAI22_X1 U757 ( .A1(n501), .A2(n386), .B1(n385), .B2(n562), .ZN(n308) );
  OAI22_X1 U758 ( .A1(n544), .A2(n387), .B1(n386), .B2(n562), .ZN(n309) );
  OAI22_X1 U759 ( .A1(n502), .A2(n507), .B1(n392), .B2(n562), .ZN(n257) );
  OAI22_X1 U760 ( .A1(n389), .A2(n12), .B1(n388), .B2(n562), .ZN(n311) );
  OAI22_X1 U761 ( .A1(n12), .A2(n388), .B1(n387), .B2(n562), .ZN(n310) );
  OAI22_X1 U762 ( .A1(n390), .A2(n501), .B1(n389), .B2(n562), .ZN(n312) );
  INV_X1 U763 ( .A(n562), .ZN(n247) );
  OAI22_X1 U764 ( .A1(n502), .A2(n391), .B1(n390), .B2(n562), .ZN(n313) );
  BUF_X4 U765 ( .A(n43), .Z(n564) );
  INV_X1 U766 ( .A(n574), .ZN(n572) );
  INV_X1 U767 ( .A(n574), .ZN(n573) );
  INV_X1 U768 ( .A(n580), .ZN(n579) );
  INV_X1 U769 ( .A(n31), .ZN(n580) );
  INV_X1 U770 ( .A(n582), .ZN(n581) );
  INV_X1 U771 ( .A(n36), .ZN(n582) );
  INV_X1 U772 ( .A(n40), .ZN(n583) );
  XOR2_X1 U773 ( .A(n259), .B(n251), .Z(n148) );
  XOR2_X1 U774 ( .A(n289), .B(n279), .Z(n146) );
  XOR2_X1 U775 ( .A(n159), .B(n150), .Z(n142) );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_13_DW01_add_2 ( A, B, CI, 
        SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n18, n20, n22, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n44, n45, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n65, n67, n68, n69, n70,
         n71, n73, n75, n76, n77, n78, n79, n81, n83, n84, n86, n88, n91, n94,
         n95, n96, n98, n100, n157, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183;

  OR2_X2 U122 ( .A1(A[10]), .A2(B[10]), .ZN(n165) );
  NOR2_X1 U123 ( .A1(A[14]), .A2(B[14]), .ZN(n157) );
  NOR2_X1 U124 ( .A1(A[14]), .A2(B[14]), .ZN(n25) );
  OR2_X1 U125 ( .A1(n18), .A2(n180), .ZN(n2) );
  AND2_X1 U126 ( .A1(n175), .A2(n86), .ZN(SUM[0]) );
  CLKBUF_X1 U127 ( .A(n58), .Z(n159) );
  OR2_X2 U128 ( .A1(A[9]), .A2(B[9]), .ZN(n160) );
  AND2_X1 U129 ( .A1(A[9]), .A2(B[9]), .ZN(n161) );
  NOR2_X1 U130 ( .A1(n163), .A2(n57), .ZN(n162) );
  NOR2_X2 U131 ( .A1(A[8]), .A2(B[8]), .ZN(n163) );
  NOR2_X1 U132 ( .A1(A[8]), .A2(B[8]), .ZN(n54) );
  XNOR2_X1 U133 ( .A(n174), .B(n164), .ZN(SUM[13]) );
  AND2_X1 U134 ( .A1(n166), .A2(n29), .ZN(n164) );
  XNOR2_X1 U135 ( .A(n38), .B(n6), .ZN(SUM[11]) );
  OR2_X1 U136 ( .A1(A[13]), .A2(B[13]), .ZN(n166) );
  OAI21_X1 U137 ( .B1(n58), .B2(n54), .A(n55), .ZN(n167) );
  NOR2_X1 U138 ( .A1(A[12]), .A2(B[12]), .ZN(n168) );
  AOI21_X1 U139 ( .B1(n52), .B2(n60), .A(n167), .ZN(n169) );
  AOI21_X1 U140 ( .B1(n162), .B2(n60), .A(n167), .ZN(n170) );
  AOI21_X1 U141 ( .B1(n162), .B2(n60), .A(n53), .ZN(n51) );
  INV_X1 U142 ( .A(n166), .ZN(n171) );
  AOI21_X1 U143 ( .B1(n165), .B2(n161), .A(n183), .ZN(n172) );
  NOR2_X1 U144 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  OAI21_X1 U145 ( .B1(n39), .B2(n169), .A(n40), .ZN(n173) );
  AOI21_X1 U146 ( .B1(n173), .B2(n30), .A(n31), .ZN(n174) );
  AOI21_X1 U147 ( .B1(n173), .B2(n30), .A(n31), .ZN(n1) );
  NOR2_X1 U148 ( .A1(A[7]), .A2(B[7]), .ZN(n57) );
  OR2_X1 U149 ( .A1(A[0]), .A2(B[0]), .ZN(n175) );
  INV_X1 U150 ( .A(n170), .ZN(n50) );
  INV_X1 U151 ( .A(n38), .ZN(n37) );
  AOI21_X1 U152 ( .B1(n178), .B2(n76), .A(n73), .ZN(n71) );
  AOI21_X1 U153 ( .B1(n179), .B2(n84), .A(n81), .ZN(n79) );
  INV_X1 U154 ( .A(n83), .ZN(n81) );
  AOI21_X1 U155 ( .B1(n177), .B2(n68), .A(n65), .ZN(n63) );
  INV_X1 U156 ( .A(n67), .ZN(n65) );
  OR2_X1 U157 ( .A1(n157), .A2(n28), .ZN(n176) );
  OAI21_X1 U158 ( .B1(n79), .B2(n77), .A(n78), .ZN(n76) );
  AOI21_X1 U159 ( .B1(n50), .B2(n160), .A(n161), .ZN(n45) );
  NAND2_X1 U160 ( .A1(n94), .A2(n55), .ZN(n9) );
  INV_X1 U161 ( .A(n86), .ZN(n84) );
  OAI21_X1 U162 ( .B1(n59), .B2(n57), .A(n159), .ZN(n56) );
  NAND2_X1 U163 ( .A1(n160), .A2(n49), .ZN(n8) );
  NAND2_X1 U164 ( .A1(n95), .A2(n58), .ZN(n10) );
  INV_X1 U165 ( .A(n57), .ZN(n95) );
  NAND2_X1 U166 ( .A1(n100), .A2(n78), .ZN(n15) );
  INV_X1 U167 ( .A(n77), .ZN(n100) );
  NAND2_X1 U168 ( .A1(n98), .A2(n70), .ZN(n13) );
  INV_X1 U169 ( .A(n69), .ZN(n98) );
  NAND2_X1 U170 ( .A1(n177), .A2(n67), .ZN(n12) );
  NAND2_X1 U171 ( .A1(n178), .A2(n75), .ZN(n14) );
  NAND2_X1 U172 ( .A1(n179), .A2(n83), .ZN(n16) );
  NAND2_X1 U173 ( .A1(n96), .A2(n62), .ZN(n11) );
  INV_X1 U174 ( .A(n61), .ZN(n96) );
  NAND2_X1 U175 ( .A1(n91), .A2(n36), .ZN(n6) );
  XNOR2_X1 U176 ( .A(n50), .B(n8), .ZN(SUM[9]) );
  XOR2_X1 U177 ( .A(n59), .B(n10), .Z(SUM[7]) );
  XOR2_X1 U178 ( .A(n15), .B(n79), .Z(SUM[2]) );
  NOR2_X1 U179 ( .A1(A[12]), .A2(B[12]), .ZN(n32) );
  OR2_X1 U180 ( .A1(A[5]), .A2(B[5]), .ZN(n177) );
  OR2_X1 U181 ( .A1(A[3]), .A2(B[3]), .ZN(n178) );
  NOR2_X1 U182 ( .A1(A[2]), .A2(B[2]), .ZN(n77) );
  NAND2_X1 U183 ( .A1(n88), .A2(n26), .ZN(n3) );
  NAND2_X1 U184 ( .A1(n182), .A2(n33), .ZN(n5) );
  XOR2_X1 U185 ( .A(n45), .B(n7), .Z(SUM[10]) );
  OR2_X1 U186 ( .A1(A[1]), .A2(B[1]), .ZN(n179) );
  AND2_X1 U187 ( .A1(A[15]), .A2(B[15]), .ZN(n180) );
  NAND2_X1 U188 ( .A1(A[14]), .A2(B[14]), .ZN(n26) );
  XNOR2_X1 U189 ( .A(n56), .B(n9), .ZN(SUM[8]) );
  XNOR2_X1 U190 ( .A(n16), .B(n84), .ZN(SUM[1]) );
  NOR2_X1 U191 ( .A1(A[6]), .A2(B[6]), .ZN(n61) );
  NOR2_X1 U192 ( .A1(A[4]), .A2(B[4]), .ZN(n69) );
  NAND2_X1 U193 ( .A1(A[7]), .A2(B[7]), .ZN(n58) );
  NAND2_X1 U194 ( .A1(A[2]), .A2(B[2]), .ZN(n78) );
  NAND2_X1 U195 ( .A1(A[5]), .A2(B[5]), .ZN(n67) );
  NAND2_X1 U196 ( .A1(A[1]), .A2(B[1]), .ZN(n83) );
  NAND2_X1 U197 ( .A1(A[0]), .A2(B[0]), .ZN(n86) );
  NAND2_X1 U198 ( .A1(A[3]), .A2(B[3]), .ZN(n75) );
  NAND2_X1 U199 ( .A1(A[6]), .A2(B[6]), .ZN(n62) );
  NAND2_X1 U200 ( .A1(A[4]), .A2(B[4]), .ZN(n70) );
  XNOR2_X1 U201 ( .A(n12), .B(n68), .ZN(SUM[5]) );
  XOR2_X1 U202 ( .A(n13), .B(n71), .Z(SUM[4]) );
  XNOR2_X1 U203 ( .A(n14), .B(n76), .ZN(SUM[3]) );
  INV_X1 U204 ( .A(n91), .ZN(n181) );
  INV_X1 U205 ( .A(n35), .ZN(n91) );
  OR2_X1 U206 ( .A1(A[12]), .A2(B[12]), .ZN(n182) );
  INV_X1 U207 ( .A(n24), .ZN(n22) );
  INV_X1 U208 ( .A(n60), .ZN(n59) );
  OAI21_X1 U209 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  XOR2_X1 U210 ( .A(n11), .B(n63), .Z(SUM[6]) );
  INV_X1 U211 ( .A(n163), .ZN(n94) );
  NOR2_X1 U212 ( .A1(n163), .A2(n57), .ZN(n52) );
  OAI21_X1 U213 ( .B1(n163), .B2(n58), .A(n55), .ZN(n53) );
  NAND2_X1 U214 ( .A1(A[8]), .A2(B[8]), .ZN(n55) );
  INV_X1 U215 ( .A(n183), .ZN(n44) );
  NAND2_X1 U216 ( .A1(A[11]), .A2(B[11]), .ZN(n36) );
  NOR2_X1 U217 ( .A1(B[11]), .A2(A[11]), .ZN(n35) );
  NAND2_X1 U218 ( .A1(A[9]), .A2(B[9]), .ZN(n49) );
  NAND2_X1 U219 ( .A1(A[12]), .A2(B[12]), .ZN(n33) );
  AND2_X1 U220 ( .A1(A[10]), .A2(B[10]), .ZN(n183) );
  NAND2_X1 U221 ( .A1(A[13]), .A2(B[13]), .ZN(n29) );
  OAI21_X1 U222 ( .B1(n37), .B2(n181), .A(n36), .ZN(n34) );
  INV_X1 U223 ( .A(n75), .ZN(n73) );
  OAI21_X1 U224 ( .B1(n71), .B2(n69), .A(n70), .ZN(n68) );
  XNOR2_X1 U225 ( .A(n20), .B(n2), .ZN(SUM[15]) );
  INV_X1 U226 ( .A(n157), .ZN(n88) );
  OAI21_X1 U227 ( .B1(n25), .B2(n29), .A(n26), .ZN(n24) );
  OAI21_X1 U228 ( .B1(n39), .B2(n51), .A(n172), .ZN(n38) );
  AOI21_X1 U229 ( .B1(n165), .B2(n161), .A(n183), .ZN(n40) );
  NOR2_X1 U230 ( .A1(A[15]), .A2(B[15]), .ZN(n18) );
  NOR2_X1 U231 ( .A1(n168), .A2(n35), .ZN(n30) );
  OAI21_X1 U232 ( .B1(n32), .B2(n36), .A(n33), .ZN(n31) );
  NAND2_X1 U233 ( .A1(n165), .A2(n44), .ZN(n7) );
  NAND2_X1 U234 ( .A1(n165), .A2(n160), .ZN(n39) );
  XNOR2_X1 U235 ( .A(n34), .B(n5), .ZN(SUM[12]) );
  XNOR2_X1 U236 ( .A(n27), .B(n3), .ZN(SUM[14]) );
  OAI21_X1 U237 ( .B1(n176), .B2(n174), .A(n22), .ZN(n20) );
  OAI21_X1 U238 ( .B1(n1), .B2(n171), .A(n29), .ZN(n27) );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_13 ( clk, clear_acc, 
        data_out_x, data_out, data_out_w, data_out_b, wr_en_y, m_valid, 
        m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [4:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
         N39, N40, N41, N42, N43, N44, n1, n2, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n85, n102, n111, n112, n113, n114, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n24), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n226), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n227), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n228), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n229), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n230), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n231), .CK(clk), .Q(n34) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n232), .CK(clk), .Q(n35) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n233), .CK(clk), .Q(n36) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n234), .CK(clk), .Q(n37) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n235), .CK(clk), .Q(n38) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n236), .CK(clk), .Q(n39) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n237), .CK(clk), .Q(n40) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n238), .CK(clk), .Q(n41) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n239), .CK(clk), .Q(n42) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n240), .CK(clk), .Q(n43) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n241), .CK(clk), .Q(n44) );
  DFF_X1 \f_reg[0]  ( .D(n114), .CK(clk), .Q(f[0]), .QN(n215) );
  DFF_X1 \f_reg[1]  ( .D(n113), .CK(clk), .Q(f[1]), .QN(n216) );
  DFF_X1 \f_reg[2]  ( .D(n112), .CK(clk), .Q(f[2]), .QN(n217) );
  DFF_X1 \f_reg[7]  ( .D(n82), .CK(clk), .Q(f[7]), .QN(n218) );
  DFF_X1 \f_reg[8]  ( .D(n81), .CK(clk), .Q(f[8]), .QN(n219) );
  DFF_X1 \f_reg[9]  ( .D(n80), .CK(clk), .Q(f[9]), .QN(n220) );
  DFF_X1 \f_reg[10]  ( .D(n79), .CK(clk), .Q(n54), .QN(n221) );
  DFF_X1 \f_reg[11]  ( .D(n78), .CK(clk), .Q(n52), .QN(n222) );
  DFF_X1 \f_reg[12]  ( .D(n5), .CK(clk), .Q(n51), .QN(n223) );
  DFF_X1 \f_reg[14]  ( .D(n11), .CK(clk), .Q(n49), .QN(n225) );
  DFF_X1 \f_reg[15]  ( .D(n18), .CK(clk), .Q(f[15]), .QN(n75) );
  DFF_X1 \data_out_reg[15]  ( .D(n167), .CK(clk), .Q(data_out[15]), .QN(n198)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n168), .CK(clk), .Q(data_out[14]), .QN(n197)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n169), .CK(clk), .Q(data_out[13]), .QN(n196)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n170), .CK(clk), .Q(data_out[12]), .QN(n195)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n171), .CK(clk), .Q(data_out[11]), .QN(n194)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n172), .CK(clk), .Q(data_out[10]), .QN(n193)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n173), .CK(clk), .Q(data_out[9]), .QN(n192) );
  DFF_X1 \data_out_reg[8]  ( .D(n174), .CK(clk), .Q(data_out[8]), .QN(n191) );
  DFF_X1 \data_out_reg[7]  ( .D(n175), .CK(clk), .Q(data_out[7]), .QN(n190) );
  DFF_X1 \data_out_reg[6]  ( .D(n176), .CK(clk), .Q(data_out[6]), .QN(n189) );
  DFF_X1 \data_out_reg[5]  ( .D(n177), .CK(clk), .Q(data_out[5]), .QN(n188) );
  DFF_X1 \data_out_reg[4]  ( .D(n178), .CK(clk), .Q(data_out[4]), .QN(n187) );
  DFF_X1 \data_out_reg[3]  ( .D(n179), .CK(clk), .Q(data_out[3]), .QN(n186) );
  DFF_X1 \data_out_reg[2]  ( .D(n180), .CK(clk), .Q(data_out[2]), .QN(n185) );
  DFF_X1 \data_out_reg[1]  ( .D(n181), .CK(clk), .Q(data_out[1]), .QN(n184) );
  DFF_X1 \data_out_reg[0]  ( .D(n182), .CK(clk), .Q(data_out[0]), .QN(n183) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_13_DW_mult_tc_1 mult_2021 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_13_DW01_add_2 add_2022 ( .A({
        n205, n204, n203, n202, n201, n200, n214, n213, n212, n211, n210, n209, 
        n208, n207, n206, n199}), .B({f[15], n49, n50, n51, n52, n54, f[9:0]}), 
        .CI(1'b0), .SUM(adder) );
  DFF_X1 \f_reg[3]  ( .D(n111), .CK(clk), .Q(f[3]), .QN(n67) );
  DFF_X1 \f_reg[4]  ( .D(n102), .CK(clk), .Q(f[4]), .QN(n68) );
  DFF_X1 \f_reg[5]  ( .D(n85), .CK(clk), .Q(f[5]), .QN(n69) );
  DFF_X1 \f_reg[6]  ( .D(n83), .CK(clk), .Q(f[6]), .QN(n70) );
  DFF_X1 \f_reg[13]  ( .D(n6), .CK(clk), .Q(n50), .QN(n224) );
  DFF_X2 delay_reg ( .D(n166), .CK(clk), .Q(n46), .QN(n242) );
  MUX2_X1 U3 ( .A(N44), .B(n27), .S(n46), .Z(n205) );
  AND2_X1 U4 ( .A1(clear_acc_delay), .A2(n242), .ZN(n1) );
  INV_X1 U5 ( .A(n48), .ZN(n65) );
  AND2_X1 U6 ( .A1(n48), .A2(n25), .ZN(n22) );
  AND2_X1 U8 ( .A1(n21), .A2(n19), .ZN(n2) );
  CLKBUF_X1 U9 ( .A(N36), .Z(n4) );
  MUX2_X2 U10 ( .A(n33), .B(N40), .S(n242), .Z(n201) );
  MUX2_X2 U11 ( .A(n35), .B(N38), .S(n242), .Z(n214) );
  NAND3_X1 U12 ( .A1(n13), .A2(n12), .A3(n14), .ZN(n5) );
  MUX2_X2 U13 ( .A(n34), .B(N39), .S(n242), .Z(n200) );
  NAND3_X1 U14 ( .A1(n9), .A2(n8), .A3(n10), .ZN(n6) );
  MUX2_X2 U15 ( .A(n29), .B(N42), .S(n242), .Z(n203) );
  CLKBUF_X1 U16 ( .A(N43), .Z(n7) );
  NAND2_X1 U17 ( .A1(n20), .A2(n2), .ZN(n18) );
  NAND2_X1 U18 ( .A1(n65), .A2(f[15]), .ZN(n21) );
  MUX2_X2 U19 ( .A(n36), .B(N37), .S(n242), .Z(n213) );
  NAND2_X1 U20 ( .A1(data_out_b[13]), .A2(n24), .ZN(n8) );
  NAND2_X1 U21 ( .A1(adder[13]), .A2(n22), .ZN(n9) );
  NAND2_X1 U22 ( .A1(n65), .A2(n50), .ZN(n10) );
  NAND3_X1 U23 ( .A1(n16), .A2(n15), .A3(n17), .ZN(n11) );
  NAND2_X1 U24 ( .A1(data_out_b[12]), .A2(n24), .ZN(n12) );
  NAND2_X1 U25 ( .A1(adder[12]), .A2(n22), .ZN(n13) );
  NAND2_X1 U26 ( .A1(n65), .A2(n51), .ZN(n14) );
  NAND2_X1 U27 ( .A1(data_out_b[14]), .A2(n24), .ZN(n15) );
  NAND2_X1 U28 ( .A1(adder[14]), .A2(n22), .ZN(n16) );
  NAND2_X1 U29 ( .A1(n65), .A2(n49), .ZN(n17) );
  MUX2_X2 U30 ( .A(n32), .B(N41), .S(n242), .Z(n202) );
  MUX2_X2 U31 ( .A(n28), .B(N43), .S(n242), .Z(n204) );
  NAND2_X1 U32 ( .A1(data_out_b[15]), .A2(n24), .ZN(n19) );
  NAND2_X1 U33 ( .A1(adder[15]), .A2(n22), .ZN(n20) );
  INV_X1 U34 ( .A(n25), .ZN(n24) );
  NAND2_X1 U35 ( .A1(n166), .A2(n23), .ZN(n244) );
  INV_X1 U36 ( .A(clear_acc), .ZN(n25) );
  OAI22_X1 U37 ( .A1(n186), .A2(n244), .B1(n67), .B2(n243), .ZN(n179) );
  OAI22_X1 U38 ( .A1(n187), .A2(n244), .B1(n68), .B2(n243), .ZN(n178) );
  OAI22_X1 U39 ( .A1(n188), .A2(n244), .B1(n69), .B2(n243), .ZN(n177) );
  OAI22_X1 U40 ( .A1(n189), .A2(n244), .B1(n70), .B2(n243), .ZN(n176) );
  OAI22_X1 U41 ( .A1(n190), .A2(n244), .B1(n218), .B2(n243), .ZN(n175) );
  OAI22_X1 U42 ( .A1(n191), .A2(n244), .B1(n219), .B2(n243), .ZN(n174) );
  OAI22_X1 U43 ( .A1(n192), .A2(n244), .B1(n220), .B2(n243), .ZN(n173) );
  INV_X1 U44 ( .A(wr_en_y), .ZN(n23) );
  INV_X1 U45 ( .A(m_ready), .ZN(n26) );
  NAND2_X1 U46 ( .A1(m_valid), .A2(n26), .ZN(n45) );
  OAI21_X1 U47 ( .B1(sel[4]), .B2(n77), .A(n45), .ZN(n166) );
  MUX2_X1 U48 ( .A(n27), .B(N44), .S(n1), .Z(n226) );
  MUX2_X1 U49 ( .A(n28), .B(n7), .S(n1), .Z(n227) );
  MUX2_X1 U50 ( .A(n29), .B(N42), .S(n1), .Z(n228) );
  MUX2_X1 U51 ( .A(n32), .B(N41), .S(n1), .Z(n229) );
  MUX2_X1 U52 ( .A(n33), .B(N40), .S(n1), .Z(n230) );
  MUX2_X1 U53 ( .A(n34), .B(N39), .S(n1), .Z(n231) );
  MUX2_X1 U54 ( .A(n35), .B(N38), .S(n1), .Z(n232) );
  MUX2_X1 U55 ( .A(n36), .B(N37), .S(n1), .Z(n233) );
  MUX2_X1 U56 ( .A(n37), .B(n4), .S(n1), .Z(n234) );
  MUX2_X1 U57 ( .A(n37), .B(N36), .S(n242), .Z(n212) );
  MUX2_X1 U58 ( .A(n38), .B(N35), .S(n1), .Z(n235) );
  MUX2_X1 U59 ( .A(n38), .B(N35), .S(n242), .Z(n211) );
  MUX2_X1 U60 ( .A(n39), .B(N34), .S(n1), .Z(n236) );
  MUX2_X1 U61 ( .A(n39), .B(N34), .S(n242), .Z(n210) );
  MUX2_X1 U62 ( .A(n40), .B(N33), .S(n1), .Z(n237) );
  MUX2_X1 U63 ( .A(n40), .B(N33), .S(n242), .Z(n209) );
  MUX2_X1 U64 ( .A(n41), .B(N32), .S(n1), .Z(n238) );
  MUX2_X1 U65 ( .A(n41), .B(N32), .S(n242), .Z(n208) );
  MUX2_X1 U66 ( .A(n42), .B(N31), .S(n1), .Z(n239) );
  MUX2_X1 U67 ( .A(n42), .B(N31), .S(n242), .Z(n207) );
  MUX2_X1 U68 ( .A(n43), .B(N30), .S(n1), .Z(n240) );
  MUX2_X1 U69 ( .A(n43), .B(N30), .S(n242), .Z(n206) );
  MUX2_X1 U70 ( .A(n44), .B(N29), .S(n1), .Z(n241) );
  MUX2_X1 U71 ( .A(n44), .B(N29), .S(n242), .Z(n199) );
  INV_X1 U72 ( .A(n45), .ZN(n47) );
  OAI21_X1 U73 ( .B1(n47), .B2(n46), .A(n25), .ZN(n48) );
  AOI222_X1 U74 ( .A1(data_out_b[11]), .A2(n24), .B1(adder[11]), .B2(n22), 
        .C1(n65), .C2(n52), .ZN(n53) );
  INV_X1 U75 ( .A(n53), .ZN(n78) );
  AOI222_X1 U76 ( .A1(data_out_b[10]), .A2(n24), .B1(adder[10]), .B2(n22), 
        .C1(n65), .C2(n54), .ZN(n55) );
  INV_X1 U77 ( .A(n55), .ZN(n79) );
  AOI222_X1 U78 ( .A1(data_out_b[8]), .A2(n24), .B1(adder[8]), .B2(n22), .C1(
        n65), .C2(f[8]), .ZN(n56) );
  INV_X1 U79 ( .A(n56), .ZN(n81) );
  AOI222_X1 U80 ( .A1(data_out_b[7]), .A2(n24), .B1(adder[7]), .B2(n22), .C1(
        n65), .C2(f[7]), .ZN(n57) );
  INV_X1 U81 ( .A(n57), .ZN(n82) );
  AOI222_X1 U82 ( .A1(data_out_b[6]), .A2(n24), .B1(adder[6]), .B2(n22), .C1(
        n65), .C2(f[6]), .ZN(n58) );
  INV_X1 U83 ( .A(n58), .ZN(n83) );
  AOI222_X1 U84 ( .A1(data_out_b[5]), .A2(n24), .B1(adder[5]), .B2(n22), .C1(
        n65), .C2(f[5]), .ZN(n59) );
  INV_X1 U85 ( .A(n59), .ZN(n85) );
  AOI222_X1 U86 ( .A1(data_out_b[4]), .A2(n24), .B1(adder[4]), .B2(n22), .C1(
        n65), .C2(f[4]), .ZN(n60) );
  INV_X1 U87 ( .A(n60), .ZN(n102) );
  AOI222_X1 U88 ( .A1(data_out_b[3]), .A2(n24), .B1(adder[3]), .B2(n22), .C1(
        n65), .C2(f[3]), .ZN(n61) );
  INV_X1 U89 ( .A(n61), .ZN(n111) );
  AOI222_X1 U90 ( .A1(data_out_b[2]), .A2(n24), .B1(adder[2]), .B2(n22), .C1(
        n65), .C2(f[2]), .ZN(n62) );
  INV_X1 U91 ( .A(n62), .ZN(n112) );
  AOI222_X1 U92 ( .A1(data_out_b[1]), .A2(n24), .B1(adder[1]), .B2(n22), .C1(
        n65), .C2(f[1]), .ZN(n63) );
  INV_X1 U93 ( .A(n63), .ZN(n113) );
  AOI222_X1 U94 ( .A1(data_out_b[0]), .A2(n24), .B1(adder[0]), .B2(n22), .C1(
        n65), .C2(f[0]), .ZN(n64) );
  INV_X1 U95 ( .A(n64), .ZN(n114) );
  AOI222_X1 U96 ( .A1(data_out_b[9]), .A2(n24), .B1(adder[9]), .B2(n22), .C1(
        n65), .C2(f[9]), .ZN(n66) );
  INV_X1 U97 ( .A(n66), .ZN(n80) );
  NOR4_X1 U98 ( .A1(n52), .A2(n51), .A3(n50), .A4(n49), .ZN(n74) );
  NOR4_X1 U99 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n54), .ZN(n73) );
  NAND4_X1 U100 ( .A1(n70), .A2(n69), .A3(n68), .A4(n67), .ZN(n71) );
  NOR4_X1 U101 ( .A1(n71), .A2(f[0]), .A3(f[1]), .A4(f[2]), .ZN(n72) );
  NAND3_X1 U102 ( .A1(n74), .A2(n73), .A3(n72), .ZN(n76) );
  NAND3_X1 U103 ( .A1(wr_en_y), .A2(n76), .A3(n75), .ZN(n243) );
  OAI22_X1 U104 ( .A1(n183), .A2(n244), .B1(n215), .B2(n243), .ZN(n182) );
  OAI22_X1 U105 ( .A1(n184), .A2(n244), .B1(n216), .B2(n243), .ZN(n181) );
  OAI22_X1 U106 ( .A1(n185), .A2(n244), .B1(n217), .B2(n243), .ZN(n180) );
  OAI22_X1 U107 ( .A1(n193), .A2(n244), .B1(n221), .B2(n243), .ZN(n172) );
  OAI22_X1 U108 ( .A1(n194), .A2(n244), .B1(n222), .B2(n243), .ZN(n171) );
  OAI22_X1 U109 ( .A1(n195), .A2(n244), .B1(n223), .B2(n243), .ZN(n170) );
  OAI22_X1 U110 ( .A1(n196), .A2(n244), .B1(n224), .B2(n243), .ZN(n169) );
  OAI22_X1 U111 ( .A1(n197), .A2(n244), .B1(n225), .B2(n243), .ZN(n168) );
  OAI22_X1 U112 ( .A1(n198), .A2(n244), .B1(n75), .B2(n243), .ZN(n167) );
  AND4_X1 U113 ( .A1(sel[3]), .A2(sel[2]), .A3(sel[1]), .A4(sel[0]), .ZN(n77)
         );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_12_DW_mult_tc_1 ( a, b, 
        product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n9, n12, n13, n16, n18, n19, n21, n25, n27, n29, n31, n32,
         n34, n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n50, n53,
         n55, n56, n57, n58, n59, n62, n63, n64, n65, n67, n69, n70, n72, n73,
         n74, n75, n76, n77, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n93, n95, n96, n97, n98, n99, n103, n104, n105, n106,
         n107, n109, n111, n112, n113, n114, n115, n117, n119, n120, n122,
         n127, n131, n133, n135, n139, n141, n142, n143, n144, n145, n147,
         n148, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n237,
         n239, n245, n247, n249, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n418, n419,
         n420, n421, n422, n423, n424, n426, n427, n428, n431, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U148 ( .A(n265), .B(n144), .Z(n145) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n272), .CI(n302), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n263), .CI(n291), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n317), .B(n252), .CO(n173), .S(n174) );
  FA_X1 U167 ( .A(n180), .B(n187), .CI(n178), .CO(n175), .S(n176) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U169 ( .A(n193), .B(n282), .CI(n191), .CO(n179), .S(n180) );
  FA_X1 U170 ( .A(n268), .B(n274), .CI(n292), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U172 ( .A(n197), .B(n190), .CI(n188), .CO(n185), .S(n186) );
  FA_X1 U173 ( .A(n199), .B(n201), .CI(n192), .CO(n187), .S(n188) );
  FA_X1 U174 ( .A(n275), .B(n293), .CI(n194), .CO(n189), .S(n190) );
  FA_X1 U175 ( .A(n305), .B(n253), .CI(n283), .CO(n191), .S(n192) );
  HA_X1 U176 ( .A(n319), .B(n269), .CO(n193), .S(n194) );
  FA_X1 U177 ( .A(n205), .B(n200), .CI(n198), .CO(n195), .S(n196) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U179 ( .A(n276), .B(n294), .CI(n284), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n320), .B(n270), .CI(n306), .CO(n201), .S(n202) );
  FA_X1 U182 ( .A(n215), .B(n307), .CI(n210), .CO(n205), .S(n206) );
  FA_X1 U183 ( .A(n295), .B(n254), .CI(n285), .CO(n207), .S(n208) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U185 ( .A(n216), .B(n219), .CI(n214), .CO(n211), .S(n212) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n322), .B(n278), .CI(n308), .CO(n215), .S(n216) );
  FA_X1 U188 ( .A(n225), .B(n222), .CI(n220), .CO(n217), .S(n218) );
  FA_X1 U189 ( .A(n297), .B(n309), .CI(n255), .CO(n219), .S(n220) );
  HA_X1 U190 ( .A(n323), .B(n287), .CO(n221), .S(n222) );
  FA_X1 U191 ( .A(n229), .B(n298), .CI(n226), .CO(n223), .S(n224) );
  FA_X1 U192 ( .A(n324), .B(n288), .CI(n310), .CO(n225), .S(n226) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  HA_X1 U194 ( .A(n325), .B(n311), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n326), .B(n300), .CI(n312), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  XNOR2_X1 U414 ( .A(n549), .B(n490), .ZN(product[7]) );
  AND2_X1 U415 ( .A1(n131), .A2(n98), .ZN(n490) );
  BUF_X2 U416 ( .A(n16), .Z(n584) );
  NOR2_X1 U417 ( .A1(n228), .A2(n231), .ZN(n105) );
  OR2_X1 U418 ( .A1(n164), .A2(n175), .ZN(n491) );
  OR2_X1 U419 ( .A1(n329), .A2(n258), .ZN(n492) );
  OR2_X1 U420 ( .A1(n176), .A2(n185), .ZN(n493) );
  CLKBUF_X1 U421 ( .A(n86), .Z(n494) );
  NOR2_X1 U422 ( .A1(n218), .A2(n223), .ZN(n495) );
  NOR2_X1 U423 ( .A1(n218), .A2(n223), .ZN(n97) );
  OR2_X1 U424 ( .A1(n196), .A2(n203), .ZN(n496) );
  OR2_X1 U425 ( .A1(n224), .A2(n227), .ZN(n497) );
  AND2_X1 U426 ( .A1(n224), .A2(n227), .ZN(n498) );
  XNOR2_X1 U427 ( .A(n603), .B(a[10]), .ZN(n428) );
  CLKBUF_X1 U428 ( .A(n558), .Z(n499) );
  BUF_X2 U429 ( .A(n9), .Z(n500) );
  XOR2_X1 U430 ( .A(n602), .B(a[10]), .Z(n501) );
  NAND2_X1 U431 ( .A1(n583), .A2(n431), .ZN(n502) );
  NAND2_X1 U432 ( .A1(n431), .A2(n583), .ZN(n520) );
  OR2_X1 U433 ( .A1(n554), .A2(n572), .ZN(n503) );
  OR2_X2 U434 ( .A1(n554), .A2(n572), .ZN(n504) );
  OR2_X1 U435 ( .A1(n554), .A2(n572), .ZN(n552) );
  XNOR2_X1 U436 ( .A(n505), .B(n147), .ZN(n144) );
  XNOR2_X1 U437 ( .A(n301), .B(n148), .ZN(n505) );
  XOR2_X1 U438 ( .A(n535), .B(n419), .Z(n385) );
  OR2_X1 U439 ( .A1(n75), .A2(n553), .ZN(n506) );
  BUF_X1 U440 ( .A(n37), .Z(n507) );
  INV_X2 U441 ( .A(n605), .ZN(n604) );
  INV_X1 U442 ( .A(n594), .ZN(n593) );
  XNOR2_X1 U443 ( .A(n508), .B(n166), .ZN(n164) );
  XNOR2_X1 U444 ( .A(n177), .B(n168), .ZN(n508) );
  XOR2_X1 U445 ( .A(n170), .B(n172), .Z(n509) );
  XOR2_X1 U446 ( .A(n509), .B(n179), .Z(n166) );
  NAND2_X1 U447 ( .A1(n170), .A2(n172), .ZN(n510) );
  NAND2_X1 U448 ( .A1(n170), .A2(n179), .ZN(n511) );
  NAND2_X1 U449 ( .A1(n172), .A2(n179), .ZN(n512) );
  NAND3_X1 U450 ( .A1(n510), .A2(n511), .A3(n512), .ZN(n165) );
  NAND2_X1 U451 ( .A1(n177), .A2(n168), .ZN(n513) );
  NAND2_X1 U452 ( .A1(n177), .A2(n166), .ZN(n514) );
  NAND2_X1 U453 ( .A1(n168), .A2(n166), .ZN(n515) );
  NAND3_X1 U454 ( .A1(n513), .A2(n514), .A3(n515), .ZN(n163) );
  XOR2_X1 U455 ( .A(n594), .B(a[4]), .Z(n16) );
  NAND2_X1 U456 ( .A1(n501), .A2(n32), .ZN(n516) );
  BUF_X1 U457 ( .A(n16), .Z(n583) );
  NAND2_X1 U458 ( .A1(n573), .A2(n527), .ZN(n558) );
  XNOR2_X1 U459 ( .A(n88), .B(n517), .ZN(product[10]) );
  NAND2_X1 U460 ( .A1(n496), .A2(n86), .ZN(n517) );
  XOR2_X1 U461 ( .A(n601), .B(a[8]), .Z(n559) );
  XNOR2_X1 U462 ( .A(n597), .B(a[6]), .ZN(n518) );
  XNOR2_X1 U463 ( .A(n91), .B(n519), .ZN(product[9]) );
  AND2_X1 U464 ( .A1(n560), .A2(n90), .ZN(n519) );
  BUF_X1 U465 ( .A(n599), .Z(n521) );
  BUF_X1 U466 ( .A(n597), .Z(n522) );
  BUF_X2 U467 ( .A(n9), .Z(n585) );
  CLKBUF_X1 U468 ( .A(n584), .Z(n523) );
  INV_X1 U469 ( .A(n589), .ZN(n524) );
  BUF_X2 U470 ( .A(n600), .Z(n525) );
  BUF_X2 U471 ( .A(n600), .Z(n526) );
  INV_X1 U472 ( .A(n601), .ZN(n600) );
  XOR2_X1 U473 ( .A(n591), .B(a[2]), .Z(n527) );
  AOI21_X1 U474 ( .B1(n577), .B2(n112), .A(n109), .ZN(n528) );
  INV_X1 U475 ( .A(n533), .ZN(n529) );
  XNOR2_X1 U476 ( .A(n522), .B(a[4]), .ZN(n431) );
  INV_X1 U477 ( .A(n597), .ZN(n595) );
  INV_X1 U478 ( .A(n544), .ZN(n530) );
  INV_X1 U479 ( .A(n544), .ZN(n590) );
  OR2_X2 U480 ( .A1(n562), .A2(n249), .ZN(n531) );
  OR2_X1 U481 ( .A1(n562), .A2(n249), .ZN(n6) );
  XNOR2_X1 U482 ( .A(n271), .B(n532), .ZN(n147) );
  XNOR2_X1 U483 ( .A(n289), .B(n279), .ZN(n532) );
  INV_X1 U484 ( .A(n521), .ZN(n533) );
  INV_X1 U485 ( .A(n526), .ZN(n534) );
  INV_X1 U486 ( .A(n592), .ZN(n535) );
  OAI21_X1 U487 ( .B1(n105), .B2(n107), .A(n106), .ZN(n536) );
  OR2_X1 U488 ( .A1(n559), .A2(n566), .ZN(n542) );
  INV_X1 U489 ( .A(n603), .ZN(n537) );
  INV_X1 U490 ( .A(n603), .ZN(n538) );
  CLKBUF_X1 U491 ( .A(n528), .Z(n539) );
  XOR2_X1 U492 ( .A(n591), .B(a[2]), .Z(n9) );
  NAND2_X1 U493 ( .A1(n431), .A2(n583), .ZN(n18) );
  INV_X1 U494 ( .A(n521), .ZN(n540) );
  INV_X1 U495 ( .A(n599), .ZN(n598) );
  XOR2_X1 U496 ( .A(n601), .B(a[10]), .Z(n541) );
  XOR2_X1 U497 ( .A(n601), .B(a[10]), .Z(n32) );
  INV_X1 U498 ( .A(n25), .ZN(n601) );
  CLKBUF_X1 U499 ( .A(n536), .Z(n543) );
  INV_X1 U500 ( .A(n1), .ZN(n544) );
  BUF_X2 U501 ( .A(n12), .Z(n557) );
  XOR2_X1 U502 ( .A(n208), .B(n213), .Z(n545) );
  XOR2_X1 U503 ( .A(n206), .B(n545), .Z(n204) );
  NAND2_X1 U504 ( .A1(n206), .A2(n208), .ZN(n546) );
  NAND2_X1 U505 ( .A1(n206), .A2(n213), .ZN(n547) );
  NAND2_X1 U506 ( .A1(n208), .A2(n213), .ZN(n548) );
  NAND3_X1 U507 ( .A1(n546), .A2(n547), .A3(n548), .ZN(n203) );
  CLKBUF_X1 U508 ( .A(n570), .Z(n549) );
  CLKBUF_X1 U509 ( .A(n571), .Z(n550) );
  CLKBUF_X1 U510 ( .A(n585), .Z(n551) );
  NOR2_X1 U511 ( .A1(n196), .A2(n203), .ZN(n85) );
  NOR2_X1 U512 ( .A1(n176), .A2(n185), .ZN(n553) );
  XNOR2_X1 U513 ( .A(n598), .B(a[6]), .ZN(n554) );
  OAI21_X1 U514 ( .B1(n99), .B2(n97), .A(n98), .ZN(n555) );
  OAI21_X1 U515 ( .B1(n495), .B2(n99), .A(n98), .ZN(n556) );
  OAI21_X1 U516 ( .B1(n570), .B2(n97), .A(n98), .ZN(n96) );
  NAND2_X1 U517 ( .A1(n573), .A2(n527), .ZN(n12) );
  OR2_X2 U518 ( .A1(n559), .A2(n566), .ZN(n29) );
  INV_X1 U519 ( .A(n566), .ZN(n27) );
  XNOR2_X1 U520 ( .A(n594), .B(a[2]), .ZN(n573) );
  OR2_X1 U521 ( .A1(n204), .A2(n211), .ZN(n560) );
  AOI21_X1 U522 ( .B1(n563), .B2(n80), .A(n81), .ZN(n571) );
  XNOR2_X1 U523 ( .A(n45), .B(n561), .ZN(product[12]) );
  AND2_X1 U524 ( .A1(n493), .A2(n79), .ZN(n561) );
  XOR2_X1 U525 ( .A(n591), .B(n249), .Z(n562) );
  INV_X1 U526 ( .A(n249), .ZN(n588) );
  OAI21_X1 U527 ( .B1(n91), .B2(n89), .A(n90), .ZN(n563) );
  AOI21_X1 U528 ( .B1(n96), .B2(n575), .A(n93), .ZN(n564) );
  OAI21_X1 U529 ( .B1(n564), .B2(n89), .A(n90), .ZN(n88) );
  NOR2_X1 U530 ( .A1(n164), .A2(n175), .ZN(n565) );
  NOR2_X1 U531 ( .A1(n164), .A2(n175), .ZN(n75) );
  INV_X1 U532 ( .A(n544), .ZN(n589) );
  INV_X1 U533 ( .A(n594), .ZN(n592) );
  XNOR2_X1 U534 ( .A(n599), .B(a[8]), .ZN(n566) );
  NOR2_X1 U535 ( .A1(n186), .A2(n195), .ZN(n567) );
  NOR2_X1 U536 ( .A1(n186), .A2(n195), .ZN(n82) );
  OR2_X1 U537 ( .A1(n542), .A2(n352), .ZN(n568) );
  OR2_X1 U538 ( .A1(n351), .A2(n27), .ZN(n569) );
  NAND2_X1 U539 ( .A1(n568), .A2(n569), .ZN(n277) );
  INV_X2 U540 ( .A(n518), .ZN(n21) );
  AOI21_X1 U541 ( .B1(n497), .B2(n104), .A(n498), .ZN(n570) );
  XNOR2_X1 U542 ( .A(n597), .B(a[6]), .ZN(n572) );
  BUF_X1 U543 ( .A(n43), .Z(n586) );
  NAND2_X1 U544 ( .A1(n574), .A2(n69), .ZN(n47) );
  NAND2_X1 U545 ( .A1(n73), .A2(n574), .ZN(n64) );
  INV_X1 U546 ( .A(n69), .ZN(n67) );
  INV_X1 U547 ( .A(n95), .ZN(n93) );
  AOI21_X1 U548 ( .B1(n563), .B2(n80), .A(n81), .ZN(n45) );
  NOR2_X1 U549 ( .A1(n567), .A2(n85), .ZN(n80) );
  NOR2_X1 U550 ( .A1(n75), .A2(n553), .ZN(n73) );
  XNOR2_X1 U551 ( .A(n77), .B(n48), .ZN(product[13]) );
  NAND2_X1 U552 ( .A1(n491), .A2(n76), .ZN(n48) );
  XNOR2_X1 U553 ( .A(n84), .B(n50), .ZN(product[11]) );
  NAND2_X1 U554 ( .A1(n127), .A2(n83), .ZN(n50) );
  OAI21_X1 U555 ( .B1(n87), .B2(n85), .A(n494), .ZN(n84) );
  INV_X1 U556 ( .A(n567), .ZN(n127) );
  OAI21_X1 U557 ( .B1(n565), .B2(n79), .A(n76), .ZN(n74) );
  OR2_X1 U558 ( .A1(n152), .A2(n163), .ZN(n574) );
  NAND2_X1 U559 ( .A1(n152), .A2(n163), .ZN(n69) );
  NAND2_X1 U560 ( .A1(n575), .A2(n95), .ZN(n53) );
  OAI21_X1 U561 ( .B1(n113), .B2(n115), .A(n114), .ZN(n112) );
  INV_X1 U562 ( .A(n495), .ZN(n131) );
  AOI21_X1 U563 ( .B1(n577), .B2(n112), .A(n109), .ZN(n107) );
  INV_X1 U564 ( .A(n111), .ZN(n109) );
  NAND2_X1 U565 ( .A1(n577), .A2(n111), .ZN(n57) );
  INV_X1 U566 ( .A(n122), .ZN(n120) );
  NAND2_X1 U567 ( .A1(n176), .A2(n185), .ZN(n79) );
  NAND2_X1 U568 ( .A1(n164), .A2(n175), .ZN(n76) );
  NAND2_X1 U569 ( .A1(n196), .A2(n203), .ZN(n86) );
  NAND2_X1 U570 ( .A1(n186), .A2(n195), .ZN(n83) );
  NAND2_X1 U571 ( .A1(n212), .A2(n217), .ZN(n95) );
  OR2_X1 U572 ( .A1(n212), .A2(n217), .ZN(n575) );
  NAND2_X1 U573 ( .A1(n204), .A2(n211), .ZN(n90) );
  INV_X1 U574 ( .A(n113), .ZN(n135) );
  NAND2_X1 U575 ( .A1(n576), .A2(n62), .ZN(n46) );
  NAND2_X1 U576 ( .A1(n133), .A2(n106), .ZN(n56) );
  AOI21_X1 U577 ( .B1(n582), .B2(n120), .A(n117), .ZN(n115) );
  INV_X1 U578 ( .A(n119), .ZN(n117) );
  OR2_X1 U579 ( .A1(n151), .A2(n139), .ZN(n576) );
  XNOR2_X1 U580 ( .A(n59), .B(n120), .ZN(product[2]) );
  NAND2_X1 U581 ( .A1(n582), .A2(n119), .ZN(n59) );
  OR2_X1 U582 ( .A1(n232), .A2(n233), .ZN(n577) );
  NAND2_X1 U583 ( .A1(n218), .A2(n223), .ZN(n98) );
  INV_X1 U584 ( .A(n37), .ZN(n237) );
  NAND2_X1 U585 ( .A1(n228), .A2(n231), .ZN(n106) );
  INV_X1 U586 ( .A(n41), .ZN(n235) );
  OR2_X1 U587 ( .A1(n224), .A2(n227), .ZN(n578) );
  AND2_X1 U588 ( .A1(n492), .A2(n122), .ZN(product[1]) );
  XNOR2_X1 U589 ( .A(n602), .B(a[12]), .ZN(n37) );
  XNOR2_X1 U590 ( .A(n604), .B(a[14]), .ZN(n41) );
  OR2_X1 U591 ( .A1(n586), .A2(n535), .ZN(n392) );
  XNOR2_X1 U592 ( .A(n593), .B(n586), .ZN(n391) );
  XNOR2_X1 U593 ( .A(n537), .B(n586), .ZN(n343) );
  AND2_X1 U594 ( .A1(n587), .A2(n572), .ZN(n288) );
  XNOR2_X1 U595 ( .A(n525), .B(n586), .ZN(n352) );
  OAI22_X1 U596 ( .A1(n42), .A2(n607), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U597 ( .A1(n586), .A2(n607), .ZN(n332) );
  XOR2_X1 U598 ( .A(n315), .B(n261), .Z(n150) );
  XNOR2_X1 U599 ( .A(n155), .B(n580), .ZN(n139) );
  XNOR2_X1 U600 ( .A(n153), .B(n141), .ZN(n580) );
  XNOR2_X1 U601 ( .A(n157), .B(n581), .ZN(n141) );
  XNOR2_X1 U602 ( .A(n145), .B(n143), .ZN(n581) );
  XNOR2_X1 U603 ( .A(n596), .B(n586), .ZN(n376) );
  XNOR2_X1 U604 ( .A(n604), .B(n586), .ZN(n336) );
  AND2_X1 U605 ( .A1(n587), .A2(n247), .ZN(n314) );
  NAND2_X1 U606 ( .A1(n427), .A2(n37), .ZN(n39) );
  XOR2_X1 U607 ( .A(n604), .B(a[12]), .Z(n427) );
  OR2_X1 U608 ( .A1(n328), .A2(n314), .ZN(n582) );
  AND2_X1 U609 ( .A1(n587), .A2(n566), .ZN(n278) );
  OAI22_X1 U610 ( .A1(n39), .A2(n336), .B1(n507), .B2(n335), .ZN(n263) );
  AND2_X1 U611 ( .A1(n587), .A2(n237), .ZN(n264) );
  AND2_X1 U612 ( .A1(n587), .A2(n245), .ZN(n300) );
  AND2_X1 U613 ( .A1(n587), .A2(n239), .ZN(n270) );
  AND2_X1 U614 ( .A1(n587), .A2(n235), .ZN(n260) );
  OAI22_X1 U615 ( .A1(n39), .A2(n335), .B1(n507), .B2(n334), .ZN(n262) );
  NAND2_X1 U616 ( .A1(n328), .A2(n314), .ZN(n119) );
  INV_X1 U617 ( .A(n19), .ZN(n599) );
  NAND2_X1 U618 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U619 ( .A(n606), .B(a[14]), .Z(n426) );
  OAI22_X1 U620 ( .A1(n39), .A2(n605), .B1(n337), .B2(n507), .ZN(n252) );
  OR2_X1 U621 ( .A1(n586), .A2(n605), .ZN(n337) );
  AND2_X1 U622 ( .A1(n587), .A2(n249), .ZN(product[0]) );
  OR2_X1 U623 ( .A1(n586), .A2(n529), .ZN(n364) );
  OR2_X1 U624 ( .A1(n586), .A2(n534), .ZN(n353) );
  OR2_X1 U625 ( .A1(n586), .A2(n603), .ZN(n344) );
  OR2_X1 U626 ( .A1(n586), .A2(n522), .ZN(n377) );
  OAI22_X1 U627 ( .A1(n39), .A2(n334), .B1(n507), .B2(n333), .ZN(n261) );
  XNOR2_X1 U628 ( .A(n604), .B(n422), .ZN(n333) );
  XNOR2_X1 U629 ( .A(n596), .B(b[11]), .ZN(n365) );
  XNOR2_X1 U630 ( .A(n604), .B(n424), .ZN(n335) );
  XNOR2_X1 U631 ( .A(n604), .B(n423), .ZN(n334) );
  OAI22_X1 U632 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U633 ( .A(n606), .B(n424), .ZN(n330) );
  XNOR2_X1 U634 ( .A(n606), .B(n586), .ZN(n331) );
  XNOR2_X1 U635 ( .A(n525), .B(n418), .ZN(n345) );
  XNOR2_X1 U636 ( .A(n537), .B(n420), .ZN(n338) );
  XNOR2_X1 U637 ( .A(n592), .B(b[13]), .ZN(n378) );
  XNOR2_X1 U638 ( .A(n538), .B(n424), .ZN(n342) );
  XNOR2_X1 U639 ( .A(n593), .B(n424), .ZN(n390) );
  XNOR2_X1 U640 ( .A(n525), .B(n424), .ZN(n351) );
  XNOR2_X1 U641 ( .A(n538), .B(n423), .ZN(n341) );
  XNOR2_X1 U642 ( .A(n537), .B(n422), .ZN(n340) );
  XNOR2_X1 U643 ( .A(n538), .B(n421), .ZN(n339) );
  XNOR2_X1 U644 ( .A(n592), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U645 ( .A(n592), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U646 ( .A(n593), .B(n418), .ZN(n384) );
  XNOR2_X1 U647 ( .A(n593), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U648 ( .A(n593), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U649 ( .A(n593), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U650 ( .A(n593), .B(n423), .ZN(n389) );
  XNOR2_X1 U651 ( .A(n592), .B(n422), .ZN(n388) );
  XNOR2_X1 U652 ( .A(n526), .B(n423), .ZN(n350) );
  XNOR2_X1 U653 ( .A(n526), .B(n422), .ZN(n349) );
  XNOR2_X1 U654 ( .A(n596), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U655 ( .A(n596), .B(n418), .ZN(n369) );
  XNOR2_X1 U656 ( .A(n596), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U657 ( .A(n596), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U658 ( .A(n530), .B(b[11]), .ZN(n397) );
  XNOR2_X1 U659 ( .A(n530), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U660 ( .A(n590), .B(b[13]), .ZN(n395) );
  XNOR2_X1 U661 ( .A(n530), .B(b[14]), .ZN(n394) );
  XNOR2_X1 U662 ( .A(n592), .B(n421), .ZN(n387) );
  XNOR2_X1 U663 ( .A(n525), .B(n421), .ZN(n348) );
  XNOR2_X1 U664 ( .A(n593), .B(n420), .ZN(n386) );
  XNOR2_X1 U665 ( .A(n525), .B(n420), .ZN(n347) );
  XNOR2_X1 U666 ( .A(n526), .B(n419), .ZN(n346) );
  XNOR2_X1 U667 ( .A(n590), .B(b[15]), .ZN(n393) );
  BUF_X1 U668 ( .A(n43), .Z(n587) );
  OAI22_X1 U669 ( .A1(n516), .A2(n339), .B1(n338), .B2(n541), .ZN(n265) );
  OAI22_X1 U670 ( .A1(n34), .A2(n340), .B1(n339), .B2(n541), .ZN(n266) );
  OAI22_X1 U671 ( .A1(n516), .A2(n341), .B1(n340), .B2(n541), .ZN(n267) );
  OAI22_X1 U672 ( .A1(n34), .A2(n342), .B1(n341), .B2(n541), .ZN(n268) );
  OAI22_X1 U673 ( .A1(n516), .A2(n343), .B1(n342), .B2(n541), .ZN(n269) );
  INV_X1 U674 ( .A(n32), .ZN(n239) );
  OAI22_X1 U675 ( .A1(n34), .A2(n603), .B1(n344), .B2(n541), .ZN(n253) );
  NAND2_X1 U676 ( .A1(n428), .A2(n32), .ZN(n34) );
  INV_X1 U677 ( .A(n13), .ZN(n597) );
  INV_X1 U678 ( .A(n105), .ZN(n133) );
  AOI21_X1 U679 ( .B1(n74), .B2(n574), .A(n67), .ZN(n65) );
  INV_X1 U680 ( .A(n74), .ZN(n72) );
  OAI22_X1 U681 ( .A1(n503), .A2(n362), .B1(n361), .B2(n21), .ZN(n286) );
  OAI22_X1 U682 ( .A1(n503), .A2(n358), .B1(n357), .B2(n21), .ZN(n282) );
  OAI22_X1 U683 ( .A1(n504), .A2(n356), .B1(n355), .B2(n21), .ZN(n280) );
  OAI22_X1 U684 ( .A1(n503), .A2(n360), .B1(n359), .B2(n21), .ZN(n284) );
  OAI22_X1 U685 ( .A1(n361), .A2(n503), .B1(n360), .B2(n21), .ZN(n285) );
  OAI22_X1 U686 ( .A1(n504), .A2(n529), .B1(n364), .B2(n21), .ZN(n255) );
  OAI22_X1 U687 ( .A1(n552), .A2(n363), .B1(n362), .B2(n21), .ZN(n287) );
  OAI22_X1 U688 ( .A1(n504), .A2(n357), .B1(n356), .B2(n21), .ZN(n281) );
  OAI22_X1 U689 ( .A1(n504), .A2(n355), .B1(n354), .B2(n21), .ZN(n279) );
  NAND2_X1 U690 ( .A1(n232), .A2(n233), .ZN(n111) );
  NAND2_X1 U691 ( .A1(n497), .A2(n103), .ZN(n55) );
  NAND2_X1 U692 ( .A1(n224), .A2(n227), .ZN(n103) );
  OAI22_X1 U693 ( .A1(n552), .A2(n359), .B1(n358), .B2(n21), .ZN(n283) );
  NOR2_X1 U694 ( .A1(n204), .A2(n211), .ZN(n89) );
  OAI22_X1 U695 ( .A1(n542), .A2(n346), .B1(n345), .B2(n27), .ZN(n271) );
  OAI22_X1 U696 ( .A1(n29), .A2(n347), .B1(n346), .B2(n27), .ZN(n272) );
  OAI22_X1 U697 ( .A1(n542), .A2(n350), .B1(n349), .B2(n27), .ZN(n275) );
  OAI22_X1 U698 ( .A1(n542), .A2(n351), .B1(n350), .B2(n27), .ZN(n276) );
  OAI22_X1 U699 ( .A1(n29), .A2(n348), .B1(n347), .B2(n27), .ZN(n273) );
  OAI22_X1 U700 ( .A1(n29), .A2(n349), .B1(n348), .B2(n27), .ZN(n274) );
  OAI22_X1 U701 ( .A1(n29), .A2(n534), .B1(n353), .B2(n27), .ZN(n254) );
  XNOR2_X1 U702 ( .A(n533), .B(n586), .ZN(n363) );
  XNOR2_X1 U703 ( .A(n540), .B(n419), .ZN(n357) );
  XNOR2_X1 U704 ( .A(n540), .B(n418), .ZN(n356) );
  XNOR2_X1 U705 ( .A(n540), .B(b[9]), .ZN(n354) );
  XNOR2_X1 U706 ( .A(n598), .B(n424), .ZN(n362) );
  XNOR2_X1 U707 ( .A(n540), .B(n422), .ZN(n360) );
  XNOR2_X1 U708 ( .A(n540), .B(n423), .ZN(n361) );
  XNOR2_X1 U709 ( .A(n540), .B(b[8]), .ZN(n355) );
  XNOR2_X1 U710 ( .A(n533), .B(n420), .ZN(n358) );
  XNOR2_X1 U711 ( .A(n533), .B(n421), .ZN(n359) );
  XNOR2_X1 U712 ( .A(n63), .B(n46), .ZN(product[15]) );
  INV_X1 U713 ( .A(n7), .ZN(n594) );
  NOR2_X1 U714 ( .A1(n234), .A2(n257), .ZN(n113) );
  NAND2_X1 U715 ( .A1(n135), .A2(n114), .ZN(n58) );
  XNOR2_X1 U716 ( .A(n595), .B(n424), .ZN(n375) );
  XNOR2_X1 U717 ( .A(n595), .B(n421), .ZN(n372) );
  XNOR2_X1 U718 ( .A(n595), .B(n419), .ZN(n370) );
  XNOR2_X1 U719 ( .A(n595), .B(n420), .ZN(n371) );
  XNOR2_X1 U720 ( .A(n595), .B(n423), .ZN(n374) );
  XNOR2_X1 U721 ( .A(n595), .B(n422), .ZN(n373) );
  INV_X1 U722 ( .A(n1), .ZN(n591) );
  OR2_X1 U723 ( .A1(n586), .A2(n544), .ZN(n409) );
  XNOR2_X1 U724 ( .A(n589), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U725 ( .A(n590), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U726 ( .A(n590), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U727 ( .A(n530), .B(n418), .ZN(n401) );
  XNOR2_X1 U728 ( .A(n530), .B(n586), .ZN(n408) );
  XNOR2_X1 U729 ( .A(n589), .B(n422), .ZN(n405) );
  XNOR2_X1 U730 ( .A(n590), .B(n420), .ZN(n403) );
  XNOR2_X1 U731 ( .A(n589), .B(n421), .ZN(n404) );
  XNOR2_X1 U732 ( .A(n589), .B(n419), .ZN(n402) );
  XNOR2_X1 U733 ( .A(n530), .B(n424), .ZN(n407) );
  XNOR2_X1 U734 ( .A(n530), .B(n423), .ZN(n406) );
  XNOR2_X1 U735 ( .A(n70), .B(n47), .ZN(product[14]) );
  OAI21_X1 U736 ( .B1(n82), .B2(n86), .A(n83), .ZN(n81) );
  OAI21_X1 U737 ( .B1(n105), .B2(n528), .A(n106), .ZN(n104) );
  AOI21_X1 U738 ( .B1(n536), .B2(n578), .A(n498), .ZN(n99) );
  XNOR2_X1 U739 ( .A(n55), .B(n543), .ZN(product[6]) );
  NAND2_X1 U740 ( .A1(n151), .A2(n139), .ZN(n62) );
  OAI22_X1 U741 ( .A1(n520), .A2(n370), .B1(n369), .B2(n584), .ZN(n293) );
  OAI22_X1 U742 ( .A1(n520), .A2(n367), .B1(n366), .B2(n523), .ZN(n290) );
  OAI22_X1 U743 ( .A1(n520), .A2(n375), .B1(n374), .B2(n523), .ZN(n298) );
  OAI22_X1 U744 ( .A1(n502), .A2(n368), .B1(n367), .B2(n584), .ZN(n291) );
  OAI22_X1 U745 ( .A1(n502), .A2(n369), .B1(n368), .B2(n584), .ZN(n292) );
  OAI22_X1 U746 ( .A1(n520), .A2(n373), .B1(n372), .B2(n584), .ZN(n296) );
  OAI22_X1 U747 ( .A1(n18), .A2(n372), .B1(n371), .B2(n584), .ZN(n295) );
  OAI22_X1 U748 ( .A1(n502), .A2(n374), .B1(n373), .B2(n584), .ZN(n297) );
  OAI22_X1 U749 ( .A1(n502), .A2(n522), .B1(n377), .B2(n584), .ZN(n256) );
  OAI22_X1 U750 ( .A1(n18), .A2(n371), .B1(n370), .B2(n584), .ZN(n294) );
  OAI22_X1 U751 ( .A1(n520), .A2(n376), .B1(n375), .B2(n584), .ZN(n299) );
  OAI22_X1 U752 ( .A1(n520), .A2(n366), .B1(n365), .B2(n584), .ZN(n289) );
  INV_X1 U753 ( .A(n584), .ZN(n245) );
  INV_X1 U754 ( .A(n88), .ZN(n87) );
  XOR2_X1 U755 ( .A(n56), .B(n539), .Z(product[5]) );
  XNOR2_X1 U756 ( .A(n57), .B(n112), .ZN(product[4]) );
  OAI21_X1 U757 ( .B1(n64), .B2(n550), .A(n65), .ZN(n63) );
  OAI21_X1 U758 ( .B1(n45), .B2(n506), .A(n72), .ZN(n70) );
  OAI21_X1 U759 ( .B1(n571), .B2(n553), .A(n79), .ZN(n77) );
  XNOR2_X1 U760 ( .A(n556), .B(n53), .ZN(product[8]) );
  AOI21_X1 U761 ( .B1(n555), .B2(n575), .A(n93), .ZN(n91) );
  XOR2_X1 U762 ( .A(n58), .B(n115), .Z(product[3]) );
  OAI22_X1 U763 ( .A1(n531), .A2(n395), .B1(n394), .B2(n588), .ZN(n316) );
  OAI22_X1 U764 ( .A1(n531), .A2(n394), .B1(n393), .B2(n588), .ZN(n315) );
  OAI22_X1 U765 ( .A1(n6), .A2(n396), .B1(n395), .B2(n588), .ZN(n317) );
  OAI22_X1 U766 ( .A1(n531), .A2(n397), .B1(n396), .B2(n588), .ZN(n318) );
  OAI22_X1 U767 ( .A1(n531), .A2(n398), .B1(n397), .B2(n588), .ZN(n319) );
  OAI22_X1 U768 ( .A1(n531), .A2(n400), .B1(n399), .B2(n588), .ZN(n321) );
  OAI22_X1 U769 ( .A1(n6), .A2(n399), .B1(n398), .B2(n588), .ZN(n320) );
  OAI22_X1 U770 ( .A1(n531), .A2(n401), .B1(n400), .B2(n588), .ZN(n322) );
  OAI22_X1 U771 ( .A1(n531), .A2(n402), .B1(n401), .B2(n588), .ZN(n323) );
  NAND2_X1 U772 ( .A1(n329), .A2(n258), .ZN(n122) );
  OAI22_X1 U773 ( .A1(n6), .A2(n404), .B1(n403), .B2(n588), .ZN(n325) );
  OAI22_X1 U774 ( .A1(n6), .A2(n403), .B1(n402), .B2(n588), .ZN(n324) );
  OAI22_X1 U775 ( .A1(n531), .A2(n406), .B1(n405), .B2(n588), .ZN(n327) );
  OAI22_X1 U776 ( .A1(n531), .A2(n405), .B1(n404), .B2(n588), .ZN(n326) );
  OAI22_X1 U777 ( .A1(n531), .A2(n407), .B1(n406), .B2(n588), .ZN(n328) );
  OAI22_X1 U778 ( .A1(n531), .A2(n408), .B1(n407), .B2(n588), .ZN(n329) );
  OAI22_X1 U779 ( .A1(n531), .A2(n524), .B1(n409), .B2(n588), .ZN(n258) );
  OAI22_X1 U780 ( .A1(n557), .A2(n379), .B1(n378), .B2(n551), .ZN(n301) );
  OAI22_X1 U781 ( .A1(n557), .A2(n380), .B1(n379), .B2(n551), .ZN(n302) );
  OAI22_X1 U782 ( .A1(n557), .A2(n385), .B1(n384), .B2(n551), .ZN(n307) );
  OAI22_X1 U783 ( .A1(n557), .A2(n382), .B1(n381), .B2(n585), .ZN(n304) );
  OAI22_X1 U784 ( .A1(n557), .A2(n381), .B1(n380), .B2(n585), .ZN(n303) );
  NAND2_X1 U785 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U786 ( .A1(n383), .A2(n558), .B1(n382), .B2(n500), .ZN(n305) );
  OAI22_X1 U787 ( .A1(n558), .A2(n384), .B1(n383), .B2(n500), .ZN(n306) );
  OAI22_X1 U788 ( .A1(n557), .A2(n386), .B1(n385), .B2(n500), .ZN(n308) );
  OAI22_X1 U789 ( .A1(n557), .A2(n387), .B1(n386), .B2(n500), .ZN(n309) );
  OAI22_X1 U790 ( .A1(n557), .A2(n535), .B1(n392), .B2(n551), .ZN(n257) );
  OAI22_X1 U791 ( .A1(n558), .A2(n389), .B1(n388), .B2(n585), .ZN(n311) );
  OAI22_X1 U792 ( .A1(n558), .A2(n388), .B1(n387), .B2(n585), .ZN(n310) );
  OAI22_X1 U793 ( .A1(n558), .A2(n390), .B1(n389), .B2(n500), .ZN(n312) );
  INV_X1 U794 ( .A(n500), .ZN(n247) );
  OAI22_X1 U795 ( .A1(n499), .A2(n391), .B1(n390), .B2(n585), .ZN(n313) );
  INV_X1 U796 ( .A(n597), .ZN(n596) );
  INV_X1 U797 ( .A(n603), .ZN(n602) );
  INV_X1 U798 ( .A(n31), .ZN(n603) );
  INV_X1 U799 ( .A(n36), .ZN(n605) );
  INV_X1 U800 ( .A(n607), .ZN(n606) );
  INV_X1 U801 ( .A(n40), .ZN(n607) );
  XOR2_X1 U802 ( .A(n259), .B(n251), .Z(n148) );
  XOR2_X1 U803 ( .A(n159), .B(n150), .Z(n142) );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_12_DW01_add_2 ( A, B, CI, 
        SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n5, n8, n9, n10, n11, n12, n13, n14, n15, n16, n19, n20, n22,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n44, n45, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n65, n67, n68, n69, n70, n71, n73, n75,
         n76, n77, n78, n79, n81, n83, n84, n86, n88, n89, n90, n94, n95, n96,
         n98, n100, n157, n158, n159, n160, n161, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181;

  NOR2_X1 U122 ( .A1(A[8]), .A2(B[8]), .ZN(n157) );
  NOR2_X1 U123 ( .A1(A[8]), .A2(B[8]), .ZN(n54) );
  XNOR2_X1 U124 ( .A(n45), .B(n158), .ZN(SUM[10]) );
  AND2_X1 U125 ( .A1(n165), .A2(n44), .ZN(n158) );
  AOI21_X1 U126 ( .B1(n60), .B2(n52), .A(n53), .ZN(n159) );
  NOR2_X1 U127 ( .A1(A[11]), .A2(B[11]), .ZN(n160) );
  XNOR2_X1 U128 ( .A(n37), .B(n161), .ZN(SUM[11]) );
  AND2_X1 U129 ( .A1(n164), .A2(n36), .ZN(n161) );
  AND2_X1 U130 ( .A1(n173), .A2(n86), .ZN(SUM[0]) );
  OR2_X1 U131 ( .A1(A[15]), .A2(B[15]), .ZN(n163) );
  OR2_X2 U132 ( .A1(A[9]), .A2(B[9]), .ZN(n177) );
  INV_X1 U133 ( .A(n160), .ZN(n164) );
  OR2_X1 U134 ( .A1(A[10]), .A2(B[10]), .ZN(n165) );
  OR2_X1 U135 ( .A1(A[10]), .A2(B[10]), .ZN(n179) );
  AND2_X1 U136 ( .A1(A[9]), .A2(B[9]), .ZN(n166) );
  XNOR2_X1 U137 ( .A(n172), .B(n167), .ZN(SUM[13]) );
  AND2_X1 U138 ( .A1(n89), .A2(n29), .ZN(n167) );
  BUF_X1 U139 ( .A(n33), .Z(n168) );
  NOR2_X1 U140 ( .A1(A[12]), .A2(B[12]), .ZN(n169) );
  NOR2_X1 U141 ( .A1(A[12]), .A2(B[12]), .ZN(n32) );
  NOR2_X1 U142 ( .A1(A[14]), .A2(B[14]), .ZN(n170) );
  AOI21_X1 U143 ( .B1(n38), .B2(n30), .A(n31), .ZN(n171) );
  AOI21_X1 U144 ( .B1(n38), .B2(n30), .A(n31), .ZN(n172) );
  INV_X1 U145 ( .A(n24), .ZN(n22) );
  OR2_X1 U146 ( .A1(A[0]), .A2(B[0]), .ZN(n173) );
  INV_X1 U147 ( .A(n60), .ZN(n59) );
  INV_X1 U148 ( .A(n159), .ZN(n50) );
  INV_X1 U149 ( .A(n38), .ZN(n37) );
  AOI21_X1 U150 ( .B1(n175), .B2(n76), .A(n73), .ZN(n71) );
  INV_X1 U151 ( .A(n75), .ZN(n73) );
  OAI21_X1 U152 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  AOI21_X1 U153 ( .B1(n178), .B2(n84), .A(n81), .ZN(n79) );
  INV_X1 U154 ( .A(n83), .ZN(n81) );
  AOI21_X1 U155 ( .B1(n52), .B2(n60), .A(n53), .ZN(n51) );
  OAI21_X1 U156 ( .B1(n71), .B2(n69), .A(n70), .ZN(n68) );
  OR2_X1 U157 ( .A1(n170), .A2(n28), .ZN(n174) );
  OAI21_X1 U158 ( .B1(n79), .B2(n77), .A(n78), .ZN(n76) );
  AOI21_X1 U159 ( .B1(n176), .B2(n68), .A(n65), .ZN(n63) );
  INV_X1 U160 ( .A(n67), .ZN(n65) );
  AOI21_X1 U161 ( .B1(n50), .B2(n177), .A(n166), .ZN(n45) );
  NAND2_X1 U162 ( .A1(n94), .A2(n55), .ZN(n9) );
  INV_X1 U163 ( .A(n86), .ZN(n84) );
  OAI21_X1 U164 ( .B1(n59), .B2(n57), .A(n58), .ZN(n56) );
  NAND2_X1 U165 ( .A1(n98), .A2(n70), .ZN(n13) );
  INV_X1 U166 ( .A(n69), .ZN(n98) );
  NAND2_X1 U167 ( .A1(n96), .A2(n62), .ZN(n11) );
  INV_X1 U168 ( .A(n61), .ZN(n96) );
  INV_X1 U169 ( .A(n169), .ZN(n90) );
  NAND2_X1 U170 ( .A1(n177), .A2(n49), .ZN(n8) );
  NAND2_X1 U171 ( .A1(n176), .A2(n67), .ZN(n12) );
  NAND2_X1 U172 ( .A1(n95), .A2(n58), .ZN(n10) );
  INV_X1 U173 ( .A(n57), .ZN(n95) );
  NAND2_X1 U174 ( .A1(n100), .A2(n78), .ZN(n15) );
  INV_X1 U175 ( .A(n77), .ZN(n100) );
  NAND2_X1 U176 ( .A1(n175), .A2(n75), .ZN(n14) );
  NAND2_X1 U177 ( .A1(n178), .A2(n83), .ZN(n16) );
  XNOR2_X1 U178 ( .A(n56), .B(n9), .ZN(SUM[8]) );
  XNOR2_X1 U179 ( .A(n50), .B(n8), .ZN(SUM[9]) );
  XOR2_X1 U180 ( .A(n59), .B(n10), .Z(SUM[7]) );
  OR2_X1 U181 ( .A1(A[3]), .A2(B[3]), .ZN(n175) );
  OR2_X1 U182 ( .A1(A[5]), .A2(B[5]), .ZN(n176) );
  NOR2_X1 U183 ( .A1(A[7]), .A2(B[7]), .ZN(n57) );
  NOR2_X1 U184 ( .A1(A[14]), .A2(B[14]), .ZN(n25) );
  NOR2_X1 U185 ( .A1(A[2]), .A2(B[2]), .ZN(n77) );
  NOR2_X1 U186 ( .A1(A[4]), .A2(B[4]), .ZN(n69) );
  NAND2_X1 U187 ( .A1(n88), .A2(n26), .ZN(n3) );
  NAND2_X1 U188 ( .A1(n90), .A2(n168), .ZN(n5) );
  OR2_X1 U189 ( .A1(A[1]), .A2(B[1]), .ZN(n178) );
  NOR2_X1 U190 ( .A1(A[6]), .A2(B[6]), .ZN(n61) );
  XNOR2_X1 U191 ( .A(n12), .B(n68), .ZN(SUM[5]) );
  XNOR2_X1 U192 ( .A(n16), .B(n84), .ZN(SUM[1]) );
  NAND2_X1 U193 ( .A1(A[7]), .A2(B[7]), .ZN(n58) );
  NAND2_X1 U194 ( .A1(A[2]), .A2(B[2]), .ZN(n78) );
  NAND2_X1 U195 ( .A1(A[4]), .A2(B[4]), .ZN(n70) );
  NAND2_X1 U196 ( .A1(A[1]), .A2(B[1]), .ZN(n83) );
  NAND2_X1 U197 ( .A1(A[0]), .A2(B[0]), .ZN(n86) );
  NAND2_X1 U198 ( .A1(A[6]), .A2(B[6]), .ZN(n62) );
  NAND2_X1 U199 ( .A1(A[3]), .A2(B[3]), .ZN(n75) );
  NAND2_X1 U200 ( .A1(A[14]), .A2(B[14]), .ZN(n26) );
  XOR2_X1 U201 ( .A(n13), .B(n71), .Z(SUM[4]) );
  XNOR2_X1 U202 ( .A(n14), .B(n76), .ZN(SUM[3]) );
  XOR2_X1 U203 ( .A(n15), .B(n79), .Z(SUM[2]) );
  NAND2_X1 U204 ( .A1(n163), .A2(n19), .ZN(n2) );
  NAND2_X1 U205 ( .A1(A[15]), .A2(B[15]), .ZN(n19) );
  XOR2_X1 U206 ( .A(n11), .B(n63), .Z(SUM[6]) );
  NAND2_X1 U207 ( .A1(A[5]), .A2(B[5]), .ZN(n67) );
  XNOR2_X1 U208 ( .A(n34), .B(n5), .ZN(SUM[12]) );
  INV_X1 U209 ( .A(n181), .ZN(n44) );
  NAND2_X1 U210 ( .A1(A[13]), .A2(B[13]), .ZN(n29) );
  AOI21_X1 U211 ( .B1(n179), .B2(n166), .A(n181), .ZN(n40) );
  INV_X1 U212 ( .A(n89), .ZN(n180) );
  INV_X1 U213 ( .A(n28), .ZN(n89) );
  NOR2_X1 U214 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  NAND2_X1 U215 ( .A1(A[12]), .A2(B[12]), .ZN(n33) );
  NAND2_X1 U216 ( .A1(A[9]), .A2(B[9]), .ZN(n49) );
  AND2_X1 U217 ( .A1(A[10]), .A2(B[10]), .ZN(n181) );
  INV_X1 U218 ( .A(n157), .ZN(n94) );
  NOR2_X1 U219 ( .A1(n157), .A2(n57), .ZN(n52) );
  OAI21_X1 U220 ( .B1(n54), .B2(n58), .A(n55), .ZN(n53) );
  NAND2_X1 U221 ( .A1(A[8]), .A2(B[8]), .ZN(n55) );
  OAI21_X1 U222 ( .B1(n32), .B2(n36), .A(n33), .ZN(n31) );
  NAND2_X1 U223 ( .A1(A[11]), .A2(B[11]), .ZN(n36) );
  INV_X1 U224 ( .A(n170), .ZN(n88) );
  OAI21_X1 U225 ( .B1(n25), .B2(n29), .A(n26), .ZN(n24) );
  NOR2_X1 U226 ( .A1(A[11]), .A2(B[11]), .ZN(n35) );
  NOR2_X1 U227 ( .A1(n169), .A2(n35), .ZN(n30) );
  OAI21_X1 U228 ( .B1(n37), .B2(n35), .A(n36), .ZN(n34) );
  OAI21_X1 U229 ( .B1(n39), .B2(n51), .A(n40), .ZN(n38) );
  NAND2_X1 U230 ( .A1(n165), .A2(n177), .ZN(n39) );
  XNOR2_X1 U231 ( .A(n20), .B(n2), .ZN(SUM[15]) );
  XNOR2_X1 U232 ( .A(n27), .B(n3), .ZN(SUM[14]) );
  OAI21_X1 U233 ( .B1(n171), .B2(n180), .A(n29), .ZN(n27) );
  OAI21_X1 U234 ( .B1(n172), .B2(n174), .A(n22), .ZN(n20) );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_12 ( clk, clear_acc, 
        data_out_x, data_out, data_out_w, data_out_b, wr_en_y, m_valid, 
        m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [4:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
         N39, N40, N41, N42, N43, N44, n1, n2, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n85, n102, n111, n112, n113, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n21), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n224), .CK(clk), .Q(n25) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n225), .CK(clk), .Q(n26) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n226), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n227), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n228), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n229), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n230), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n231), .CK(clk), .Q(n34) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n232), .CK(clk), .Q(n35) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n233), .CK(clk), .Q(n36) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n234), .CK(clk), .Q(n37) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n235), .CK(clk), .Q(n38) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n236), .CK(clk), .Q(n39) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n237), .CK(clk), .Q(n40) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n238), .CK(clk), .Q(n41) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n239), .CK(clk), .Q(n43) );
  DFF_X1 \f_reg[0]  ( .D(n111), .CK(clk), .Q(f[0]), .QN(n212) );
  DFF_X1 \f_reg[1]  ( .D(n102), .CK(clk), .Q(f[1]), .QN(n213) );
  DFF_X1 \f_reg[2]  ( .D(n85), .CK(clk), .Q(f[2]), .QN(n214) );
  DFF_X1 \f_reg[3]  ( .D(n83), .CK(clk), .Q(f[3]), .QN(n215) );
  DFF_X1 \f_reg[7]  ( .D(n79), .CK(clk), .Q(f[7]), .QN(n216) );
  DFF_X1 \f_reg[8]  ( .D(n78), .CK(clk), .Q(f[8]), .QN(n217) );
  DFF_X1 \f_reg[9]  ( .D(n77), .CK(clk), .Q(f[9]), .QN(n218) );
  DFF_X1 \f_reg[10]  ( .D(n76), .CK(clk), .Q(n52), .QN(n219) );
  DFF_X1 \f_reg[11]  ( .D(n75), .CK(clk), .Q(n50), .QN(n220) );
  DFF_X1 \f_reg[12]  ( .D(n1), .CK(clk), .Q(n49), .QN(n221) );
  DFF_X1 \f_reg[13]  ( .D(n16), .CK(clk), .Q(n48), .QN(n222) );
  DFF_X1 \f_reg[14]  ( .D(n4), .CK(clk), .Q(n47), .QN(n223) );
  DFF_X1 \f_reg[15]  ( .D(n5), .CK(clk), .Q(f[15]), .QN(n72) );
  DFF_X1 \data_out_reg[15]  ( .D(n113), .CK(clk), .Q(data_out[15]), .QN(n195)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n165), .CK(clk), .Q(data_out[14]), .QN(n194)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n166), .CK(clk), .Q(data_out[13]), .QN(n193)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n167), .CK(clk), .Q(data_out[12]), .QN(n192)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n168), .CK(clk), .Q(data_out[11]), .QN(n191)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n169), .CK(clk), .Q(data_out[10]), .QN(n190)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n170), .CK(clk), .Q(data_out[9]), .QN(n189) );
  DFF_X1 \data_out_reg[8]  ( .D(n171), .CK(clk), .Q(data_out[8]), .QN(n188) );
  DFF_X1 \data_out_reg[7]  ( .D(n172), .CK(clk), .Q(data_out[7]), .QN(n187) );
  DFF_X1 \data_out_reg[6]  ( .D(n173), .CK(clk), .Q(data_out[6]), .QN(n186) );
  DFF_X1 \data_out_reg[5]  ( .D(n174), .CK(clk), .Q(data_out[5]), .QN(n185) );
  DFF_X1 \data_out_reg[4]  ( .D(n175), .CK(clk), .Q(data_out[4]), .QN(n184) );
  DFF_X1 \data_out_reg[3]  ( .D(n176), .CK(clk), .Q(data_out[3]), .QN(n183) );
  DFF_X1 \data_out_reg[2]  ( .D(n177), .CK(clk), .Q(data_out[2]), .QN(n182) );
  DFF_X1 \data_out_reg[1]  ( .D(n178), .CK(clk), .Q(data_out[1]), .QN(n181) );
  DFF_X1 \data_out_reg[0]  ( .D(n179), .CK(clk), .Q(data_out[0]), .QN(n180) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_12_DW_mult_tc_1 mult_2021 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_12_DW01_add_2 add_2022 ( .A({
        n202, n201, n200, n199, n198, n197, n211, n210, n209, n208, n207, n206, 
        n205, n204, n203, n196}), .B({f[15], n47, n48, n49, n50, n52, f[9:0]}), 
        .CI(1'b0), .SUM(adder) );
  DFF_X1 \f_reg[4]  ( .D(n82), .CK(clk), .Q(f[4]), .QN(n65) );
  DFF_X1 \f_reg[5]  ( .D(n81), .CK(clk), .Q(f[5]), .QN(n66) );
  DFF_X1 \f_reg[6]  ( .D(n80), .CK(clk), .Q(f[6]), .QN(n67) );
  DFF_X2 delay_reg ( .D(n112), .CK(clk), .Q(n2), .QN(n240) );
  MUX2_X2 U3 ( .A(n29), .B(N40), .S(n240), .Z(n198) );
  MUX2_X1 U4 ( .A(N39), .B(n32), .S(n2), .Z(n197) );
  AND2_X1 U5 ( .A1(n46), .A2(n22), .ZN(n15) );
  NAND3_X1 U6 ( .A1(n13), .A2(n12), .A3(n14), .ZN(n1) );
  MUX2_X2 U8 ( .A(n33), .B(N38), .S(n240), .Z(n211) );
  MUX2_X2 U9 ( .A(N41), .B(n28), .S(n2), .Z(n199) );
  NAND3_X1 U10 ( .A1(n7), .A2(n6), .A3(n8), .ZN(n4) );
  MUX2_X2 U11 ( .A(n34), .B(N37), .S(n240), .Z(n210) );
  NAND3_X1 U12 ( .A1(n10), .A2(n9), .A3(n11), .ZN(n5) );
  NAND2_X1 U13 ( .A1(data_out_b[14]), .A2(n21), .ZN(n6) );
  NAND2_X1 U14 ( .A1(adder[14]), .A2(n15), .ZN(n7) );
  NAND2_X1 U15 ( .A1(n63), .A2(n47), .ZN(n8) );
  NAND2_X1 U16 ( .A1(data_out_b[15]), .A2(n21), .ZN(n9) );
  NAND2_X1 U17 ( .A1(adder[15]), .A2(n15), .ZN(n10) );
  NAND2_X1 U18 ( .A1(n63), .A2(f[15]), .ZN(n11) );
  MUX2_X2 U19 ( .A(n26), .B(N43), .S(n240), .Z(n201) );
  NAND2_X1 U20 ( .A1(data_out_b[12]), .A2(n21), .ZN(n12) );
  NAND2_X1 U21 ( .A1(adder[12]), .A2(n15), .ZN(n13) );
  NAND2_X1 U22 ( .A1(n63), .A2(n49), .ZN(n14) );
  NAND2_X1 U23 ( .A1(n112), .A2(n20), .ZN(n242) );
  INV_X1 U24 ( .A(clear_acc), .ZN(n22) );
  INV_X1 U25 ( .A(n24), .ZN(n42) );
  OAI22_X1 U26 ( .A1(n183), .A2(n242), .B1(n215), .B2(n241), .ZN(n176) );
  OAI22_X1 U27 ( .A1(n184), .A2(n242), .B1(n65), .B2(n241), .ZN(n175) );
  OAI22_X1 U28 ( .A1(n185), .A2(n242), .B1(n66), .B2(n241), .ZN(n174) );
  OAI22_X1 U29 ( .A1(n186), .A2(n242), .B1(n67), .B2(n241), .ZN(n173) );
  OAI22_X1 U30 ( .A1(n187), .A2(n242), .B1(n216), .B2(n241), .ZN(n172) );
  OAI22_X1 U31 ( .A1(n188), .A2(n242), .B1(n217), .B2(n241), .ZN(n171) );
  OAI22_X1 U32 ( .A1(n189), .A2(n242), .B1(n218), .B2(n241), .ZN(n170) );
  MUX2_X1 U33 ( .A(n39), .B(N32), .S(n240), .Z(n205) );
  NAND3_X1 U34 ( .A1(n18), .A2(n17), .A3(n19), .ZN(n16) );
  NAND2_X1 U35 ( .A1(data_out_b[13]), .A2(n21), .ZN(n17) );
  NAND2_X1 U36 ( .A1(adder[13]), .A2(n15), .ZN(n18) );
  NAND2_X1 U37 ( .A1(n63), .A2(n48), .ZN(n19) );
  INV_X1 U38 ( .A(n22), .ZN(n21) );
  INV_X1 U39 ( .A(n46), .ZN(n63) );
  INV_X1 U40 ( .A(wr_en_y), .ZN(n20) );
  INV_X1 U41 ( .A(m_ready), .ZN(n23) );
  NAND2_X1 U42 ( .A1(m_valid), .A2(n23), .ZN(n44) );
  OAI21_X1 U43 ( .B1(sel[4]), .B2(n74), .A(n44), .ZN(n112) );
  NAND2_X1 U44 ( .A1(clear_acc_delay), .A2(n240), .ZN(n24) );
  MUX2_X1 U45 ( .A(n25), .B(N44), .S(n42), .Z(n224) );
  MUX2_X1 U46 ( .A(n25), .B(N44), .S(n240), .Z(n202) );
  MUX2_X1 U47 ( .A(n26), .B(N43), .S(n42), .Z(n225) );
  MUX2_X1 U48 ( .A(n27), .B(N42), .S(n42), .Z(n226) );
  MUX2_X1 U49 ( .A(n27), .B(N42), .S(n240), .Z(n200) );
  MUX2_X1 U50 ( .A(n28), .B(N41), .S(n42), .Z(n227) );
  MUX2_X1 U51 ( .A(n29), .B(N40), .S(n42), .Z(n228) );
  MUX2_X1 U52 ( .A(n32), .B(N39), .S(n42), .Z(n229) );
  MUX2_X1 U53 ( .A(n33), .B(N38), .S(n42), .Z(n230) );
  MUX2_X1 U54 ( .A(n34), .B(N37), .S(n42), .Z(n231) );
  MUX2_X1 U55 ( .A(n35), .B(N36), .S(n42), .Z(n232) );
  MUX2_X1 U56 ( .A(n35), .B(N36), .S(n240), .Z(n209) );
  MUX2_X1 U57 ( .A(n36), .B(N35), .S(n42), .Z(n233) );
  MUX2_X1 U58 ( .A(n36), .B(N35), .S(n240), .Z(n208) );
  MUX2_X1 U59 ( .A(n37), .B(N34), .S(n42), .Z(n234) );
  MUX2_X1 U60 ( .A(n37), .B(N34), .S(n240), .Z(n207) );
  MUX2_X1 U61 ( .A(n38), .B(N33), .S(n42), .Z(n235) );
  MUX2_X1 U62 ( .A(n38), .B(N33), .S(n240), .Z(n206) );
  MUX2_X1 U63 ( .A(n39), .B(N32), .S(n42), .Z(n236) );
  MUX2_X1 U64 ( .A(n40), .B(N31), .S(n42), .Z(n237) );
  MUX2_X1 U65 ( .A(n40), .B(N31), .S(n240), .Z(n204) );
  MUX2_X1 U66 ( .A(n41), .B(N30), .S(n42), .Z(n238) );
  MUX2_X1 U67 ( .A(n41), .B(N30), .S(n240), .Z(n203) );
  MUX2_X1 U68 ( .A(n43), .B(N29), .S(n42), .Z(n239) );
  MUX2_X1 U69 ( .A(n43), .B(N29), .S(n240), .Z(n196) );
  INV_X1 U70 ( .A(n44), .ZN(n45) );
  OAI21_X1 U71 ( .B1(n45), .B2(n2), .A(n22), .ZN(n46) );
  AOI222_X1 U72 ( .A1(data_out_b[11]), .A2(n21), .B1(adder[11]), .B2(n15), 
        .C1(n63), .C2(n50), .ZN(n51) );
  INV_X1 U73 ( .A(n51), .ZN(n75) );
  AOI222_X1 U74 ( .A1(data_out_b[10]), .A2(n21), .B1(adder[10]), .B2(n15), 
        .C1(n63), .C2(n52), .ZN(n53) );
  INV_X1 U75 ( .A(n53), .ZN(n76) );
  AOI222_X1 U76 ( .A1(data_out_b[8]), .A2(n21), .B1(adder[8]), .B2(n15), .C1(
        n63), .C2(f[8]), .ZN(n54) );
  INV_X1 U77 ( .A(n54), .ZN(n78) );
  AOI222_X1 U78 ( .A1(data_out_b[7]), .A2(n21), .B1(adder[7]), .B2(n15), .C1(
        n63), .C2(f[7]), .ZN(n55) );
  INV_X1 U79 ( .A(n55), .ZN(n79) );
  AOI222_X1 U80 ( .A1(data_out_b[6]), .A2(n21), .B1(adder[6]), .B2(n15), .C1(
        n63), .C2(f[6]), .ZN(n56) );
  INV_X1 U81 ( .A(n56), .ZN(n80) );
  AOI222_X1 U82 ( .A1(data_out_b[5]), .A2(n21), .B1(adder[5]), .B2(n15), .C1(
        n63), .C2(f[5]), .ZN(n57) );
  INV_X1 U83 ( .A(n57), .ZN(n81) );
  AOI222_X1 U84 ( .A1(data_out_b[4]), .A2(n21), .B1(adder[4]), .B2(n15), .C1(
        n63), .C2(f[4]), .ZN(n58) );
  INV_X1 U85 ( .A(n58), .ZN(n82) );
  AOI222_X1 U86 ( .A1(data_out_b[3]), .A2(n21), .B1(adder[3]), .B2(n15), .C1(
        n63), .C2(f[3]), .ZN(n59) );
  INV_X1 U87 ( .A(n59), .ZN(n83) );
  AOI222_X1 U88 ( .A1(data_out_b[2]), .A2(n21), .B1(adder[2]), .B2(n15), .C1(
        n63), .C2(f[2]), .ZN(n60) );
  INV_X1 U89 ( .A(n60), .ZN(n85) );
  AOI222_X1 U90 ( .A1(data_out_b[1]), .A2(n21), .B1(adder[1]), .B2(n15), .C1(
        n63), .C2(f[1]), .ZN(n61) );
  INV_X1 U91 ( .A(n61), .ZN(n102) );
  AOI222_X1 U92 ( .A1(data_out_b[0]), .A2(n21), .B1(adder[0]), .B2(n15), .C1(
        n63), .C2(f[0]), .ZN(n62) );
  INV_X1 U93 ( .A(n62), .ZN(n111) );
  AOI222_X1 U94 ( .A1(data_out_b[9]), .A2(n21), .B1(adder[9]), .B2(n15), .C1(
        n63), .C2(f[9]), .ZN(n64) );
  INV_X1 U95 ( .A(n64), .ZN(n77) );
  NOR4_X1 U96 ( .A1(n50), .A2(n49), .A3(n48), .A4(n47), .ZN(n71) );
  NOR4_X1 U97 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n52), .ZN(n70) );
  NAND4_X1 U98 ( .A1(n67), .A2(n66), .A3(n65), .A4(n215), .ZN(n68) );
  NOR4_X1 U99 ( .A1(n68), .A2(f[0]), .A3(f[1]), .A4(f[2]), .ZN(n69) );
  NAND3_X1 U100 ( .A1(n71), .A2(n70), .A3(n69), .ZN(n73) );
  NAND3_X1 U101 ( .A1(wr_en_y), .A2(n73), .A3(n72), .ZN(n241) );
  OAI22_X1 U102 ( .A1(n180), .A2(n242), .B1(n212), .B2(n241), .ZN(n179) );
  OAI22_X1 U103 ( .A1(n181), .A2(n242), .B1(n213), .B2(n241), .ZN(n178) );
  OAI22_X1 U104 ( .A1(n182), .A2(n242), .B1(n214), .B2(n241), .ZN(n177) );
  OAI22_X1 U105 ( .A1(n190), .A2(n242), .B1(n219), .B2(n241), .ZN(n169) );
  OAI22_X1 U106 ( .A1(n191), .A2(n242), .B1(n220), .B2(n241), .ZN(n168) );
  OAI22_X1 U107 ( .A1(n192), .A2(n242), .B1(n221), .B2(n241), .ZN(n167) );
  OAI22_X1 U108 ( .A1(n193), .A2(n242), .B1(n222), .B2(n241), .ZN(n166) );
  OAI22_X1 U109 ( .A1(n194), .A2(n242), .B1(n223), .B2(n241), .ZN(n165) );
  OAI22_X1 U110 ( .A1(n195), .A2(n242), .B1(n72), .B2(n241), .ZN(n113) );
  AND4_X1 U111 ( .A1(sel[3]), .A2(sel[2]), .A3(sel[1]), .A4(sel[0]), .ZN(n74)
         );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_11_DW_mult_tc_1 ( a, b, 
        product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n9, n12, n13, n16, n18, n19, n21, n23, n25, n29, n31, n32,
         n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n50, n53, n54,
         n55, n56, n57, n58, n59, n62, n63, n64, n65, n67, n69, n70, n71, n72,
         n73, n74, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n93, n95, n96, n97, n98, n99, n101, n103, n104,
         n105, n106, n107, n109, n111, n112, n113, n114, n115, n117, n119,
         n120, n122, n127, n131, n135, n139, n141, n142, n143, n144, n145,
         n146, n148, n149, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n245, n247, n249, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n418, n419, n420,
         n421, n422, n423, n424, n426, n427, n428, n429, n433, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U148 ( .A(n265), .B(n144), .Z(n145) );
  XOR2_X1 U152 ( .A(n301), .B(n148), .Z(n149) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U162 ( .A(n170), .B(n172), .CI(n179), .CO(n165), .S(n166) );
  FA_X1 U163 ( .A(n181), .B(n174), .CI(n183), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n263), .CI(n291), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n252), .B(n317), .CO(n173), .S(n174) );
  FA_X1 U167 ( .A(n180), .B(n187), .CI(n178), .CO(n175), .S(n176) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U169 ( .A(n193), .B(n282), .CI(n191), .CO(n179), .S(n180) );
  FA_X1 U170 ( .A(n268), .B(n274), .CI(n292), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n304), .B(n264), .CI(n318), .CO(n183), .S(n184) );
  FA_X1 U172 ( .A(n197), .B(n190), .CI(n188), .CO(n185), .S(n186) );
  FA_X1 U173 ( .A(n199), .B(n201), .CI(n192), .CO(n187), .S(n188) );
  FA_X1 U174 ( .A(n275), .B(n293), .CI(n194), .CO(n189), .S(n190) );
  FA_X1 U175 ( .A(n253), .B(n305), .CI(n283), .CO(n191), .S(n192) );
  HA_X1 U176 ( .A(n319), .B(n269), .CO(n193), .S(n194) );
  FA_X1 U177 ( .A(n205), .B(n200), .CI(n198), .CO(n195), .S(n196) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U179 ( .A(n276), .B(n284), .CI(n294), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n320), .B(n270), .CI(n306), .CO(n201), .S(n202) );
  FA_X1 U181 ( .A(n208), .B(n213), .CI(n206), .CO(n203), .S(n204) );
  FA_X1 U182 ( .A(n210), .B(n307), .CI(n215), .CO(n205), .S(n206) );
  FA_X1 U183 ( .A(n285), .B(n254), .CI(n295), .CO(n207), .S(n208) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n322), .B(n278), .CI(n308), .CO(n215), .S(n216) );
  FA_X1 U188 ( .A(n225), .B(n222), .CI(n220), .CO(n217), .S(n218) );
  FA_X1 U189 ( .A(n255), .B(n309), .CI(n297), .CO(n219), .S(n220) );
  HA_X1 U190 ( .A(n287), .B(n323), .CO(n221), .S(n222) );
  FA_X1 U192 ( .A(n324), .B(n288), .CI(n310), .CO(n225), .S(n226) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  HA_X1 U194 ( .A(n311), .B(n325), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n326), .B(n300), .CI(n312), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  INV_X1 U414 ( .A(n529), .ZN(n490) );
  CLKBUF_X1 U415 ( .A(n18), .Z(n491) );
  BUF_X2 U416 ( .A(n18), .Z(n492) );
  NAND2_X1 U417 ( .A1(n16), .A2(n567), .ZN(n18) );
  XOR2_X1 U418 ( .A(n158), .B(n160), .Z(n493) );
  XOR2_X1 U419 ( .A(n493), .B(n167), .Z(n154) );
  XOR2_X1 U420 ( .A(n156), .B(n165), .Z(n494) );
  XOR2_X1 U421 ( .A(n494), .B(n154), .Z(n152) );
  NAND2_X1 U422 ( .A1(n158), .A2(n160), .ZN(n495) );
  NAND2_X1 U423 ( .A1(n158), .A2(n167), .ZN(n496) );
  NAND2_X1 U424 ( .A1(n160), .A2(n167), .ZN(n497) );
  NAND3_X1 U425 ( .A1(n495), .A2(n496), .A3(n497), .ZN(n153) );
  NAND2_X1 U426 ( .A1(n156), .A2(n165), .ZN(n498) );
  NAND2_X1 U427 ( .A1(n156), .A2(n154), .ZN(n499) );
  NAND2_X1 U428 ( .A1(n165), .A2(n154), .ZN(n500) );
  NAND3_X1 U429 ( .A1(n498), .A2(n499), .A3(n500), .ZN(n151) );
  BUF_X1 U430 ( .A(n86), .Z(n501) );
  OR2_X1 U431 ( .A1(n164), .A2(n175), .ZN(n502) );
  OR2_X1 U432 ( .A1(n329), .A2(n258), .ZN(n503) );
  CLKBUF_X1 U433 ( .A(n12), .Z(n509) );
  BUF_X1 U434 ( .A(n96), .Z(n557) );
  XOR2_X1 U435 ( .A(n600), .B(a[14]), .Z(n41) );
  INV_X1 U436 ( .A(n600), .ZN(n599) );
  OR2_X1 U437 ( .A1(n204), .A2(n211), .ZN(n504) );
  OAI21_X1 U438 ( .B1(n553), .B2(n79), .A(n76), .ZN(n505) );
  BUF_X1 U439 ( .A(n12), .Z(n535) );
  XOR2_X1 U440 ( .A(n594), .B(a[8]), .Z(n506) );
  OAI21_X1 U441 ( .B1(n99), .B2(n97), .A(n98), .ZN(n96) );
  AND2_X1 U442 ( .A1(n427), .A2(n507), .ZN(n515) );
  NOR2_X1 U443 ( .A1(n528), .A2(n600), .ZN(n507) );
  INV_X1 U444 ( .A(n524), .ZN(n508) );
  BUF_X1 U445 ( .A(n588), .Z(n524) );
  INV_X1 U446 ( .A(n596), .ZN(n510) );
  XNOR2_X1 U447 ( .A(n88), .B(n511), .ZN(product[10]) );
  NAND2_X1 U448 ( .A1(n547), .A2(n86), .ZN(n511) );
  AOI21_X1 U449 ( .B1(n96), .B2(n572), .A(n93), .ZN(n512) );
  INV_X1 U450 ( .A(n514), .ZN(n513) );
  CLKBUF_X1 U451 ( .A(n528), .Z(n514) );
  NOR2_X1 U452 ( .A1(n337), .A2(n37), .ZN(n516) );
  OR2_X1 U453 ( .A1(n515), .A2(n516), .ZN(n252) );
  INV_X1 U454 ( .A(n528), .ZN(n37) );
  OR2_X2 U455 ( .A1(n152), .A2(n163), .ZN(n571) );
  XOR2_X1 U456 ( .A(n512), .B(n517), .Z(product[9]) );
  NAND2_X1 U457 ( .A1(n504), .A2(n90), .ZN(n517) );
  XOR2_X1 U458 ( .A(n588), .B(a[2]), .Z(n518) );
  BUF_X2 U459 ( .A(n518), .Z(n519) );
  BUF_X2 U460 ( .A(n518), .Z(n520) );
  INV_X1 U461 ( .A(n570), .ZN(n21) );
  INV_X2 U462 ( .A(n593), .ZN(n592) );
  INV_X1 U463 ( .A(n524), .ZN(n521) );
  XNOR2_X1 U464 ( .A(n596), .B(a[10]), .ZN(n522) );
  BUF_X2 U465 ( .A(n518), .Z(n582) );
  INV_X1 U466 ( .A(n592), .ZN(n523) );
  CLKBUF_X1 U467 ( .A(n587), .Z(n525) );
  CLKBUF_X1 U468 ( .A(n16), .Z(n526) );
  CLKBUF_X1 U469 ( .A(n104), .Z(n527) );
  XNOR2_X1 U470 ( .A(n598), .B(a[12]), .ZN(n528) );
  INV_X1 U471 ( .A(n598), .ZN(n597) );
  INV_X1 U472 ( .A(n589), .ZN(n529) );
  CLKBUF_X1 U473 ( .A(n107), .Z(n530) );
  CLKBUF_X1 U474 ( .A(n569), .Z(n531) );
  XNOR2_X1 U475 ( .A(n598), .B(a[10]), .ZN(n428) );
  XNOR2_X1 U476 ( .A(n149), .B(n532), .ZN(n144) );
  XNOR2_X1 U477 ( .A(n271), .B(n146), .ZN(n532) );
  XNOR2_X1 U478 ( .A(n588), .B(n249), .ZN(n433) );
  CLKBUF_X1 U479 ( .A(n12), .Z(n533) );
  BUF_X1 U480 ( .A(n12), .Z(n534) );
  NAND2_X1 U481 ( .A1(n9), .A2(n568), .ZN(n12) );
  INV_X1 U482 ( .A(n594), .ZN(n536) );
  INV_X1 U483 ( .A(n594), .ZN(n537) );
  INV_X1 U484 ( .A(n559), .ZN(n538) );
  INV_X1 U485 ( .A(n522), .ZN(n539) );
  XOR2_X1 U486 ( .A(n596), .B(a[10]), .Z(n32) );
  XOR2_X1 U487 ( .A(n219), .B(n216), .Z(n540) );
  XOR2_X1 U488 ( .A(n214), .B(n540), .Z(n212) );
  NAND2_X1 U489 ( .A1(n214), .A2(n219), .ZN(n541) );
  NAND2_X1 U490 ( .A1(n214), .A2(n216), .ZN(n542) );
  NAND2_X1 U491 ( .A1(n219), .A2(n216), .ZN(n543) );
  NAND3_X1 U492 ( .A1(n541), .A2(n542), .A3(n543), .ZN(n211) );
  OR2_X1 U493 ( .A1(n228), .A2(n231), .ZN(n544) );
  XNOR2_X1 U494 ( .A(n593), .B(a[4]), .ZN(n567) );
  XOR2_X1 U495 ( .A(n588), .B(a[2]), .Z(n9) );
  XNOR2_X1 U496 ( .A(n596), .B(a[8]), .ZN(n429) );
  INV_X1 U497 ( .A(n596), .ZN(n595) );
  XNOR2_X1 U498 ( .A(n166), .B(n545), .ZN(n164) );
  XNOR2_X1 U499 ( .A(n177), .B(n168), .ZN(n545) );
  XNOR2_X1 U500 ( .A(n569), .B(n546), .ZN(product[12]) );
  AND2_X1 U501 ( .A1(n552), .A2(n79), .ZN(n546) );
  OR2_X1 U502 ( .A1(n196), .A2(n203), .ZN(n547) );
  NAND2_X1 U503 ( .A1(n166), .A2(n177), .ZN(n548) );
  NAND2_X1 U504 ( .A1(n166), .A2(n168), .ZN(n549) );
  NAND2_X1 U505 ( .A1(n177), .A2(n168), .ZN(n550) );
  NAND3_X1 U506 ( .A1(n548), .A2(n549), .A3(n550), .ZN(n163) );
  NAND2_X1 U507 ( .A1(n428), .A2(n32), .ZN(n551) );
  OR2_X1 U508 ( .A1(n176), .A2(n185), .ZN(n552) );
  NOR2_X1 U509 ( .A1(n164), .A2(n175), .ZN(n553) );
  INV_X1 U510 ( .A(n537), .ZN(n554) );
  CLKBUF_X2 U511 ( .A(n16), .Z(n581) );
  OR2_X2 U512 ( .A1(n555), .A2(n570), .ZN(n23) );
  XNOR2_X1 U513 ( .A(n19), .B(a[6]), .ZN(n555) );
  BUF_X1 U514 ( .A(n83), .Z(n556) );
  NOR2_X1 U515 ( .A1(n186), .A2(n195), .ZN(n558) );
  NOR2_X1 U516 ( .A1(n186), .A2(n195), .ZN(n82) );
  XNOR2_X1 U517 ( .A(n591), .B(a[2]), .ZN(n568) );
  INV_X1 U518 ( .A(n591), .ZN(n589) );
  XNOR2_X1 U519 ( .A(n594), .B(a[8]), .ZN(n559) );
  OAI21_X1 U520 ( .B1(n512), .B2(n89), .A(n90), .ZN(n560) );
  NAND2_X2 U521 ( .A1(n429), .A2(n506), .ZN(n29) );
  XOR2_X1 U522 ( .A(n591), .B(a[4]), .Z(n16) );
  XOR2_X1 U523 ( .A(n229), .B(n298), .Z(n561) );
  XOR2_X1 U524 ( .A(n226), .B(n561), .Z(n224) );
  NAND2_X1 U525 ( .A1(n226), .A2(n229), .ZN(n562) );
  NAND2_X1 U526 ( .A1(n226), .A2(n298), .ZN(n563) );
  NAND2_X1 U527 ( .A1(n229), .A2(n298), .ZN(n564) );
  NAND3_X1 U528 ( .A1(n562), .A2(n563), .A3(n564), .ZN(n223) );
  INV_X2 U529 ( .A(n588), .ZN(n587) );
  INV_X2 U530 ( .A(n249), .ZN(n586) );
  NAND2_X1 U531 ( .A1(n433), .A2(n586), .ZN(n565) );
  NAND2_X1 U532 ( .A1(n433), .A2(n586), .ZN(n566) );
  BUF_X1 U533 ( .A(n43), .Z(n584) );
  AOI21_X1 U534 ( .B1(n80), .B2(n560), .A(n81), .ZN(n569) );
  XNOR2_X1 U535 ( .A(n593), .B(a[6]), .ZN(n570) );
  AOI21_X1 U536 ( .B1(n505), .B2(n571), .A(n67), .ZN(n65) );
  INV_X1 U537 ( .A(n69), .ZN(n67) );
  NAND2_X1 U538 ( .A1(n571), .A2(n69), .ZN(n47) );
  INV_X1 U539 ( .A(n73), .ZN(n71) );
  NAND2_X1 U540 ( .A1(n73), .A2(n571), .ZN(n64) );
  INV_X1 U541 ( .A(n74), .ZN(n72) );
  INV_X1 U542 ( .A(n95), .ZN(n93) );
  AOI21_X1 U543 ( .B1(n560), .B2(n80), .A(n81), .ZN(n45) );
  OAI21_X1 U544 ( .B1(n91), .B2(n89), .A(n90), .ZN(n88) );
  NAND2_X1 U545 ( .A1(n127), .A2(n556), .ZN(n50) );
  NAND2_X1 U546 ( .A1(n572), .A2(n95), .ZN(n53) );
  OAI21_X1 U547 ( .B1(n553), .B2(n79), .A(n76), .ZN(n74) );
  NAND2_X1 U548 ( .A1(n502), .A2(n76), .ZN(n48) );
  NOR2_X1 U549 ( .A1(n553), .A2(n78), .ZN(n73) );
  NAND2_X1 U550 ( .A1(n152), .A2(n163), .ZN(n69) );
  NAND2_X1 U551 ( .A1(n131), .A2(n98), .ZN(n54) );
  INV_X1 U552 ( .A(n97), .ZN(n131) );
  NAND2_X1 U553 ( .A1(n135), .A2(n114), .ZN(n58) );
  NAND2_X1 U554 ( .A1(n544), .A2(n106), .ZN(n56) );
  AOI21_X1 U555 ( .B1(n575), .B2(n112), .A(n109), .ZN(n107) );
  INV_X1 U556 ( .A(n111), .ZN(n109) );
  NOR2_X1 U557 ( .A1(n176), .A2(n185), .ZN(n78) );
  AOI21_X1 U558 ( .B1(n573), .B2(n120), .A(n117), .ZN(n115) );
  INV_X1 U559 ( .A(n119), .ZN(n117) );
  INV_X1 U560 ( .A(n122), .ZN(n120) );
  NOR2_X1 U561 ( .A1(n196), .A2(n203), .ZN(n85) );
  XNOR2_X1 U562 ( .A(n57), .B(n112), .ZN(product[4]) );
  NAND2_X1 U563 ( .A1(n575), .A2(n111), .ZN(n57) );
  NAND2_X1 U564 ( .A1(n176), .A2(n185), .ZN(n79) );
  NAND2_X1 U565 ( .A1(n164), .A2(n175), .ZN(n76) );
  NAND2_X1 U566 ( .A1(n212), .A2(n217), .ZN(n95) );
  OR2_X1 U567 ( .A1(n212), .A2(n217), .ZN(n572) );
  NAND2_X1 U568 ( .A1(n196), .A2(n203), .ZN(n86) );
  XNOR2_X1 U569 ( .A(n59), .B(n120), .ZN(product[2]) );
  NAND2_X1 U570 ( .A1(n573), .A2(n119), .ZN(n59) );
  OR2_X1 U571 ( .A1(n328), .A2(n314), .ZN(n573) );
  OR2_X1 U572 ( .A1(n139), .A2(n151), .ZN(n574) );
  XNOR2_X1 U573 ( .A(n63), .B(n46), .ZN(product[15]) );
  NAND2_X1 U574 ( .A1(n574), .A2(n62), .ZN(n46) );
  NOR2_X1 U575 ( .A1(n218), .A2(n223), .ZN(n97) );
  OR2_X1 U576 ( .A1(n232), .A2(n233), .ZN(n575) );
  NAND2_X1 U577 ( .A1(n218), .A2(n223), .ZN(n98) );
  NAND2_X1 U578 ( .A1(n228), .A2(n231), .ZN(n106) );
  OR2_X1 U579 ( .A1(n224), .A2(n227), .ZN(n576) );
  INV_X1 U580 ( .A(n41), .ZN(n235) );
  AND2_X1 U581 ( .A1(n503), .A2(n122), .ZN(product[1]) );
  OR2_X1 U582 ( .A1(n584), .A2(n529), .ZN(n392) );
  AND2_X1 U583 ( .A1(n585), .A2(n245), .ZN(n300) );
  AND2_X1 U584 ( .A1(n585), .A2(n570), .ZN(n288) );
  AND2_X1 U585 ( .A1(n585), .A2(n522), .ZN(n270) );
  XNOR2_X1 U586 ( .A(n595), .B(n584), .ZN(n352) );
  OR2_X1 U587 ( .A1(n584), .A2(n600), .ZN(n337) );
  OAI22_X1 U588 ( .A1(n42), .A2(n602), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U589 ( .A1(n584), .A2(n602), .ZN(n332) );
  XNOR2_X1 U590 ( .A(n597), .B(n584), .ZN(n343) );
  NAND2_X1 U591 ( .A1(n433), .A2(n586), .ZN(n6) );
  XNOR2_X1 U592 ( .A(n155), .B(n578), .ZN(n139) );
  XNOR2_X1 U593 ( .A(n153), .B(n141), .ZN(n578) );
  XNOR2_X1 U594 ( .A(n157), .B(n579), .ZN(n141) );
  XNOR2_X1 U595 ( .A(n145), .B(n143), .ZN(n579) );
  XNOR2_X1 U596 ( .A(n159), .B(n580), .ZN(n142) );
  XNOR2_X1 U597 ( .A(n315), .B(n261), .ZN(n580) );
  XNOR2_X1 U598 ( .A(n592), .B(n584), .ZN(n376) );
  XNOR2_X1 U599 ( .A(n599), .B(n584), .ZN(n336) );
  NAND2_X1 U600 ( .A1(n427), .A2(n37), .ZN(n39) );
  XOR2_X1 U601 ( .A(n599), .B(a[12]), .Z(n427) );
  OAI22_X1 U602 ( .A1(n39), .A2(n336), .B1(n513), .B2(n335), .ZN(n263) );
  AND2_X1 U603 ( .A1(n585), .A2(n528), .ZN(n264) );
  AND2_X1 U604 ( .A1(n585), .A2(n235), .ZN(n260) );
  OAI22_X1 U605 ( .A1(n39), .A2(n335), .B1(n513), .B2(n334), .ZN(n262) );
  INV_X1 U606 ( .A(n19), .ZN(n594) );
  INV_X1 U607 ( .A(n25), .ZN(n596) );
  AND2_X1 U608 ( .A1(n585), .A2(n559), .ZN(n278) );
  INV_X1 U609 ( .A(n1), .ZN(n588) );
  NAND2_X1 U610 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U611 ( .A(n601), .B(a[14]), .Z(n426) );
  INV_X1 U612 ( .A(n7), .ZN(n591) );
  XNOR2_X1 U613 ( .A(n537), .B(n584), .ZN(n363) );
  AND2_X1 U614 ( .A1(n585), .A2(n247), .ZN(n314) );
  AND2_X1 U615 ( .A1(n585), .A2(n249), .ZN(product[0]) );
  OR2_X1 U616 ( .A1(n584), .A2(n554), .ZN(n364) );
  OR2_X1 U617 ( .A1(n584), .A2(n598), .ZN(n344) );
  OR2_X1 U618 ( .A1(n584), .A2(n596), .ZN(n353) );
  OR2_X1 U619 ( .A1(n584), .A2(n523), .ZN(n377) );
  XNOR2_X1 U620 ( .A(n537), .B(b[9]), .ZN(n354) );
  OAI22_X1 U621 ( .A1(n39), .A2(n334), .B1(n513), .B2(n333), .ZN(n261) );
  XNOR2_X1 U622 ( .A(n599), .B(n422), .ZN(n333) );
  XNOR2_X1 U623 ( .A(n592), .B(b[11]), .ZN(n365) );
  XNOR2_X1 U624 ( .A(n599), .B(n424), .ZN(n335) );
  XNOR2_X1 U625 ( .A(n599), .B(n423), .ZN(n334) );
  OAI22_X1 U626 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U627 ( .A(n601), .B(n424), .ZN(n330) );
  XNOR2_X1 U628 ( .A(n601), .B(n584), .ZN(n331) );
  XNOR2_X1 U629 ( .A(n510), .B(n418), .ZN(n345) );
  XNOR2_X1 U630 ( .A(n597), .B(n420), .ZN(n338) );
  XNOR2_X1 U631 ( .A(n490), .B(b[13]), .ZN(n378) );
  XNOR2_X1 U632 ( .A(n597), .B(n424), .ZN(n342) );
  XNOR2_X1 U633 ( .A(n536), .B(n424), .ZN(n362) );
  XNOR2_X1 U634 ( .A(n595), .B(n424), .ZN(n351) );
  XNOR2_X1 U635 ( .A(n597), .B(n423), .ZN(n341) );
  XNOR2_X1 U636 ( .A(n597), .B(n422), .ZN(n340) );
  XNOR2_X1 U637 ( .A(n597), .B(n421), .ZN(n339) );
  XNOR2_X1 U638 ( .A(n590), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U639 ( .A(n590), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U640 ( .A(n590), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U641 ( .A(n590), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U642 ( .A(n590), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U643 ( .A(n590), .B(n418), .ZN(n384) );
  XNOR2_X1 U644 ( .A(n590), .B(n419), .ZN(n385) );
  XNOR2_X1 U645 ( .A(n536), .B(n423), .ZN(n361) );
  XNOR2_X1 U646 ( .A(n510), .B(n423), .ZN(n350) );
  XNOR2_X1 U647 ( .A(n595), .B(n422), .ZN(n349) );
  XNOR2_X1 U648 ( .A(n537), .B(n422), .ZN(n360) );
  XNOR2_X1 U649 ( .A(n592), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U650 ( .A(n592), .B(n418), .ZN(n369) );
  XNOR2_X1 U651 ( .A(n592), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U652 ( .A(n592), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U653 ( .A(n536), .B(n420), .ZN(n358) );
  XNOR2_X1 U654 ( .A(n510), .B(n420), .ZN(n347) );
  XNOR2_X1 U655 ( .A(n536), .B(n418), .ZN(n356) );
  XNOR2_X1 U656 ( .A(n521), .B(b[11]), .ZN(n397) );
  XNOR2_X1 U657 ( .A(n525), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U658 ( .A(n508), .B(b[13]), .ZN(n395) );
  XNOR2_X1 U659 ( .A(n508), .B(b[14]), .ZN(n394) );
  XNOR2_X1 U660 ( .A(n537), .B(n421), .ZN(n359) );
  XNOR2_X1 U661 ( .A(n595), .B(n421), .ZN(n348) );
  XNOR2_X1 U662 ( .A(n536), .B(n419), .ZN(n357) );
  XNOR2_X1 U663 ( .A(n510), .B(n419), .ZN(n346) );
  XNOR2_X1 U664 ( .A(n536), .B(b[8]), .ZN(n355) );
  BUF_X1 U665 ( .A(n43), .Z(n585) );
  XNOR2_X1 U666 ( .A(n508), .B(b[15]), .ZN(n393) );
  OAI22_X1 U667 ( .A1(n551), .A2(n339), .B1(n338), .B2(n539), .ZN(n265) );
  OAI22_X1 U668 ( .A1(n551), .A2(n340), .B1(n339), .B2(n539), .ZN(n266) );
  OAI22_X1 U669 ( .A1(n551), .A2(n341), .B1(n340), .B2(n539), .ZN(n267) );
  OAI22_X1 U670 ( .A1(n551), .A2(n342), .B1(n341), .B2(n539), .ZN(n268) );
  OAI22_X1 U671 ( .A1(n551), .A2(n343), .B1(n342), .B2(n539), .ZN(n269) );
  OAI22_X1 U672 ( .A1(n551), .A2(n598), .B1(n344), .B2(n539), .ZN(n253) );
  INV_X1 U673 ( .A(n558), .ZN(n127) );
  NOR2_X1 U674 ( .A1(n558), .A2(n85), .ZN(n80) );
  OAI21_X1 U675 ( .B1(n82), .B2(n86), .A(n83), .ZN(n81) );
  NAND2_X1 U676 ( .A1(n186), .A2(n195), .ZN(n83) );
  INV_X1 U677 ( .A(n13), .ZN(n593) );
  NAND2_X1 U678 ( .A1(n232), .A2(n233), .ZN(n111) );
  NAND2_X1 U679 ( .A1(n576), .A2(n103), .ZN(n55) );
  INV_X1 U680 ( .A(n103), .ZN(n101) );
  NAND2_X1 U681 ( .A1(n224), .A2(n227), .ZN(n103) );
  XNOR2_X1 U682 ( .A(n84), .B(n50), .ZN(product[11]) );
  NOR2_X1 U683 ( .A1(n228), .A2(n231), .ZN(n105) );
  NAND2_X1 U684 ( .A1(n204), .A2(n211), .ZN(n90) );
  NOR2_X1 U685 ( .A1(n204), .A2(n211), .ZN(n89) );
  OAI22_X1 U686 ( .A1(n29), .A2(n350), .B1(n349), .B2(n538), .ZN(n275) );
  OAI22_X1 U687 ( .A1(n29), .A2(n346), .B1(n345), .B2(n538), .ZN(n271) );
  OAI22_X1 U688 ( .A1(n29), .A2(n347), .B1(n346), .B2(n538), .ZN(n272) );
  OAI22_X1 U689 ( .A1(n29), .A2(n348), .B1(n347), .B2(n538), .ZN(n273) );
  OAI22_X1 U690 ( .A1(n29), .A2(n349), .B1(n348), .B2(n538), .ZN(n274) );
  OAI22_X1 U691 ( .A1(n29), .A2(n596), .B1(n353), .B2(n538), .ZN(n254) );
  OAI22_X1 U692 ( .A1(n29), .A2(n351), .B1(n350), .B2(n538), .ZN(n276) );
  OAI22_X1 U693 ( .A1(n29), .A2(n352), .B1(n351), .B2(n538), .ZN(n277) );
  OAI21_X1 U694 ( .B1(n113), .B2(n115), .A(n114), .ZN(n112) );
  INV_X1 U695 ( .A(n113), .ZN(n135) );
  XNOR2_X1 U696 ( .A(n77), .B(n48), .ZN(product[13]) );
  XNOR2_X1 U697 ( .A(n589), .B(n420), .ZN(n386) );
  XNOR2_X1 U698 ( .A(n589), .B(n584), .ZN(n391) );
  XNOR2_X1 U699 ( .A(n589), .B(n423), .ZN(n389) );
  XNOR2_X1 U700 ( .A(n589), .B(n424), .ZN(n390) );
  XNOR2_X1 U701 ( .A(n589), .B(n422), .ZN(n388) );
  XNOR2_X1 U702 ( .A(n589), .B(n421), .ZN(n387) );
  CLKBUF_X1 U703 ( .A(n99), .Z(n583) );
  AOI21_X1 U704 ( .B1(n104), .B2(n576), .A(n101), .ZN(n99) );
  OAI21_X1 U705 ( .B1(n87), .B2(n85), .A(n501), .ZN(n84) );
  XNOR2_X1 U706 ( .A(n557), .B(n53), .ZN(product[8]) );
  XOR2_X1 U707 ( .A(n583), .B(n54), .Z(product[7]) );
  AOI21_X1 U708 ( .B1(n96), .B2(n572), .A(n93), .ZN(n91) );
  OR2_X1 U709 ( .A1(n584), .A2(n524), .ZN(n409) );
  XNOR2_X1 U710 ( .A(n70), .B(n47), .ZN(product[14]) );
  OAI22_X1 U711 ( .A1(n23), .A2(n358), .B1(n357), .B2(n21), .ZN(n282) );
  OAI22_X1 U712 ( .A1(n23), .A2(n356), .B1(n355), .B2(n21), .ZN(n280) );
  OAI22_X1 U713 ( .A1(n23), .A2(n362), .B1(n361), .B2(n21), .ZN(n286) );
  OAI22_X1 U714 ( .A1(n23), .A2(n360), .B1(n359), .B2(n21), .ZN(n284) );
  OAI22_X1 U715 ( .A1(n23), .A2(n554), .B1(n364), .B2(n21), .ZN(n255) );
  OAI22_X1 U716 ( .A1(n23), .A2(n361), .B1(n360), .B2(n21), .ZN(n285) );
  OAI22_X1 U717 ( .A1(n23), .A2(n357), .B1(n356), .B2(n21), .ZN(n281) );
  OAI22_X1 U718 ( .A1(n23), .A2(n355), .B1(n354), .B2(n21), .ZN(n279) );
  XNOR2_X1 U719 ( .A(n592), .B(n424), .ZN(n375) );
  OAI22_X1 U720 ( .A1(n23), .A2(n363), .B1(n362), .B2(n21), .ZN(n287) );
  XNOR2_X1 U721 ( .A(n592), .B(n423), .ZN(n374) );
  XNOR2_X1 U722 ( .A(n592), .B(n421), .ZN(n372) );
  OAI22_X1 U723 ( .A1(n23), .A2(n359), .B1(n358), .B2(n21), .ZN(n283) );
  XNOR2_X1 U724 ( .A(n592), .B(n422), .ZN(n373) );
  XNOR2_X1 U725 ( .A(n592), .B(n419), .ZN(n370) );
  XNOR2_X1 U726 ( .A(n592), .B(n420), .ZN(n371) );
  INV_X1 U727 ( .A(n88), .ZN(n87) );
  XNOR2_X1 U728 ( .A(n587), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U729 ( .A(n587), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U730 ( .A(n587), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U731 ( .A(n587), .B(n418), .ZN(n401) );
  XNOR2_X1 U732 ( .A(n521), .B(n423), .ZN(n406) );
  XNOR2_X1 U733 ( .A(n521), .B(n584), .ZN(n408) );
  XNOR2_X1 U734 ( .A(n587), .B(n422), .ZN(n405) );
  XNOR2_X1 U735 ( .A(n587), .B(n421), .ZN(n404) );
  XNOR2_X1 U736 ( .A(n587), .B(n420), .ZN(n403) );
  XNOR2_X1 U737 ( .A(n587), .B(n424), .ZN(n407) );
  XNOR2_X1 U738 ( .A(n587), .B(n419), .ZN(n402) );
  NAND2_X1 U739 ( .A1(n151), .A2(n139), .ZN(n62) );
  OAI22_X1 U740 ( .A1(n492), .A2(n370), .B1(n369), .B2(n581), .ZN(n293) );
  OAI22_X1 U741 ( .A1(n492), .A2(n367), .B1(n366), .B2(n581), .ZN(n290) );
  OAI22_X1 U742 ( .A1(n492), .A2(n375), .B1(n374), .B2(n581), .ZN(n298) );
  OAI22_X1 U743 ( .A1(n492), .A2(n368), .B1(n367), .B2(n581), .ZN(n291) );
  OAI22_X1 U744 ( .A1(n492), .A2(n373), .B1(n372), .B2(n581), .ZN(n296) );
  OAI22_X1 U745 ( .A1(n491), .A2(n369), .B1(n581), .B2(n368), .ZN(n292) );
  OAI22_X1 U746 ( .A1(n492), .A2(n523), .B1(n377), .B2(n581), .ZN(n256) );
  OAI22_X1 U747 ( .A1(n492), .A2(n372), .B1(n371), .B2(n581), .ZN(n295) );
  OAI22_X1 U748 ( .A1(n492), .A2(n371), .B1(n370), .B2(n581), .ZN(n294) );
  OAI22_X1 U749 ( .A1(n492), .A2(n376), .B1(n375), .B2(n581), .ZN(n299) );
  OAI22_X1 U750 ( .A1(n492), .A2(n374), .B1(n373), .B2(n581), .ZN(n297) );
  OAI22_X1 U751 ( .A1(n491), .A2(n366), .B1(n365), .B2(n581), .ZN(n289) );
  INV_X1 U752 ( .A(n526), .ZN(n245) );
  OAI21_X1 U753 ( .B1(n64), .B2(n531), .A(n65), .ZN(n63) );
  OAI21_X1 U754 ( .B1(n71), .B2(n45), .A(n72), .ZN(n70) );
  OAI21_X1 U755 ( .B1(n45), .B2(n78), .A(n79), .ZN(n77) );
  XNOR2_X1 U756 ( .A(n527), .B(n55), .ZN(product[6]) );
  NAND2_X1 U757 ( .A1(n328), .A2(n314), .ZN(n119) );
  OAI21_X1 U758 ( .B1(n105), .B2(n107), .A(n106), .ZN(n104) );
  NOR2_X1 U759 ( .A1(n234), .A2(n257), .ZN(n113) );
  XOR2_X1 U760 ( .A(n56), .B(n530), .Z(product[5]) );
  XOR2_X1 U761 ( .A(n58), .B(n115), .Z(product[3]) );
  OAI22_X1 U762 ( .A1(n566), .A2(n395), .B1(n394), .B2(n586), .ZN(n316) );
  OAI22_X1 U763 ( .A1(n6), .A2(n394), .B1(n393), .B2(n586), .ZN(n315) );
  OAI22_X1 U764 ( .A1(n565), .A2(n396), .B1(n395), .B2(n586), .ZN(n317) );
  OAI22_X1 U765 ( .A1(n6), .A2(n397), .B1(n396), .B2(n586), .ZN(n318) );
  OAI22_X1 U766 ( .A1(n565), .A2(n398), .B1(n397), .B2(n586), .ZN(n319) );
  OAI22_X1 U767 ( .A1(n6), .A2(n400), .B1(n399), .B2(n586), .ZN(n321) );
  OAI22_X1 U768 ( .A1(n565), .A2(n399), .B1(n398), .B2(n586), .ZN(n320) );
  OAI22_X1 U769 ( .A1(n566), .A2(n401), .B1(n400), .B2(n586), .ZN(n322) );
  OAI22_X1 U770 ( .A1(n6), .A2(n402), .B1(n401), .B2(n586), .ZN(n323) );
  NAND2_X1 U771 ( .A1(n329), .A2(n258), .ZN(n122) );
  OAI22_X1 U772 ( .A1(n565), .A2(n404), .B1(n403), .B2(n586), .ZN(n325) );
  OAI22_X1 U773 ( .A1(n6), .A2(n403), .B1(n402), .B2(n586), .ZN(n324) );
  OAI22_X1 U774 ( .A1(n566), .A2(n406), .B1(n405), .B2(n586), .ZN(n327) );
  OAI22_X1 U775 ( .A1(n566), .A2(n405), .B1(n404), .B2(n586), .ZN(n326) );
  OAI22_X1 U776 ( .A1(n566), .A2(n407), .B1(n406), .B2(n586), .ZN(n328) );
  OAI22_X1 U777 ( .A1(n6), .A2(n408), .B1(n407), .B2(n586), .ZN(n329) );
  OAI22_X1 U778 ( .A1(n565), .A2(n524), .B1(n409), .B2(n586), .ZN(n258) );
  OAI22_X1 U779 ( .A1(n509), .A2(n379), .B1(n378), .B2(n520), .ZN(n301) );
  OAI22_X1 U780 ( .A1(n509), .A2(n380), .B1(n379), .B2(n520), .ZN(n302) );
  OAI22_X1 U781 ( .A1(n533), .A2(n385), .B1(n384), .B2(n519), .ZN(n307) );
  OAI22_X1 U782 ( .A1(n509), .A2(n382), .B1(n381), .B2(n582), .ZN(n304) );
  OAI22_X1 U783 ( .A1(n535), .A2(n381), .B1(n380), .B2(n519), .ZN(n303) );
  NAND2_X1 U784 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U785 ( .A1(n534), .A2(n383), .B1(n382), .B2(n519), .ZN(n305) );
  OAI22_X1 U786 ( .A1(n534), .A2(n384), .B1(n383), .B2(n520), .ZN(n306) );
  OAI22_X1 U787 ( .A1(n533), .A2(n386), .B1(n385), .B2(n519), .ZN(n308) );
  OAI22_X1 U788 ( .A1(n509), .A2(n387), .B1(n386), .B2(n582), .ZN(n309) );
  OAI22_X1 U789 ( .A1(n535), .A2(n529), .B1(n392), .B2(n582), .ZN(n257) );
  OAI22_X1 U790 ( .A1(n534), .A2(n389), .B1(n582), .B2(n388), .ZN(n311) );
  OAI22_X1 U791 ( .A1(n535), .A2(n388), .B1(n387), .B2(n582), .ZN(n310) );
  OAI22_X1 U792 ( .A1(n535), .A2(n390), .B1(n389), .B2(n519), .ZN(n312) );
  INV_X1 U793 ( .A(n520), .ZN(n247) );
  OAI22_X1 U794 ( .A1(n533), .A2(n391), .B1(n390), .B2(n520), .ZN(n313) );
  INV_X1 U795 ( .A(n591), .ZN(n590) );
  INV_X1 U796 ( .A(n31), .ZN(n598) );
  INV_X1 U797 ( .A(n36), .ZN(n600) );
  INV_X1 U798 ( .A(n602), .ZN(n601) );
  INV_X1 U799 ( .A(n40), .ZN(n602) );
  XOR2_X1 U800 ( .A(n259), .B(n251), .Z(n148) );
  XOR2_X1 U801 ( .A(n289), .B(n279), .Z(n146) );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_11_DW01_add_2 ( A, B, CI, 
        SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n8, n9, n10, n11, n12, n13, n14, n15, n16, n19,
         n20, n22, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n44, n45, n47, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n65, n67, n68, n69, n70,
         n71, n73, n75, n76, n77, n78, n79, n81, n83, n84, n86, n88, n89, n90,
         n91, n94, n95, n96, n98, n100, n157, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179;

  BUF_X1 U122 ( .A(n168), .Z(n157) );
  AND2_X1 U123 ( .A1(n172), .A2(n86), .ZN(SUM[0]) );
  BUF_X1 U124 ( .A(n55), .Z(n159) );
  XNOR2_X1 U125 ( .A(n45), .B(n160), .ZN(SUM[10]) );
  AND2_X1 U126 ( .A1(n44), .A2(n166), .ZN(n160) );
  BUF_X1 U127 ( .A(n36), .Z(n168) );
  BUF_X1 U128 ( .A(n29), .Z(n162) );
  XNOR2_X1 U129 ( .A(n38), .B(n6), .ZN(SUM[11]) );
  NOR2_X1 U130 ( .A1(A[11]), .A2(B[11]), .ZN(n35) );
  OR2_X1 U131 ( .A1(A[15]), .A2(B[15]), .ZN(n161) );
  BUF_X1 U132 ( .A(n26), .Z(n163) );
  NOR2_X1 U133 ( .A1(A[8]), .A2(B[8]), .ZN(n164) );
  CLKBUF_X1 U134 ( .A(n179), .Z(n165) );
  OR2_X1 U135 ( .A1(A[10]), .A2(B[10]), .ZN(n166) );
  OR2_X1 U136 ( .A1(A[10]), .A2(B[10]), .ZN(n178) );
  NOR2_X1 U137 ( .A1(A[12]), .A2(B[12]), .ZN(n167) );
  NOR2_X1 U138 ( .A1(A[12]), .A2(B[12]), .ZN(n32) );
  NOR2_X1 U139 ( .A1(A[14]), .A2(B[14]), .ZN(n169) );
  NOR2_X1 U140 ( .A1(A[14]), .A2(B[14]), .ZN(n25) );
  AOI21_X1 U141 ( .B1(n38), .B2(n30), .A(n31), .ZN(n170) );
  AOI21_X1 U142 ( .B1(n38), .B2(n30), .A(n31), .ZN(n171) );
  OR2_X1 U143 ( .A1(A[0]), .A2(B[0]), .ZN(n172) );
  INV_X1 U144 ( .A(n60), .ZN(n59) );
  INV_X1 U145 ( .A(n51), .ZN(n50) );
  OAI21_X1 U146 ( .B1(n71), .B2(n69), .A(n70), .ZN(n68) );
  OAI21_X1 U147 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  AOI21_X1 U148 ( .B1(n176), .B2(n84), .A(n81), .ZN(n79) );
  INV_X1 U149 ( .A(n83), .ZN(n81) );
  OAI21_X1 U150 ( .B1(n79), .B2(n77), .A(n78), .ZN(n76) );
  NAND2_X1 U151 ( .A1(n89), .A2(n162), .ZN(n4) );
  INV_X1 U152 ( .A(n28), .ZN(n89) );
  OR2_X1 U153 ( .A1(n169), .A2(n28), .ZN(n173) );
  AOI21_X1 U154 ( .B1(n177), .B2(n68), .A(n65), .ZN(n63) );
  INV_X1 U155 ( .A(n67), .ZN(n65) );
  AOI21_X1 U156 ( .B1(n175), .B2(n76), .A(n73), .ZN(n71) );
  INV_X1 U157 ( .A(n75), .ZN(n73) );
  AOI21_X1 U158 ( .B1(n52), .B2(n60), .A(n53), .ZN(n51) );
  AOI21_X1 U159 ( .B1(n50), .B2(n174), .A(n47), .ZN(n45) );
  NAND2_X1 U160 ( .A1(n94), .A2(n159), .ZN(n9) );
  INV_X1 U161 ( .A(n86), .ZN(n84) );
  OAI21_X1 U162 ( .B1(n59), .B2(n57), .A(n58), .ZN(n56) );
  INV_X1 U163 ( .A(n49), .ZN(n47) );
  NAND2_X1 U164 ( .A1(n95), .A2(n58), .ZN(n10) );
  INV_X1 U165 ( .A(n57), .ZN(n95) );
  NAND2_X1 U166 ( .A1(n96), .A2(n62), .ZN(n11) );
  INV_X1 U167 ( .A(n61), .ZN(n96) );
  NAND2_X1 U168 ( .A1(n174), .A2(n49), .ZN(n8) );
  NAND2_X1 U169 ( .A1(n177), .A2(n67), .ZN(n12) );
  NAND2_X1 U170 ( .A1(n100), .A2(n78), .ZN(n15) );
  INV_X1 U171 ( .A(n77), .ZN(n100) );
  NAND2_X1 U172 ( .A1(n175), .A2(n75), .ZN(n14) );
  NAND2_X1 U173 ( .A1(n176), .A2(n83), .ZN(n16) );
  NAND2_X1 U174 ( .A1(n98), .A2(n70), .ZN(n13) );
  INV_X1 U175 ( .A(n69), .ZN(n98) );
  NAND2_X1 U176 ( .A1(n88), .A2(n163), .ZN(n3) );
  NAND2_X1 U177 ( .A1(n91), .A2(n168), .ZN(n6) );
  NAND2_X1 U178 ( .A1(n90), .A2(n33), .ZN(n5) );
  XNOR2_X1 U179 ( .A(n50), .B(n8), .ZN(SUM[9]) );
  XOR2_X1 U180 ( .A(n59), .B(n10), .Z(SUM[7]) );
  XNOR2_X1 U181 ( .A(n14), .B(n76), .ZN(SUM[3]) );
  XOR2_X1 U182 ( .A(n15), .B(n79), .Z(SUM[2]) );
  NOR2_X1 U183 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  NOR2_X1 U184 ( .A1(A[7]), .A2(B[7]), .ZN(n57) );
  NOR2_X1 U185 ( .A1(A[8]), .A2(B[8]), .ZN(n54) );
  OR2_X1 U186 ( .A1(A[9]), .A2(B[9]), .ZN(n174) );
  NOR2_X1 U187 ( .A1(A[2]), .A2(B[2]), .ZN(n77) );
  NAND2_X1 U188 ( .A1(A[11]), .A2(B[11]), .ZN(n36) );
  OR2_X1 U189 ( .A1(A[3]), .A2(B[3]), .ZN(n175) );
  OR2_X1 U190 ( .A1(A[1]), .A2(B[1]), .ZN(n176) );
  OR2_X1 U191 ( .A1(A[5]), .A2(B[5]), .ZN(n177) );
  NOR2_X1 U192 ( .A1(A[4]), .A2(B[4]), .ZN(n69) );
  NOR2_X1 U193 ( .A1(A[6]), .A2(B[6]), .ZN(n61) );
  NAND2_X1 U194 ( .A1(A[14]), .A2(B[14]), .ZN(n26) );
  XNOR2_X1 U195 ( .A(n56), .B(n9), .ZN(SUM[8]) );
  XNOR2_X1 U196 ( .A(n16), .B(n84), .ZN(SUM[1]) );
  NAND2_X1 U197 ( .A1(A[7]), .A2(B[7]), .ZN(n58) );
  NAND2_X1 U198 ( .A1(A[2]), .A2(B[2]), .ZN(n78) );
  NAND2_X1 U199 ( .A1(A[1]), .A2(B[1]), .ZN(n83) );
  NAND2_X1 U200 ( .A1(A[3]), .A2(B[3]), .ZN(n75) );
  NAND2_X1 U201 ( .A1(A[0]), .A2(B[0]), .ZN(n86) );
  NAND2_X1 U202 ( .A1(A[4]), .A2(B[4]), .ZN(n70) );
  NAND2_X1 U203 ( .A1(A[6]), .A2(B[6]), .ZN(n62) );
  XNOR2_X1 U204 ( .A(n12), .B(n68), .ZN(SUM[5]) );
  NAND2_X1 U205 ( .A1(n161), .A2(n19), .ZN(n2) );
  INV_X1 U206 ( .A(n24), .ZN(n22) );
  INV_X1 U207 ( .A(n164), .ZN(n94) );
  NOR2_X1 U208 ( .A1(n164), .A2(n57), .ZN(n52) );
  OAI21_X1 U209 ( .B1(n54), .B2(n58), .A(n55), .ZN(n53) );
  NAND2_X1 U210 ( .A1(A[8]), .A2(B[8]), .ZN(n55) );
  INV_X1 U211 ( .A(n165), .ZN(n44) );
  AND2_X1 U212 ( .A1(A[10]), .A2(B[10]), .ZN(n179) );
  XOR2_X1 U213 ( .A(n11), .B(n63), .Z(SUM[6]) );
  NAND2_X1 U214 ( .A1(A[5]), .A2(B[5]), .ZN(n67) );
  NAND2_X1 U215 ( .A1(A[9]), .A2(B[9]), .ZN(n49) );
  XOR2_X1 U216 ( .A(n13), .B(n71), .Z(SUM[4]) );
  INV_X1 U217 ( .A(n167), .ZN(n90) );
  OAI21_X1 U218 ( .B1(n32), .B2(n36), .A(n33), .ZN(n31) );
  NAND2_X1 U219 ( .A1(A[13]), .A2(B[13]), .ZN(n29) );
  NAND2_X1 U220 ( .A1(A[15]), .A2(B[15]), .ZN(n19) );
  NAND2_X1 U221 ( .A1(A[12]), .A2(B[12]), .ZN(n33) );
  INV_X1 U222 ( .A(n38), .ZN(n37) );
  INV_X1 U223 ( .A(n169), .ZN(n88) );
  OAI21_X1 U224 ( .B1(n25), .B2(n29), .A(n26), .ZN(n24) );
  OAI21_X1 U225 ( .B1(n37), .B2(n35), .A(n157), .ZN(n34) );
  INV_X1 U226 ( .A(n35), .ZN(n91) );
  NOR2_X1 U227 ( .A1(n167), .A2(n35), .ZN(n30) );
  XNOR2_X1 U228 ( .A(n20), .B(n2), .ZN(SUM[15]) );
  OAI21_X1 U229 ( .B1(n39), .B2(n51), .A(n40), .ZN(n38) );
  NAND2_X1 U230 ( .A1(n166), .A2(n174), .ZN(n39) );
  AOI21_X1 U231 ( .B1(n178), .B2(n47), .A(n179), .ZN(n40) );
  XNOR2_X1 U232 ( .A(n34), .B(n5), .ZN(SUM[12]) );
  XNOR2_X1 U233 ( .A(n27), .B(n3), .ZN(SUM[14]) );
  XOR2_X1 U234 ( .A(n4), .B(n170), .Z(SUM[13]) );
  OAI21_X1 U235 ( .B1(n171), .B2(n173), .A(n22), .ZN(n20) );
  OAI21_X1 U236 ( .B1(n170), .B2(n28), .A(n162), .ZN(n27) );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_11 ( clk, clear_acc, 
        data_out_x, data_out, data_out_w, data_out_b, wr_en_y, m_valid, 
        m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [4:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
         N39, N40, N41, N42, N43, N44, n1, n2, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n85, n102, n111, n112, n113, n114, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n23), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n225), .CK(clk), .Q(n26) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n226), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n227), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n228), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n229), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n230), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n231), .CK(clk), .Q(n34) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n232), .CK(clk), .Q(n35) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n233), .CK(clk), .Q(n36) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n234), .CK(clk), .Q(n37) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n235), .CK(clk), .Q(n38) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n236), .CK(clk), .Q(n39) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n237), .CK(clk), .Q(n40) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n238), .CK(clk), .Q(n41) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n239), .CK(clk), .Q(n42) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n240), .CK(clk), .Q(n43) );
  DFF_X1 \f_reg[0]  ( .D(n113), .CK(clk), .Q(f[0]), .QN(n214) );
  DFF_X1 \f_reg[1]  ( .D(n112), .CK(clk), .Q(f[1]), .QN(n215) );
  DFF_X1 \f_reg[2]  ( .D(n111), .CK(clk), .Q(f[2]), .QN(n216) );
  DFF_X1 \f_reg[7]  ( .D(n81), .CK(clk), .Q(f[7]), .QN(n217) );
  DFF_X1 \f_reg[8]  ( .D(n80), .CK(clk), .Q(f[8]), .QN(n218) );
  DFF_X1 \f_reg[9]  ( .D(n79), .CK(clk), .Q(f[9]), .QN(n219) );
  DFF_X1 \f_reg[10]  ( .D(n78), .CK(clk), .Q(n52), .QN(n220) );
  DFF_X1 \f_reg[11]  ( .D(n77), .CK(clk), .Q(n50), .QN(n221) );
  DFF_X1 \f_reg[12]  ( .D(n4), .CK(clk), .Q(n49), .QN(n222) );
  DFF_X1 \f_reg[13]  ( .D(n18), .CK(clk), .Q(n48), .QN(n223) );
  DFF_X1 \f_reg[14]  ( .D(n6), .CK(clk), .Q(n47), .QN(n224) );
  DFF_X1 \data_out_reg[15]  ( .D(n166), .CK(clk), .Q(data_out[15]), .QN(n197)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n167), .CK(clk), .Q(data_out[14]), .QN(n196)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n168), .CK(clk), .Q(data_out[13]), .QN(n195)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n169), .CK(clk), .Q(data_out[12]), .QN(n194)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n170), .CK(clk), .Q(data_out[11]), .QN(n193)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n171), .CK(clk), .Q(data_out[10]), .QN(n192)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n172), .CK(clk), .Q(data_out[9]), .QN(n191) );
  DFF_X1 \data_out_reg[8]  ( .D(n173), .CK(clk), .Q(data_out[8]), .QN(n190) );
  DFF_X1 \data_out_reg[7]  ( .D(n174), .CK(clk), .Q(data_out[7]), .QN(n189) );
  DFF_X1 \data_out_reg[6]  ( .D(n175), .CK(clk), .Q(data_out[6]), .QN(n188) );
  DFF_X1 \data_out_reg[5]  ( .D(n176), .CK(clk), .Q(data_out[5]), .QN(n187) );
  DFF_X1 \data_out_reg[4]  ( .D(n177), .CK(clk), .Q(data_out[4]), .QN(n186) );
  DFF_X1 \data_out_reg[3]  ( .D(n178), .CK(clk), .Q(data_out[3]), .QN(n185) );
  DFF_X1 \data_out_reg[2]  ( .D(n179), .CK(clk), .Q(data_out[2]), .QN(n184) );
  DFF_X1 \data_out_reg[1]  ( .D(n180), .CK(clk), .Q(data_out[1]), .QN(n183) );
  DFF_X1 \data_out_reg[0]  ( .D(n181), .CK(clk), .Q(data_out[0]), .QN(n182) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_11_DW_mult_tc_1 mult_2021 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_11_DW01_add_2 add_2022 ( .A({
        n204, n203, n202, n201, n200, n199, n213, n212, n211, n210, n209, n208, 
        n207, n206, n205, n198}), .B({f[15], n47, n48, n49, n50, n52, f[9:0]}), 
        .CI(1'b0), .SUM(adder) );
  DFF_X2 \f_reg[15]  ( .D(n76), .CK(clk), .Q(f[15]), .QN(n73) );
  DFF_X1 delay_reg ( .D(n114), .CK(clk), .Q(n13), .QN(n241) );
  DFF_X1 \f_reg[3]  ( .D(n102), .CK(clk), .Q(f[3]), .QN(n65) );
  DFF_X1 \f_reg[4]  ( .D(n85), .CK(clk), .Q(f[4]), .QN(n66) );
  DFF_X1 \f_reg[5]  ( .D(n83), .CK(clk), .Q(f[5]), .QN(n67) );
  DFF_X1 \f_reg[6]  ( .D(n82), .CK(clk), .Q(f[6]), .QN(n68) );
  CLKBUF_X1 U3 ( .A(N43), .Z(n1) );
  AND2_X1 U4 ( .A1(n46), .A2(n24), .ZN(n17) );
  AND2_X1 U5 ( .A1(clear_acc_delay), .A2(n241), .ZN(n2) );
  NAND3_X1 U6 ( .A1(n8), .A2(n7), .A3(n9), .ZN(n4) );
  CLKBUF_X1 U8 ( .A(N44), .Z(n5) );
  NAND3_X1 U9 ( .A1(n15), .A2(n14), .A3(n16), .ZN(n6) );
  NAND2_X1 U10 ( .A1(data_out_b[12]), .A2(n23), .ZN(n7) );
  NAND2_X1 U11 ( .A1(adder[12]), .A2(n17), .ZN(n8) );
  NAND2_X1 U12 ( .A1(n63), .A2(n49), .ZN(n9) );
  OAI222_X1 U13 ( .A1(n10), .A2(n24), .B1(n11), .B2(n12), .C1(n73), .C2(n46), 
        .ZN(n76) );
  INV_X1 U14 ( .A(data_out_b[15]), .ZN(n10) );
  INV_X1 U15 ( .A(adder[15]), .ZN(n11) );
  INV_X1 U16 ( .A(n17), .ZN(n12) );
  MUX2_X2 U17 ( .A(n35), .B(N37), .S(n241), .Z(n212) );
  MUX2_X2 U18 ( .A(n32), .B(N40), .S(n241), .Z(n200) );
  MUX2_X2 U19 ( .A(N39), .B(n33), .S(n13), .Z(n199) );
  MUX2_X2 U20 ( .A(n29), .B(N41), .S(n241), .Z(n201) );
  MUX2_X2 U21 ( .A(n27), .B(N43), .S(n241), .Z(n203) );
  NAND2_X1 U22 ( .A1(data_out_b[14]), .A2(n23), .ZN(n14) );
  NAND2_X1 U23 ( .A1(adder[14]), .A2(n17), .ZN(n15) );
  NAND2_X1 U24 ( .A1(n63), .A2(n47), .ZN(n16) );
  NAND2_X1 U25 ( .A1(n114), .A2(n22), .ZN(n243) );
  INV_X1 U26 ( .A(clear_acc), .ZN(n24) );
  OAI22_X1 U27 ( .A1(n185), .A2(n243), .B1(n65), .B2(n242), .ZN(n178) );
  OAI22_X1 U28 ( .A1(n186), .A2(n243), .B1(n66), .B2(n242), .ZN(n177) );
  OAI22_X1 U29 ( .A1(n187), .A2(n243), .B1(n67), .B2(n242), .ZN(n176) );
  OAI22_X1 U30 ( .A1(n188), .A2(n243), .B1(n68), .B2(n242), .ZN(n175) );
  OAI22_X1 U31 ( .A1(n189), .A2(n243), .B1(n217), .B2(n242), .ZN(n174) );
  OAI22_X1 U32 ( .A1(n190), .A2(n243), .B1(n218), .B2(n242), .ZN(n173) );
  OAI22_X1 U33 ( .A1(n191), .A2(n243), .B1(n219), .B2(n242), .ZN(n172) );
  NAND3_X1 U34 ( .A1(n20), .A2(n19), .A3(n21), .ZN(n18) );
  NAND2_X1 U35 ( .A1(data_out_b[13]), .A2(n23), .ZN(n19) );
  NAND2_X1 U36 ( .A1(adder[13]), .A2(n17), .ZN(n20) );
  NAND2_X1 U37 ( .A1(n63), .A2(n48), .ZN(n21) );
  INV_X1 U38 ( .A(n46), .ZN(n63) );
  INV_X1 U39 ( .A(wr_en_y), .ZN(n22) );
  INV_X1 U40 ( .A(n24), .ZN(n23) );
  INV_X1 U41 ( .A(m_ready), .ZN(n25) );
  NAND2_X1 U42 ( .A1(m_valid), .A2(n25), .ZN(n44) );
  OAI21_X1 U43 ( .B1(sel[4]), .B2(n75), .A(n44), .ZN(n114) );
  MUX2_X1 U44 ( .A(n26), .B(n5), .S(n2), .Z(n225) );
  MUX2_X1 U45 ( .A(n26), .B(N44), .S(n241), .Z(n204) );
  MUX2_X1 U46 ( .A(n27), .B(n1), .S(n2), .Z(n226) );
  MUX2_X1 U47 ( .A(n28), .B(N42), .S(n2), .Z(n227) );
  MUX2_X1 U48 ( .A(n28), .B(N42), .S(n241), .Z(n202) );
  MUX2_X1 U49 ( .A(n29), .B(N41), .S(n2), .Z(n228) );
  MUX2_X1 U50 ( .A(n32), .B(N40), .S(n2), .Z(n229) );
  MUX2_X1 U51 ( .A(n33), .B(N39), .S(n2), .Z(n230) );
  MUX2_X1 U52 ( .A(n34), .B(N38), .S(n2), .Z(n231) );
  MUX2_X1 U53 ( .A(n34), .B(N38), .S(n241), .Z(n213) );
  MUX2_X1 U54 ( .A(n35), .B(N37), .S(n2), .Z(n232) );
  MUX2_X1 U55 ( .A(n36), .B(N36), .S(n2), .Z(n233) );
  MUX2_X1 U56 ( .A(n36), .B(N36), .S(n241), .Z(n211) );
  MUX2_X1 U57 ( .A(n37), .B(N35), .S(n2), .Z(n234) );
  MUX2_X1 U58 ( .A(n37), .B(N35), .S(n241), .Z(n210) );
  MUX2_X1 U59 ( .A(n38), .B(N34), .S(n2), .Z(n235) );
  MUX2_X1 U60 ( .A(n38), .B(N34), .S(n241), .Z(n209) );
  MUX2_X1 U61 ( .A(n39), .B(N33), .S(n2), .Z(n236) );
  MUX2_X1 U62 ( .A(n39), .B(N33), .S(n241), .Z(n208) );
  MUX2_X1 U63 ( .A(n40), .B(N32), .S(n2), .Z(n237) );
  MUX2_X1 U64 ( .A(n40), .B(N32), .S(n241), .Z(n207) );
  MUX2_X1 U65 ( .A(n41), .B(N31), .S(n2), .Z(n238) );
  MUX2_X1 U66 ( .A(n41), .B(N31), .S(n241), .Z(n206) );
  MUX2_X1 U67 ( .A(n42), .B(N30), .S(n2), .Z(n239) );
  MUX2_X1 U68 ( .A(n42), .B(N30), .S(n241), .Z(n205) );
  MUX2_X1 U69 ( .A(n43), .B(N29), .S(n2), .Z(n240) );
  MUX2_X1 U70 ( .A(n43), .B(N29), .S(n241), .Z(n198) );
  INV_X1 U71 ( .A(n44), .ZN(n45) );
  OAI21_X1 U72 ( .B1(n45), .B2(n13), .A(n24), .ZN(n46) );
  AOI222_X1 U73 ( .A1(data_out_b[11]), .A2(n23), .B1(adder[11]), .B2(n17), 
        .C1(n63), .C2(n50), .ZN(n51) );
  INV_X1 U74 ( .A(n51), .ZN(n77) );
  AOI222_X1 U75 ( .A1(data_out_b[10]), .A2(n23), .B1(adder[10]), .B2(n17), 
        .C1(n63), .C2(n52), .ZN(n53) );
  INV_X1 U76 ( .A(n53), .ZN(n78) );
  AOI222_X1 U77 ( .A1(data_out_b[8]), .A2(n23), .B1(adder[8]), .B2(n17), .C1(
        n63), .C2(f[8]), .ZN(n54) );
  INV_X1 U78 ( .A(n54), .ZN(n80) );
  AOI222_X1 U79 ( .A1(data_out_b[7]), .A2(n23), .B1(adder[7]), .B2(n17), .C1(
        n63), .C2(f[7]), .ZN(n55) );
  INV_X1 U80 ( .A(n55), .ZN(n81) );
  AOI222_X1 U81 ( .A1(data_out_b[6]), .A2(n23), .B1(adder[6]), .B2(n17), .C1(
        n63), .C2(f[6]), .ZN(n56) );
  INV_X1 U82 ( .A(n56), .ZN(n82) );
  AOI222_X1 U83 ( .A1(data_out_b[5]), .A2(n23), .B1(adder[5]), .B2(n17), .C1(
        n63), .C2(f[5]), .ZN(n57) );
  INV_X1 U84 ( .A(n57), .ZN(n83) );
  AOI222_X1 U85 ( .A1(data_out_b[4]), .A2(n23), .B1(adder[4]), .B2(n17), .C1(
        n63), .C2(f[4]), .ZN(n58) );
  INV_X1 U86 ( .A(n58), .ZN(n85) );
  AOI222_X1 U87 ( .A1(data_out_b[3]), .A2(n23), .B1(adder[3]), .B2(n17), .C1(
        n63), .C2(f[3]), .ZN(n59) );
  INV_X1 U88 ( .A(n59), .ZN(n102) );
  AOI222_X1 U89 ( .A1(data_out_b[2]), .A2(n23), .B1(adder[2]), .B2(n17), .C1(
        n63), .C2(f[2]), .ZN(n60) );
  INV_X1 U90 ( .A(n60), .ZN(n111) );
  AOI222_X1 U91 ( .A1(data_out_b[1]), .A2(n23), .B1(adder[1]), .B2(n17), .C1(
        n63), .C2(f[1]), .ZN(n61) );
  INV_X1 U92 ( .A(n61), .ZN(n112) );
  AOI222_X1 U93 ( .A1(data_out_b[0]), .A2(n23), .B1(adder[0]), .B2(n17), .C1(
        n63), .C2(f[0]), .ZN(n62) );
  INV_X1 U94 ( .A(n62), .ZN(n113) );
  AOI222_X1 U95 ( .A1(data_out_b[9]), .A2(n23), .B1(adder[9]), .B2(n17), .C1(
        n63), .C2(f[9]), .ZN(n64) );
  INV_X1 U96 ( .A(n64), .ZN(n79) );
  NOR4_X1 U97 ( .A1(n50), .A2(n49), .A3(n48), .A4(n47), .ZN(n72) );
  NOR4_X1 U98 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n52), .ZN(n71) );
  NAND4_X1 U99 ( .A1(n68), .A2(n67), .A3(n66), .A4(n65), .ZN(n69) );
  NOR4_X1 U100 ( .A1(n69), .A2(f[0]), .A3(f[1]), .A4(f[2]), .ZN(n70) );
  NAND3_X1 U101 ( .A1(n72), .A2(n71), .A3(n70), .ZN(n74) );
  NAND3_X1 U102 ( .A1(wr_en_y), .A2(n74), .A3(n73), .ZN(n242) );
  OAI22_X1 U103 ( .A1(n182), .A2(n243), .B1(n214), .B2(n242), .ZN(n181) );
  OAI22_X1 U104 ( .A1(n183), .A2(n243), .B1(n215), .B2(n242), .ZN(n180) );
  OAI22_X1 U105 ( .A1(n184), .A2(n243), .B1(n216), .B2(n242), .ZN(n179) );
  OAI22_X1 U106 ( .A1(n192), .A2(n243), .B1(n220), .B2(n242), .ZN(n171) );
  OAI22_X1 U107 ( .A1(n193), .A2(n243), .B1(n221), .B2(n242), .ZN(n170) );
  OAI22_X1 U108 ( .A1(n194), .A2(n243), .B1(n222), .B2(n242), .ZN(n169) );
  OAI22_X1 U109 ( .A1(n195), .A2(n243), .B1(n223), .B2(n242), .ZN(n168) );
  OAI22_X1 U110 ( .A1(n196), .A2(n243), .B1(n224), .B2(n242), .ZN(n167) );
  OAI22_X1 U111 ( .A1(n197), .A2(n243), .B1(n73), .B2(n242), .ZN(n166) );
  AND4_X1 U112 ( .A1(sel[3]), .A2(sel[2]), .A3(sel[1]), .A4(sel[0]), .ZN(n75)
         );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_10_DW_mult_tc_1 ( a, b, 
        product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n9, n13, n16, n18, n19, n23, n25, n27, n29, n31, n34, n36,
         n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n50, n53, n54, n55,
         n56, n57, n58, n59, n62, n63, n64, n65, n67, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n93, n95, n96, n97, n98, n99, n103, n104, n105, n106,
         n107, n109, n111, n112, n113, n114, n115, n117, n119, n120, n122,
         n127, n135, n139, n141, n142, n143, n144, n145, n147, n148, n149,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n241, n247, n249,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n418, n419, n420, n421, n422, n423,
         n424, n426, n427, n429, n432, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U148 ( .A(n265), .B(n144), .Z(n145) );
  XOR2_X1 U152 ( .A(n301), .B(n148), .Z(n149) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U161 ( .A(n177), .B(n168), .CI(n166), .CO(n163), .S(n164) );
  FA_X1 U162 ( .A(n170), .B(n172), .CI(n179), .CO(n165), .S(n166) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n263), .CI(n291), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n317), .B(n252), .CO(n173), .S(n174) );
  FA_X1 U167 ( .A(n180), .B(n187), .CI(n178), .CO(n175), .S(n176) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U169 ( .A(n193), .B(n282), .CI(n191), .CO(n179), .S(n180) );
  FA_X1 U170 ( .A(n268), .B(n274), .CI(n292), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U172 ( .A(n197), .B(n190), .CI(n188), .CO(n185), .S(n186) );
  FA_X1 U173 ( .A(n199), .B(n201), .CI(n192), .CO(n187), .S(n188) );
  FA_X1 U174 ( .A(n275), .B(n293), .CI(n194), .CO(n189), .S(n190) );
  FA_X1 U175 ( .A(n283), .B(n253), .CI(n305), .CO(n191), .S(n192) );
  HA_X1 U176 ( .A(n269), .B(n319), .CO(n193), .S(n194) );
  FA_X1 U177 ( .A(n205), .B(n200), .CI(n198), .CO(n195), .S(n196) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U179 ( .A(n276), .B(n284), .CI(n294), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n320), .B(n270), .CI(n306), .CO(n201), .S(n202) );
  FA_X1 U182 ( .A(n210), .B(n307), .CI(n215), .CO(n205), .S(n206) );
  FA_X1 U183 ( .A(n254), .B(n285), .CI(n295), .CO(n207), .S(n208) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U185 ( .A(n216), .B(n219), .CI(n214), .CO(n211), .S(n212) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n322), .B(n278), .CI(n308), .CO(n215), .S(n216) );
  FA_X1 U188 ( .A(n225), .B(n222), .CI(n220), .CO(n217), .S(n218) );
  FA_X1 U189 ( .A(n255), .B(n309), .CI(n297), .CO(n219), .S(n220) );
  HA_X1 U190 ( .A(n287), .B(n323), .CO(n221), .S(n222) );
  FA_X1 U191 ( .A(n229), .B(n298), .CI(n226), .CO(n223), .S(n224) );
  FA_X1 U192 ( .A(n324), .B(n288), .CI(n310), .CO(n225), .S(n226) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  HA_X1 U194 ( .A(n311), .B(n325), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n326), .B(n300), .CI(n312), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  OR2_X1 U414 ( .A1(n228), .A2(n231), .ZN(n490) );
  OR2_X2 U415 ( .A1(n224), .A2(n227), .ZN(n566) );
  BUF_X1 U416 ( .A(n587), .Z(n491) );
  OR2_X1 U417 ( .A1(n548), .A2(n249), .ZN(n6) );
  XOR2_X2 U418 ( .A(n587), .B(a[10]), .Z(n508) );
  CLKBUF_X1 U419 ( .A(n583), .Z(n516) );
  OR2_X1 U420 ( .A1(n545), .A2(n560), .ZN(n504) );
  OR2_X1 U421 ( .A1(n329), .A2(n258), .ZN(n492) );
  CLKBUF_X1 U422 ( .A(n550), .Z(n493) );
  OR2_X1 U423 ( .A1(n196), .A2(n203), .ZN(n494) );
  XNOR2_X1 U424 ( .A(n271), .B(n495), .ZN(n147) );
  XNOR2_X1 U425 ( .A(n289), .B(n279), .ZN(n495) );
  XNOR2_X1 U426 ( .A(n45), .B(n496), .ZN(product[12]) );
  AND2_X1 U427 ( .A1(n541), .A2(n79), .ZN(n496) );
  NOR2_X1 U428 ( .A1(n186), .A2(n195), .ZN(n497) );
  NOR2_X1 U429 ( .A1(n186), .A2(n195), .ZN(n82) );
  BUF_X2 U430 ( .A(n16), .Z(n498) );
  OR2_X1 U431 ( .A1(n218), .A2(n223), .ZN(n499) );
  AOI21_X1 U432 ( .B1(n566), .B2(n104), .A(n543), .ZN(n500) );
  INV_X1 U433 ( .A(n249), .ZN(n501) );
  XOR2_X1 U434 ( .A(n590), .B(a[14]), .Z(n41) );
  INV_X1 U435 ( .A(n580), .ZN(n502) );
  OR2_X1 U436 ( .A1(n545), .A2(n560), .ZN(n503) );
  OR2_X1 U437 ( .A1(n545), .A2(n560), .ZN(n23) );
  BUF_X1 U438 ( .A(n588), .Z(n505) );
  XNOR2_X2 U439 ( .A(n584), .B(a[8]), .ZN(n506) );
  XOR2_X1 U440 ( .A(n588), .B(a[10]), .Z(n542) );
  OAI21_X1 U441 ( .B1(n105), .B2(n107), .A(n106), .ZN(n507) );
  BUF_X1 U442 ( .A(n526), .Z(n573) );
  XNOR2_X1 U443 ( .A(n579), .B(n577), .ZN(n548) );
  XOR2_X1 U444 ( .A(n505), .B(n424), .Z(n342) );
  AND2_X2 U445 ( .A1(n224), .A2(n227), .ZN(n543) );
  XOR2_X1 U446 ( .A(n208), .B(n213), .Z(n509) );
  XOR2_X1 U447 ( .A(n206), .B(n509), .Z(n204) );
  NAND2_X1 U448 ( .A1(n206), .A2(n208), .ZN(n510) );
  NAND2_X1 U449 ( .A1(n206), .A2(n213), .ZN(n511) );
  NAND2_X1 U450 ( .A1(n208), .A2(n213), .ZN(n512) );
  NAND3_X1 U451 ( .A1(n510), .A2(n511), .A3(n512), .ZN(n203) );
  XOR2_X1 U452 ( .A(n19), .B(a[6]), .Z(n513) );
  INV_X1 U453 ( .A(n513), .ZN(n545) );
  CLKBUF_X1 U454 ( .A(n523), .Z(n514) );
  INV_X1 U455 ( .A(n586), .ZN(n515) );
  BUF_X2 U456 ( .A(n9), .Z(n572) );
  NOR2_X1 U457 ( .A1(n164), .A2(n175), .ZN(n517) );
  XOR2_X1 U458 ( .A(n583), .B(a[6]), .Z(n518) );
  CLKBUF_X1 U459 ( .A(n559), .Z(n519) );
  NAND2_X1 U460 ( .A1(n176), .A2(n185), .ZN(n79) );
  NOR2_X1 U461 ( .A1(n164), .A2(n175), .ZN(n75) );
  CLKBUF_X1 U462 ( .A(n504), .Z(n520) );
  CLKBUF_X1 U463 ( .A(n503), .Z(n521) );
  INV_X1 U464 ( .A(n578), .ZN(n522) );
  INV_X2 U465 ( .A(n579), .ZN(n574) );
  XNOR2_X1 U466 ( .A(n516), .B(a[4]), .ZN(n561) );
  XNOR2_X1 U467 ( .A(n491), .B(a[8]), .ZN(n429) );
  INV_X1 U468 ( .A(n581), .ZN(n523) );
  INV_X1 U469 ( .A(n581), .ZN(n580) );
  INV_X1 U470 ( .A(n531), .ZN(n524) );
  NAND2_X1 U471 ( .A1(n429), .A2(n27), .ZN(n525) );
  XOR2_X1 U472 ( .A(n579), .B(a[2]), .Z(n526) );
  CLKBUF_X1 U473 ( .A(n518), .Z(n527) );
  BUF_X2 U474 ( .A(n518), .Z(n528) );
  CLKBUF_X1 U475 ( .A(n518), .Z(n529) );
  AOI21_X1 U476 ( .B1(n566), .B2(n507), .A(n543), .ZN(n530) );
  AOI21_X1 U477 ( .B1(n566), .B2(n104), .A(n543), .ZN(n99) );
  XOR2_X1 U478 ( .A(n7), .B(a[4]), .Z(n531) );
  INV_X1 U479 ( .A(n540), .ZN(n37) );
  NAND2_X1 U480 ( .A1(n561), .A2(n16), .ZN(n532) );
  NAND2_X1 U481 ( .A1(n561), .A2(n524), .ZN(n18) );
  INV_X1 U482 ( .A(n582), .ZN(n533) );
  OAI21_X1 U483 ( .B1(n500), .B2(n97), .A(n98), .ZN(n534) );
  OAI21_X1 U484 ( .B1(n530), .B2(n97), .A(n98), .ZN(n535) );
  INV_X1 U485 ( .A(n585), .ZN(n536) );
  INV_X1 U486 ( .A(n585), .ZN(n537) );
  INV_X1 U487 ( .A(n585), .ZN(n584) );
  OAI21_X1 U488 ( .B1(n99), .B2(n97), .A(n98), .ZN(n96) );
  NAND2_X1 U489 ( .A1(n429), .A2(n27), .ZN(n29) );
  OR2_X1 U490 ( .A1(n164), .A2(n175), .ZN(n538) );
  INV_X1 U491 ( .A(n588), .ZN(n539) );
  XNOR2_X1 U492 ( .A(n588), .B(a[12]), .ZN(n540) );
  OR2_X1 U493 ( .A1(n176), .A2(n185), .ZN(n541) );
  INV_X1 U494 ( .A(n543), .ZN(n103) );
  OR2_X2 U495 ( .A1(n542), .A2(n555), .ZN(n34) );
  XNOR2_X1 U496 ( .A(n581), .B(a[2]), .ZN(n432) );
  OR2_X1 U497 ( .A1(n204), .A2(n211), .ZN(n544) );
  XNOR2_X1 U498 ( .A(n584), .B(a[8]), .ZN(n27) );
  XNOR2_X1 U499 ( .A(n554), .B(n546), .ZN(product[9]) );
  AND2_X1 U500 ( .A1(n544), .A2(n90), .ZN(n546) );
  XNOR2_X1 U501 ( .A(n88), .B(n547), .ZN(product[10]) );
  NAND2_X1 U502 ( .A1(n494), .A2(n86), .ZN(n547) );
  OR2_X2 U503 ( .A1(n548), .A2(n249), .ZN(n549) );
  INV_X2 U504 ( .A(n583), .ZN(n582) );
  INV_X1 U505 ( .A(n249), .ZN(n577) );
  NAND2_X1 U506 ( .A1(n432), .A2(n9), .ZN(n550) );
  CLKBUF_X1 U507 ( .A(n107), .Z(n551) );
  NAND2_X1 U508 ( .A1(n432), .A2(n526), .ZN(n558) );
  AOI21_X1 U509 ( .B1(n534), .B2(n563), .A(n93), .ZN(n552) );
  AOI21_X1 U510 ( .B1(n96), .B2(n563), .A(n93), .ZN(n553) );
  CLKBUF_X1 U511 ( .A(n552), .Z(n554) );
  XNOR2_X1 U512 ( .A(n587), .B(a[10]), .ZN(n555) );
  OAI21_X1 U513 ( .B1(n552), .B2(n89), .A(n90), .ZN(n556) );
  BUF_X2 U514 ( .A(n16), .Z(n557) );
  INV_X2 U515 ( .A(n587), .ZN(n586) );
  AOI21_X1 U516 ( .B1(n556), .B2(n80), .A(n81), .ZN(n559) );
  XNOR2_X1 U517 ( .A(n583), .B(a[6]), .ZN(n560) );
  BUF_X1 U518 ( .A(n43), .Z(n575) );
  AOI21_X1 U519 ( .B1(n74), .B2(n562), .A(n67), .ZN(n65) );
  INV_X1 U520 ( .A(n69), .ZN(n67) );
  NAND2_X1 U521 ( .A1(n73), .A2(n562), .ZN(n64) );
  INV_X1 U522 ( .A(n73), .ZN(n71) );
  NAND2_X1 U523 ( .A1(n562), .A2(n69), .ZN(n47) );
  INV_X1 U524 ( .A(n74), .ZN(n72) );
  INV_X1 U525 ( .A(n95), .ZN(n93) );
  NAND2_X1 U526 ( .A1(n538), .A2(n76), .ZN(n48) );
  OR2_X1 U527 ( .A1(n152), .A2(n163), .ZN(n562) );
  XNOR2_X1 U528 ( .A(n84), .B(n50), .ZN(product[11]) );
  NAND2_X1 U529 ( .A1(n127), .A2(n83), .ZN(n50) );
  NAND2_X1 U530 ( .A1(n152), .A2(n163), .ZN(n69) );
  NAND2_X1 U531 ( .A1(n563), .A2(n95), .ZN(n53) );
  INV_X1 U532 ( .A(n111), .ZN(n109) );
  OAI21_X1 U533 ( .B1(n115), .B2(n113), .A(n114), .ZN(n112) );
  NAND2_X1 U534 ( .A1(n490), .A2(n106), .ZN(n56) );
  NAND2_X1 U535 ( .A1(n499), .A2(n98), .ZN(n54) );
  AOI21_X1 U536 ( .B1(n564), .B2(n120), .A(n117), .ZN(n115) );
  INV_X1 U537 ( .A(n119), .ZN(n117) );
  NAND2_X1 U538 ( .A1(n566), .A2(n103), .ZN(n55) );
  XOR2_X1 U539 ( .A(n58), .B(n115), .Z(product[3]) );
  NAND2_X1 U540 ( .A1(n135), .A2(n114), .ZN(n58) );
  INV_X1 U541 ( .A(n113), .ZN(n135) );
  NOR2_X1 U542 ( .A1(n176), .A2(n185), .ZN(n78) );
  NOR2_X1 U543 ( .A1(n196), .A2(n203), .ZN(n85) );
  XNOR2_X1 U544 ( .A(n57), .B(n112), .ZN(product[4]) );
  NAND2_X1 U545 ( .A1(n567), .A2(n111), .ZN(n57) );
  XNOR2_X1 U546 ( .A(n59), .B(n120), .ZN(product[2]) );
  NAND2_X1 U547 ( .A1(n564), .A2(n119), .ZN(n59) );
  NAND2_X1 U548 ( .A1(n212), .A2(n217), .ZN(n95) );
  NAND2_X1 U549 ( .A1(n164), .A2(n175), .ZN(n76) );
  OR2_X1 U550 ( .A1(n212), .A2(n217), .ZN(n563) );
  NAND2_X1 U551 ( .A1(n204), .A2(n211), .ZN(n90) );
  NAND2_X1 U552 ( .A1(n196), .A2(n203), .ZN(n86) );
  XNOR2_X1 U553 ( .A(n63), .B(n46), .ZN(product[15]) );
  NAND2_X1 U554 ( .A1(n565), .A2(n62), .ZN(n46) );
  OR2_X1 U555 ( .A1(n328), .A2(n314), .ZN(n564) );
  OR2_X1 U556 ( .A1(n151), .A2(n139), .ZN(n565) );
  NOR2_X1 U557 ( .A1(n228), .A2(n231), .ZN(n105) );
  NOR2_X1 U558 ( .A1(n218), .A2(n223), .ZN(n97) );
  NAND2_X1 U559 ( .A1(n218), .A2(n223), .ZN(n98) );
  NAND2_X1 U560 ( .A1(n228), .A2(n231), .ZN(n106) );
  OR2_X1 U561 ( .A1(n233), .A2(n232), .ZN(n567) );
  INV_X1 U562 ( .A(n41), .ZN(n235) );
  AND2_X1 U563 ( .A1(n492), .A2(n122), .ZN(product[1]) );
  AND2_X1 U564 ( .A1(n576), .A2(n241), .ZN(n278) );
  OR2_X1 U565 ( .A1(n575), .A2(n502), .ZN(n392) );
  XNOR2_X1 U566 ( .A(n582), .B(n575), .ZN(n376) );
  XNOR2_X1 U567 ( .A(n586), .B(n575), .ZN(n352) );
  XNOR2_X1 U568 ( .A(n155), .B(n569), .ZN(n139) );
  XNOR2_X1 U569 ( .A(n153), .B(n141), .ZN(n569) );
  XNOR2_X1 U570 ( .A(n157), .B(n570), .ZN(n141) );
  XNOR2_X1 U571 ( .A(n145), .B(n143), .ZN(n570) );
  OAI22_X1 U572 ( .A1(n39), .A2(n590), .B1(n337), .B2(n37), .ZN(n252) );
  OR2_X1 U573 ( .A1(n575), .A2(n590), .ZN(n337) );
  XOR2_X1 U574 ( .A(n579), .B(a[2]), .Z(n9) );
  OAI22_X1 U575 ( .A1(n42), .A2(n592), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U576 ( .A1(n575), .A2(n592), .ZN(n332) );
  XNOR2_X1 U577 ( .A(n539), .B(n575), .ZN(n343) );
  AND2_X1 U578 ( .A1(n576), .A2(n531), .ZN(n300) );
  XNOR2_X1 U579 ( .A(n159), .B(n571), .ZN(n142) );
  XNOR2_X1 U580 ( .A(n315), .B(n261), .ZN(n571) );
  XNOR2_X1 U581 ( .A(n589), .B(n575), .ZN(n336) );
  NAND2_X1 U582 ( .A1(n427), .A2(n37), .ZN(n39) );
  XOR2_X1 U583 ( .A(n589), .B(a[12]), .Z(n427) );
  OAI22_X1 U584 ( .A1(n39), .A2(n336), .B1(n37), .B2(n335), .ZN(n263) );
  AND2_X1 U585 ( .A1(n576), .A2(n235), .ZN(n260) );
  OAI22_X1 U586 ( .A1(n39), .A2(n335), .B1(n37), .B2(n334), .ZN(n262) );
  AND2_X1 U587 ( .A1(n576), .A2(n560), .ZN(n288) );
  AND2_X1 U588 ( .A1(n576), .A2(n555), .ZN(n270) );
  INV_X1 U589 ( .A(n19), .ZN(n585) );
  INV_X1 U590 ( .A(n25), .ZN(n587) );
  NAND2_X1 U591 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U592 ( .A(n591), .B(a[14]), .Z(n426) );
  INV_X1 U593 ( .A(n7), .ZN(n581) );
  XNOR2_X1 U594 ( .A(n537), .B(n575), .ZN(n363) );
  AND2_X1 U595 ( .A1(n576), .A2(n247), .ZN(n314) );
  AND2_X1 U596 ( .A1(n576), .A2(n540), .ZN(n264) );
  AND2_X1 U597 ( .A1(n576), .A2(n249), .ZN(product[0]) );
  OR2_X1 U598 ( .A1(n575), .A2(n585), .ZN(n364) );
  OR2_X1 U599 ( .A1(n575), .A2(n515), .ZN(n353) );
  OR2_X1 U600 ( .A1(n505), .A2(n575), .ZN(n344) );
  OR2_X1 U601 ( .A1(n575), .A2(n533), .ZN(n377) );
  XNOR2_X1 U602 ( .A(n536), .B(b[9]), .ZN(n354) );
  OAI22_X1 U603 ( .A1(n39), .A2(n334), .B1(n37), .B2(n333), .ZN(n261) );
  XNOR2_X1 U604 ( .A(n589), .B(n422), .ZN(n333) );
  XNOR2_X1 U605 ( .A(n582), .B(b[11]), .ZN(n365) );
  XNOR2_X1 U606 ( .A(n589), .B(n423), .ZN(n334) );
  XNOR2_X1 U607 ( .A(n589), .B(n424), .ZN(n335) );
  OAI22_X1 U608 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U609 ( .A(n591), .B(n424), .ZN(n330) );
  XNOR2_X1 U610 ( .A(n591), .B(n575), .ZN(n331) );
  XNOR2_X1 U611 ( .A(n586), .B(n418), .ZN(n345) );
  XNOR2_X1 U612 ( .A(n539), .B(n420), .ZN(n338) );
  XNOR2_X1 U613 ( .A(n514), .B(b[13]), .ZN(n378) );
  XNOR2_X1 U614 ( .A(n537), .B(n424), .ZN(n362) );
  XNOR2_X1 U615 ( .A(n586), .B(n424), .ZN(n351) );
  XNOR2_X1 U616 ( .A(n539), .B(n423), .ZN(n341) );
  XNOR2_X1 U617 ( .A(n539), .B(n422), .ZN(n340) );
  XNOR2_X1 U618 ( .A(n580), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U619 ( .A(n580), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U620 ( .A(n580), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U621 ( .A(n523), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U622 ( .A(n514), .B(n419), .ZN(n385) );
  XNOR2_X1 U623 ( .A(n523), .B(n418), .ZN(n384) );
  XNOR2_X1 U624 ( .A(n580), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U625 ( .A(n537), .B(n423), .ZN(n361) );
  XNOR2_X1 U626 ( .A(n586), .B(n423), .ZN(n350) );
  XNOR2_X1 U627 ( .A(n536), .B(n422), .ZN(n360) );
  XNOR2_X1 U628 ( .A(n586), .B(n422), .ZN(n349) );
  XNOR2_X1 U629 ( .A(n582), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U630 ( .A(n582), .B(n418), .ZN(n369) );
  XNOR2_X1 U631 ( .A(n582), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U632 ( .A(n582), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U633 ( .A(n537), .B(n420), .ZN(n358) );
  XNOR2_X1 U634 ( .A(n586), .B(n420), .ZN(n347) );
  XNOR2_X1 U635 ( .A(n536), .B(n418), .ZN(n356) );
  XNOR2_X1 U636 ( .A(n574), .B(b[13]), .ZN(n395) );
  XNOR2_X1 U637 ( .A(n586), .B(n419), .ZN(n346) );
  XNOR2_X1 U638 ( .A(n536), .B(n419), .ZN(n357) );
  XNOR2_X1 U639 ( .A(n574), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U640 ( .A(n537), .B(b[8]), .ZN(n355) );
  BUF_X1 U641 ( .A(n43), .Z(n576) );
  XNOR2_X1 U642 ( .A(n574), .B(b[15]), .ZN(n393) );
  XNOR2_X1 U643 ( .A(n539), .B(n421), .ZN(n339) );
  XNOR2_X1 U644 ( .A(n586), .B(n421), .ZN(n348) );
  XNOR2_X1 U645 ( .A(n536), .B(n421), .ZN(n359) );
  XNOR2_X1 U646 ( .A(n7), .B(a[4]), .ZN(n16) );
  NOR2_X1 U647 ( .A1(n75), .A2(n78), .ZN(n73) );
  OAI21_X1 U648 ( .B1(n517), .B2(n79), .A(n76), .ZN(n74) );
  OAI22_X1 U649 ( .A1(n34), .A2(n339), .B1(n338), .B2(n508), .ZN(n265) );
  OAI22_X1 U650 ( .A1(n34), .A2(n340), .B1(n339), .B2(n508), .ZN(n266) );
  OAI22_X1 U651 ( .A1(n34), .A2(n342), .B1(n341), .B2(n508), .ZN(n268) );
  OAI22_X1 U652 ( .A1(n34), .A2(n341), .B1(n340), .B2(n508), .ZN(n267) );
  OAI22_X1 U653 ( .A1(n34), .A2(n343), .B1(n342), .B2(n508), .ZN(n269) );
  OAI22_X1 U654 ( .A1(n34), .A2(n505), .B1(n344), .B2(n508), .ZN(n253) );
  INV_X1 U655 ( .A(n13), .ZN(n583) );
  XNOR2_X1 U656 ( .A(n55), .B(n507), .ZN(product[6]) );
  NAND2_X1 U657 ( .A1(n328), .A2(n314), .ZN(n119) );
  XNOR2_X1 U658 ( .A(n574), .B(b[14]), .ZN(n394) );
  XNOR2_X1 U659 ( .A(n578), .B(b[11]), .ZN(n397) );
  INV_X1 U660 ( .A(n1), .ZN(n579) );
  NOR2_X1 U661 ( .A1(n204), .A2(n211), .ZN(n89) );
  OAI22_X1 U662 ( .A1(n525), .A2(n346), .B1(n345), .B2(n506), .ZN(n271) );
  OAI22_X1 U663 ( .A1(n525), .A2(n350), .B1(n349), .B2(n506), .ZN(n275) );
  OAI22_X1 U664 ( .A1(n29), .A2(n351), .B1(n350), .B2(n506), .ZN(n276) );
  OAI22_X1 U665 ( .A1(n525), .A2(n347), .B1(n346), .B2(n506), .ZN(n272) );
  OAI22_X1 U666 ( .A1(n29), .A2(n515), .B1(n353), .B2(n506), .ZN(n254) );
  OAI22_X1 U667 ( .A1(n525), .A2(n348), .B1(n347), .B2(n506), .ZN(n273) );
  OAI22_X1 U668 ( .A1(n525), .A2(n349), .B1(n348), .B2(n506), .ZN(n274) );
  INV_X1 U669 ( .A(n27), .ZN(n241) );
  OAI22_X1 U670 ( .A1(n29), .A2(n352), .B1(n351), .B2(n506), .ZN(n277) );
  OR2_X1 U671 ( .A1(n575), .A2(n522), .ZN(n409) );
  INV_X1 U672 ( .A(n579), .ZN(n578) );
  XNOR2_X1 U673 ( .A(n582), .B(n419), .ZN(n370) );
  XNOR2_X1 U674 ( .A(n582), .B(n424), .ZN(n375) );
  XNOR2_X1 U675 ( .A(n582), .B(n420), .ZN(n371) );
  XNOR2_X1 U676 ( .A(n582), .B(n423), .ZN(n374) );
  XNOR2_X1 U677 ( .A(n582), .B(n422), .ZN(n373) );
  XNOR2_X1 U678 ( .A(n582), .B(n421), .ZN(n372) );
  OAI21_X1 U679 ( .B1(n87), .B2(n85), .A(n86), .ZN(n84) );
  XNOR2_X1 U680 ( .A(n77), .B(n48), .ZN(product[13]) );
  INV_X1 U681 ( .A(n497), .ZN(n127) );
  NOR2_X1 U682 ( .A1(n497), .A2(n85), .ZN(n80) );
  OAI21_X1 U683 ( .B1(n86), .B2(n82), .A(n83), .ZN(n81) );
  NAND2_X1 U684 ( .A1(n186), .A2(n195), .ZN(n83) );
  OAI21_X1 U685 ( .B1(n105), .B2(n107), .A(n106), .ZN(n104) );
  AOI21_X1 U686 ( .B1(n567), .B2(n112), .A(n109), .ZN(n107) );
  AOI21_X1 U687 ( .B1(n80), .B2(n556), .A(n81), .ZN(n45) );
  INV_X1 U688 ( .A(n88), .ZN(n87) );
  OAI21_X1 U689 ( .B1(n553), .B2(n89), .A(n90), .ZN(n88) );
  NOR2_X1 U690 ( .A1(n234), .A2(n257), .ZN(n113) );
  XNOR2_X1 U691 ( .A(n70), .B(n47), .ZN(product[14]) );
  OAI22_X1 U692 ( .A1(n520), .A2(n358), .B1(n357), .B2(n529), .ZN(n282) );
  OAI22_X1 U693 ( .A1(n504), .A2(n355), .B1(n354), .B2(n528), .ZN(n279) );
  OAI22_X1 U694 ( .A1(n503), .A2(n362), .B1(n361), .B2(n528), .ZN(n286) );
  OAI22_X1 U695 ( .A1(n521), .A2(n356), .B1(n355), .B2(n528), .ZN(n280) );
  OAI22_X1 U696 ( .A1(n503), .A2(n585), .B1(n364), .B2(n528), .ZN(n255) );
  OAI22_X1 U697 ( .A1(n503), .A2(n360), .B1(n359), .B2(n529), .ZN(n284) );
  OAI22_X1 U698 ( .A1(n504), .A2(n361), .B1(n360), .B2(n529), .ZN(n285) );
  OAI22_X1 U699 ( .A1(n503), .A2(n357), .B1(n356), .B2(n528), .ZN(n281) );
  OAI22_X1 U700 ( .A1(n504), .A2(n363), .B1(n362), .B2(n528), .ZN(n287) );
  OAI22_X1 U701 ( .A1(n23), .A2(n359), .B1(n358), .B2(n527), .ZN(n283) );
  OAI21_X1 U702 ( .B1(n64), .B2(n519), .A(n65), .ZN(n63) );
  XOR2_X1 U703 ( .A(n56), .B(n551), .Z(product[5]) );
  NAND2_X1 U704 ( .A1(n232), .A2(n233), .ZN(n111) );
  NAND2_X1 U705 ( .A1(n151), .A2(n139), .ZN(n62) );
  OAI22_X1 U706 ( .A1(n18), .A2(n370), .B1(n369), .B2(n557), .ZN(n293) );
  OAI22_X1 U707 ( .A1(n18), .A2(n367), .B1(n366), .B2(n557), .ZN(n290) );
  OAI22_X1 U708 ( .A1(n18), .A2(n375), .B1(n374), .B2(n557), .ZN(n298) );
  OAI22_X1 U709 ( .A1(n532), .A2(n373), .B1(n372), .B2(n498), .ZN(n296) );
  OAI22_X1 U710 ( .A1(n532), .A2(n372), .B1(n371), .B2(n498), .ZN(n295) );
  OAI22_X1 U711 ( .A1(n18), .A2(n368), .B1(n367), .B2(n498), .ZN(n291) );
  OAI22_X1 U712 ( .A1(n18), .A2(n369), .B1(n368), .B2(n498), .ZN(n292) );
  OAI22_X1 U713 ( .A1(n532), .A2(n374), .B1(n373), .B2(n557), .ZN(n297) );
  OAI22_X1 U714 ( .A1(n532), .A2(n376), .B1(n375), .B2(n498), .ZN(n299) );
  OAI22_X1 U715 ( .A1(n532), .A2(n533), .B1(n377), .B2(n498), .ZN(n256) );
  OAI22_X1 U716 ( .A1(n532), .A2(n371), .B1(n370), .B2(n557), .ZN(n294) );
  OAI22_X1 U717 ( .A1(n18), .A2(n366), .B1(n365), .B2(n557), .ZN(n289) );
  XNOR2_X1 U718 ( .A(n523), .B(n420), .ZN(n386) );
  XNOR2_X1 U719 ( .A(n523), .B(n421), .ZN(n387) );
  XNOR2_X1 U720 ( .A(n523), .B(n422), .ZN(n388) );
  XNOR2_X1 U721 ( .A(n580), .B(n575), .ZN(n391) );
  XNOR2_X1 U722 ( .A(n523), .B(n424), .ZN(n390) );
  XNOR2_X1 U723 ( .A(n580), .B(n423), .ZN(n389) );
  XNOR2_X1 U724 ( .A(n574), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U725 ( .A(n578), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U726 ( .A(n578), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U727 ( .A(n574), .B(n418), .ZN(n401) );
  XNOR2_X1 U728 ( .A(n578), .B(n419), .ZN(n402) );
  XNOR2_X1 U729 ( .A(n578), .B(n420), .ZN(n403) );
  XNOR2_X1 U730 ( .A(n574), .B(n575), .ZN(n408) );
  XNOR2_X1 U731 ( .A(n574), .B(n422), .ZN(n405) );
  XNOR2_X1 U732 ( .A(n574), .B(n421), .ZN(n404) );
  XNOR2_X1 U733 ( .A(n574), .B(n424), .ZN(n407) );
  XNOR2_X1 U734 ( .A(n574), .B(n423), .ZN(n406) );
  OAI21_X1 U735 ( .B1(n71), .B2(n559), .A(n72), .ZN(n70) );
  OAI21_X1 U736 ( .B1(n559), .B2(n78), .A(n79), .ZN(n77) );
  XNOR2_X1 U737 ( .A(n535), .B(n53), .ZN(product[8]) );
  OAI22_X1 U738 ( .A1(n549), .A2(n395), .B1(n394), .B2(n501), .ZN(n316) );
  OAI22_X1 U739 ( .A1(n549), .A2(n394), .B1(n393), .B2(n501), .ZN(n315) );
  OAI22_X1 U740 ( .A1(n549), .A2(n396), .B1(n395), .B2(n501), .ZN(n317) );
  OAI22_X1 U741 ( .A1(n549), .A2(n397), .B1(n396), .B2(n501), .ZN(n318) );
  OAI22_X1 U742 ( .A1(n549), .A2(n398), .B1(n397), .B2(n501), .ZN(n319) );
  OAI22_X1 U743 ( .A1(n549), .A2(n400), .B1(n399), .B2(n501), .ZN(n321) );
  OAI22_X1 U744 ( .A1(n549), .A2(n401), .B1(n400), .B2(n501), .ZN(n322) );
  OAI22_X1 U745 ( .A1(n6), .A2(n399), .B1(n398), .B2(n501), .ZN(n320) );
  OAI22_X1 U746 ( .A1(n6), .A2(n402), .B1(n401), .B2(n501), .ZN(n323) );
  OAI22_X1 U747 ( .A1(n6), .A2(n404), .B1(n403), .B2(n501), .ZN(n325) );
  OAI22_X1 U748 ( .A1(n403), .A2(n6), .B1(n402), .B2(n501), .ZN(n324) );
  OAI22_X1 U749 ( .A1(n549), .A2(n406), .B1(n405), .B2(n501), .ZN(n327) );
  OAI22_X1 U750 ( .A1(n549), .A2(n405), .B1(n404), .B2(n501), .ZN(n326) );
  OAI22_X1 U751 ( .A1(n549), .A2(n407), .B1(n406), .B2(n501), .ZN(n328) );
  OAI22_X1 U752 ( .A1(n549), .A2(n408), .B1(n407), .B2(n501), .ZN(n329) );
  INV_X1 U753 ( .A(n122), .ZN(n120) );
  NAND2_X1 U754 ( .A1(n258), .A2(n329), .ZN(n122) );
  OAI22_X1 U755 ( .A1(n549), .A2(n522), .B1(n409), .B2(n501), .ZN(n258) );
  XOR2_X1 U756 ( .A(n530), .B(n54), .Z(product[7]) );
  OAI22_X1 U757 ( .A1(n550), .A2(n379), .B1(n378), .B2(n572), .ZN(n301) );
  OAI22_X1 U758 ( .A1(n550), .A2(n380), .B1(n379), .B2(n572), .ZN(n302) );
  OAI22_X1 U759 ( .A1(n493), .A2(n385), .B1(n384), .B2(n572), .ZN(n307) );
  OAI22_X1 U760 ( .A1(n550), .A2(n382), .B1(n381), .B2(n572), .ZN(n304) );
  OAI22_X1 U761 ( .A1(n558), .A2(n381), .B1(n380), .B2(n572), .ZN(n303) );
  NAND2_X1 U762 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U763 ( .A1(n558), .A2(n383), .B1(n382), .B2(n573), .ZN(n305) );
  OAI22_X1 U764 ( .A1(n558), .A2(n384), .B1(n383), .B2(n573), .ZN(n306) );
  OAI22_X1 U765 ( .A1(n550), .A2(n386), .B1(n385), .B2(n572), .ZN(n308) );
  OAI22_X1 U766 ( .A1(n550), .A2(n387), .B1(n386), .B2(n572), .ZN(n309) );
  OAI22_X1 U767 ( .A1(n493), .A2(n502), .B1(n392), .B2(n572), .ZN(n257) );
  OAI22_X1 U768 ( .A1(n558), .A2(n389), .B1(n388), .B2(n573), .ZN(n311) );
  OAI22_X1 U769 ( .A1(n558), .A2(n388), .B1(n387), .B2(n573), .ZN(n310) );
  OAI22_X1 U770 ( .A1(n558), .A2(n390), .B1(n389), .B2(n572), .ZN(n312) );
  INV_X1 U771 ( .A(n572), .ZN(n247) );
  OAI22_X1 U772 ( .A1(n550), .A2(n391), .B1(n390), .B2(n572), .ZN(n313) );
  INV_X1 U773 ( .A(n31), .ZN(n588) );
  INV_X1 U774 ( .A(n590), .ZN(n589) );
  INV_X1 U775 ( .A(n36), .ZN(n590) );
  INV_X1 U776 ( .A(n592), .ZN(n591) );
  INV_X1 U777 ( .A(n40), .ZN(n592) );
  XOR2_X1 U778 ( .A(n259), .B(n251), .Z(n148) );
  XOR2_X1 U779 ( .A(n149), .B(n147), .Z(n144) );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_10_DW01_add_2 ( A, B, CI, 
        SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n9, n10, n11, n12, n13, n14, n15, n16, n19, n20, n22,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n44, n45, n47, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n65, n67, n68, n69, n70, n71, n73,
         n75, n76, n77, n78, n79, n81, n83, n84, n86, n88, n89, n90, n91, n95,
         n96, n98, n100, n157, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182;

  OR2_X2 U122 ( .A1(A[10]), .A2(B[10]), .ZN(n178) );
  NOR2_X2 U123 ( .A1(A[11]), .A2(B[11]), .ZN(n35) );
  INV_X1 U124 ( .A(n173), .ZN(n44) );
  OR2_X1 U125 ( .A1(A[8]), .A2(B[8]), .ZN(n157) );
  AND2_X1 U126 ( .A1(n176), .A2(n86), .ZN(SUM[0]) );
  OR2_X1 U127 ( .A1(A[15]), .A2(B[15]), .ZN(n159) );
  XNOR2_X1 U128 ( .A(n51), .B(n160), .ZN(SUM[9]) );
  AND2_X1 U129 ( .A1(n179), .A2(n49), .ZN(n160) );
  NOR2_X1 U130 ( .A1(A[8]), .A2(B[8]), .ZN(n161) );
  NOR2_X1 U131 ( .A1(A[8]), .A2(B[8]), .ZN(n54) );
  XNOR2_X1 U132 ( .A(n45), .B(n162), .ZN(SUM[10]) );
  AND2_X1 U133 ( .A1(n178), .A2(n44), .ZN(n162) );
  INV_X1 U134 ( .A(n91), .ZN(n163) );
  XNOR2_X1 U135 ( .A(n164), .B(n37), .ZN(SUM[11]) );
  AND2_X1 U136 ( .A1(n91), .A2(n36), .ZN(n164) );
  AOI21_X2 U137 ( .B1(n52), .B2(n60), .A(n53), .ZN(n51) );
  NOR2_X1 U138 ( .A1(A[14]), .A2(B[14]), .ZN(n165) );
  NOR2_X1 U139 ( .A1(A[14]), .A2(B[14]), .ZN(n25) );
  AOI21_X1 U140 ( .B1(n178), .B2(n47), .A(n173), .ZN(n166) );
  CLKBUF_X1 U141 ( .A(n29), .Z(n167) );
  OAI21_X1 U142 ( .B1(n39), .B2(n51), .A(n166), .ZN(n168) );
  OAI21_X1 U143 ( .B1(n32), .B2(n36), .A(n33), .ZN(n169) );
  NOR2_X1 U144 ( .A1(n172), .A2(n35), .ZN(n170) );
  CLKBUF_X1 U145 ( .A(n36), .Z(n171) );
  NOR2_X1 U146 ( .A1(A[12]), .A2(B[12]), .ZN(n172) );
  NOR2_X1 U147 ( .A1(A[12]), .A2(B[12]), .ZN(n32) );
  AND2_X1 U148 ( .A1(A[10]), .A2(B[10]), .ZN(n173) );
  AOI21_X1 U149 ( .B1(n168), .B2(n170), .A(n169), .ZN(n174) );
  AOI21_X1 U150 ( .B1(n38), .B2(n30), .A(n31), .ZN(n175) );
  INV_X1 U151 ( .A(n24), .ZN(n22) );
  OR2_X1 U152 ( .A1(A[0]), .A2(B[0]), .ZN(n176) );
  INV_X1 U153 ( .A(n60), .ZN(n59) );
  INV_X1 U154 ( .A(n51), .ZN(n50) );
  AOI21_X1 U155 ( .B1(n178), .B2(n47), .A(n173), .ZN(n40) );
  AOI21_X1 U156 ( .B1(n180), .B2(n76), .A(n73), .ZN(n71) );
  INV_X1 U157 ( .A(n75), .ZN(n73) );
  AOI21_X1 U158 ( .B1(n181), .B2(n84), .A(n81), .ZN(n79) );
  INV_X1 U159 ( .A(n83), .ZN(n81) );
  OAI21_X1 U160 ( .B1(n79), .B2(n77), .A(n78), .ZN(n76) );
  AOI21_X1 U161 ( .B1(n182), .B2(n68), .A(n65), .ZN(n63) );
  INV_X1 U162 ( .A(n67), .ZN(n65) );
  OR2_X1 U163 ( .A1(n165), .A2(n28), .ZN(n177) );
  OAI21_X1 U164 ( .B1(n71), .B2(n69), .A(n70), .ZN(n68) );
  AOI21_X1 U165 ( .B1(n50), .B2(n179), .A(n47), .ZN(n45) );
  NAND2_X1 U166 ( .A1(n157), .A2(n55), .ZN(n9) );
  INV_X1 U167 ( .A(n86), .ZN(n84) );
  OAI21_X1 U168 ( .B1(n59), .B2(n57), .A(n58), .ZN(n56) );
  INV_X1 U169 ( .A(n49), .ZN(n47) );
  NAND2_X1 U170 ( .A1(n98), .A2(n70), .ZN(n13) );
  INV_X1 U171 ( .A(n69), .ZN(n98) );
  NAND2_X1 U172 ( .A1(n95), .A2(n58), .ZN(n10) );
  INV_X1 U173 ( .A(n57), .ZN(n95) );
  NAND2_X1 U174 ( .A1(n100), .A2(n78), .ZN(n15) );
  INV_X1 U175 ( .A(n77), .ZN(n100) );
  NAND2_X1 U176 ( .A1(n182), .A2(n67), .ZN(n12) );
  NAND2_X1 U177 ( .A1(n180), .A2(n75), .ZN(n14) );
  NAND2_X1 U178 ( .A1(n181), .A2(n83), .ZN(n16) );
  NAND2_X1 U179 ( .A1(n96), .A2(n62), .ZN(n11) );
  INV_X1 U180 ( .A(n61), .ZN(n96) );
  NAND2_X1 U181 ( .A1(n88), .A2(n26), .ZN(n3) );
  XNOR2_X1 U182 ( .A(n34), .B(n5), .ZN(SUM[12]) );
  NAND2_X1 U183 ( .A1(n90), .A2(n33), .ZN(n5) );
  XOR2_X1 U184 ( .A(n59), .B(n10), .Z(SUM[7]) );
  XOR2_X1 U185 ( .A(n13), .B(n71), .Z(SUM[4]) );
  NOR2_X1 U186 ( .A1(A[7]), .A2(B[7]), .ZN(n57) );
  NAND2_X1 U187 ( .A1(n89), .A2(n29), .ZN(n4) );
  OR2_X1 U188 ( .A1(A[9]), .A2(B[9]), .ZN(n179) );
  NOR2_X1 U189 ( .A1(A[4]), .A2(B[4]), .ZN(n69) );
  NOR2_X1 U190 ( .A1(A[2]), .A2(B[2]), .ZN(n77) );
  NAND2_X1 U191 ( .A1(A[11]), .A2(B[11]), .ZN(n36) );
  OR2_X1 U192 ( .A1(A[3]), .A2(B[3]), .ZN(n180) );
  OR2_X1 U193 ( .A1(A[1]), .A2(B[1]), .ZN(n181) );
  XNOR2_X1 U194 ( .A(n56), .B(n9), .ZN(SUM[8]) );
  XNOR2_X1 U195 ( .A(n14), .B(n76), .ZN(SUM[3]) );
  XNOR2_X1 U196 ( .A(n16), .B(n84), .ZN(SUM[1]) );
  NOR2_X1 U197 ( .A1(A[6]), .A2(B[6]), .ZN(n61) );
  NAND2_X1 U198 ( .A1(A[7]), .A2(B[7]), .ZN(n58) );
  OR2_X1 U199 ( .A1(A[5]), .A2(B[5]), .ZN(n182) );
  NAND2_X1 U200 ( .A1(A[4]), .A2(B[4]), .ZN(n70) );
  NAND2_X1 U201 ( .A1(A[2]), .A2(B[2]), .ZN(n78) );
  NAND2_X1 U202 ( .A1(A[9]), .A2(B[9]), .ZN(n49) );
  NAND2_X1 U203 ( .A1(A[5]), .A2(B[5]), .ZN(n67) );
  NAND2_X1 U204 ( .A1(A[3]), .A2(B[3]), .ZN(n75) );
  NAND2_X1 U205 ( .A1(A[1]), .A2(B[1]), .ZN(n83) );
  NAND2_X1 U206 ( .A1(A[0]), .A2(B[0]), .ZN(n86) );
  NAND2_X1 U207 ( .A1(A[8]), .A2(B[8]), .ZN(n55) );
  NAND2_X1 U208 ( .A1(A[6]), .A2(B[6]), .ZN(n62) );
  NAND2_X1 U209 ( .A1(A[13]), .A2(B[13]), .ZN(n29) );
  XNOR2_X1 U210 ( .A(n12), .B(n68), .ZN(SUM[5]) );
  XOR2_X1 U211 ( .A(n15), .B(n79), .Z(SUM[2]) );
  NAND2_X1 U212 ( .A1(n159), .A2(n19), .ZN(n2) );
  OAI21_X1 U213 ( .B1(n25), .B2(n29), .A(n26), .ZN(n24) );
  INV_X1 U214 ( .A(n172), .ZN(n90) );
  NAND2_X1 U215 ( .A1(A[12]), .A2(B[12]), .ZN(n33) );
  NOR2_X1 U216 ( .A1(n161), .A2(n57), .ZN(n52) );
  OAI21_X1 U217 ( .B1(n54), .B2(n58), .A(n55), .ZN(n53) );
  XOR2_X1 U218 ( .A(n11), .B(n63), .Z(SUM[6]) );
  OAI21_X1 U219 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  NAND2_X1 U220 ( .A1(A[14]), .A2(B[14]), .ZN(n26) );
  INV_X1 U221 ( .A(n165), .ZN(n88) );
  INV_X1 U222 ( .A(n28), .ZN(n89) );
  NOR2_X1 U223 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  OAI21_X1 U224 ( .B1(n32), .B2(n36), .A(n33), .ZN(n31) );
  INV_X1 U225 ( .A(n168), .ZN(n37) );
  OAI21_X1 U226 ( .B1(n37), .B2(n163), .A(n171), .ZN(n34) );
  INV_X1 U227 ( .A(n35), .ZN(n91) );
  NOR2_X1 U228 ( .A1(n172), .A2(n35), .ZN(n30) );
  NAND2_X1 U229 ( .A1(A[15]), .A2(B[15]), .ZN(n19) );
  OAI21_X1 U230 ( .B1(n39), .B2(n51), .A(n40), .ZN(n38) );
  XNOR2_X1 U231 ( .A(n20), .B(n2), .ZN(SUM[15]) );
  NAND2_X1 U232 ( .A1(n178), .A2(n179), .ZN(n39) );
  XNOR2_X1 U233 ( .A(n27), .B(n3), .ZN(SUM[14]) );
  XOR2_X1 U234 ( .A(n175), .B(n4), .Z(SUM[13]) );
  OAI21_X1 U235 ( .B1(n175), .B2(n28), .A(n167), .ZN(n27) );
  OAI21_X1 U236 ( .B1(n174), .B2(n177), .A(n22), .ZN(n20) );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_10 ( clk, clear_acc, 
        data_out_x, data_out, data_out_w, data_out_b, wr_en_y, m_valid, 
        m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [4:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
         N39, N40, N41, N42, N43, N44, n1, n2, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n85, n102, n111, n112, n113, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n17), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n218), .CK(clk), .Q(n20) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n219), .CK(clk), .Q(n21) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n220), .CK(clk), .Q(n22) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n221), .CK(clk), .Q(n23) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n222), .CK(clk), .Q(n24) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n223), .CK(clk), .Q(n25) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n224), .CK(clk), .Q(n26) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n225), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n226), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n227), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n228), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n229), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n230), .CK(clk), .Q(n34) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n231), .CK(clk), .Q(n35) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n232), .CK(clk), .Q(n36) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n233), .CK(clk), .Q(n37) );
  DFF_X1 \f_reg[0]  ( .D(n83), .CK(clk), .Q(f[0]), .QN(n206) );
  DFF_X1 \f_reg[1]  ( .D(n82), .CK(clk), .Q(f[1]), .QN(n207) );
  DFF_X1 \f_reg[2]  ( .D(n81), .CK(clk), .Q(f[2]), .QN(n208) );
  DFF_X1 \f_reg[3]  ( .D(n80), .CK(clk), .Q(f[3]), .QN(n209) );
  DFF_X1 \f_reg[7]  ( .D(n76), .CK(clk), .Q(f[7]), .QN(n210) );
  DFF_X1 \f_reg[8]  ( .D(n75), .CK(clk), .Q(f[8]), .QN(n211) );
  DFF_X1 \f_reg[9]  ( .D(n74), .CK(clk), .Q(f[9]), .QN(n212) );
  DFF_X1 \f_reg[10]  ( .D(n73), .CK(clk), .Q(n47), .QN(n213) );
  DFF_X1 \f_reg[11]  ( .D(n72), .CK(clk), .Q(n45), .QN(n214) );
  DFF_X1 \f_reg[12]  ( .D(n2), .CK(clk), .Q(n44), .QN(n215) );
  DFF_X1 \f_reg[13]  ( .D(n71), .CK(clk), .Q(n42), .QN(n216) );
  DFF_X1 \f_reg[14]  ( .D(n4), .CK(clk), .Q(n41), .QN(n217) );
  DFF_X1 \f_reg[15]  ( .D(n70), .CK(clk), .Q(f[15]), .QN(n67) );
  DFF_X1 \data_out_reg[15]  ( .D(n102), .CK(clk), .Q(data_out[15]), .QN(n189)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n111), .CK(clk), .Q(data_out[14]), .QN(n188)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n112), .CK(clk), .Q(data_out[13]), .QN(n187)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n113), .CK(clk), .Q(data_out[12]), .QN(n186)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n162), .CK(clk), .Q(data_out[11]), .QN(n185)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n163), .CK(clk), .Q(data_out[10]), .QN(n184)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n164), .CK(clk), .Q(data_out[9]), .QN(n183) );
  DFF_X1 \data_out_reg[8]  ( .D(n165), .CK(clk), .Q(data_out[8]), .QN(n182) );
  DFF_X1 \data_out_reg[7]  ( .D(n166), .CK(clk), .Q(data_out[7]), .QN(n181) );
  DFF_X1 \data_out_reg[6]  ( .D(n167), .CK(clk), .Q(data_out[6]), .QN(n180) );
  DFF_X1 \data_out_reg[5]  ( .D(n168), .CK(clk), .Q(data_out[5]), .QN(n179) );
  DFF_X1 \data_out_reg[4]  ( .D(n169), .CK(clk), .Q(data_out[4]), .QN(n178) );
  DFF_X1 \data_out_reg[3]  ( .D(n170), .CK(clk), .Q(data_out[3]), .QN(n177) );
  DFF_X1 \data_out_reg[2]  ( .D(n171), .CK(clk), .Q(data_out[2]), .QN(n176) );
  DFF_X1 \data_out_reg[1]  ( .D(n172), .CK(clk), .Q(data_out[1]), .QN(n175) );
  DFF_X1 \data_out_reg[0]  ( .D(n173), .CK(clk), .Q(data_out[0]), .QN(n174) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_10_DW_mult_tc_1 mult_2021 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_10_DW01_add_2 add_2022 ( .A({
        n196, n195, n194, n193, n192, n191, n205, n204, n203, n202, n201, n200, 
        n199, n198, n197, n190}), .B({f[15], n41, n42, n44, n45, n47, f[9:0]}), 
        .CI(1'b0), .SUM(adder) );
  DFF_X1 \f_reg[4]  ( .D(n79), .CK(clk), .Q(f[4]), .QN(n60) );
  DFF_X1 \f_reg[5]  ( .D(n78), .CK(clk), .Q(f[5]), .QN(n61) );
  DFF_X1 \f_reg[6]  ( .D(n77), .CK(clk), .Q(f[6]), .QN(n62) );
  DFF_X2 delay_reg ( .D(n85), .CK(clk), .Q(n14), .QN(n234) );
  MUX2_X2 U3 ( .A(N37), .B(n27), .S(n14), .Z(n204) );
  MUX2_X2 U4 ( .A(n21), .B(N43), .S(n234), .Z(n195) );
  MUX2_X1 U5 ( .A(n22), .B(N42), .S(n234), .Z(n194) );
  AND2_X1 U6 ( .A1(clear_acc_delay), .A2(n234), .ZN(n1) );
  AND2_X1 U8 ( .A1(n40), .A2(n18), .ZN(n15) );
  NAND3_X1 U9 ( .A1(n6), .A2(n5), .A3(n7), .ZN(n2) );
  NAND3_X1 U10 ( .A1(n12), .A2(n13), .A3(n11), .ZN(n70) );
  NAND3_X1 U11 ( .A1(n9), .A2(n8), .A3(n10), .ZN(n4) );
  NAND2_X1 U12 ( .A1(data_out_b[12]), .A2(n17), .ZN(n5) );
  NAND2_X1 U13 ( .A1(adder[12]), .A2(n15), .ZN(n6) );
  NAND2_X1 U14 ( .A1(n58), .A2(n44), .ZN(n7) );
  MUX2_X1 U15 ( .A(N38), .B(n26), .S(n14), .Z(n205) );
  NAND2_X1 U16 ( .A1(data_out_b[14]), .A2(n17), .ZN(n8) );
  NAND2_X1 U17 ( .A1(adder[14]), .A2(n15), .ZN(n9) );
  NAND2_X1 U18 ( .A1(n58), .A2(n41), .ZN(n10) );
  MUX2_X2 U19 ( .A(n24), .B(N40), .S(n234), .Z(n192) );
  MUX2_X1 U20 ( .A(N39), .B(n25), .S(n14), .Z(n191) );
  MUX2_X2 U21 ( .A(n23), .B(N41), .S(n234), .Z(n193) );
  NAND2_X1 U22 ( .A1(data_out_b[15]), .A2(n17), .ZN(n11) );
  NAND2_X1 U23 ( .A1(adder[15]), .A2(n15), .ZN(n12) );
  NAND2_X1 U24 ( .A1(n58), .A2(f[15]), .ZN(n13) );
  NAND2_X1 U25 ( .A1(n85), .A2(n16), .ZN(n236) );
  INV_X1 U26 ( .A(n40), .ZN(n58) );
  INV_X1 U27 ( .A(clear_acc), .ZN(n18) );
  OAI22_X1 U28 ( .A1(n177), .A2(n236), .B1(n209), .B2(n235), .ZN(n170) );
  OAI22_X1 U29 ( .A1(n178), .A2(n236), .B1(n60), .B2(n235), .ZN(n169) );
  OAI22_X1 U30 ( .A1(n179), .A2(n236), .B1(n61), .B2(n235), .ZN(n168) );
  OAI22_X1 U31 ( .A1(n180), .A2(n236), .B1(n62), .B2(n235), .ZN(n167) );
  OAI22_X1 U32 ( .A1(n181), .A2(n236), .B1(n210), .B2(n235), .ZN(n166) );
  OAI22_X1 U33 ( .A1(n182), .A2(n236), .B1(n211), .B2(n235), .ZN(n165) );
  OAI22_X1 U34 ( .A1(n183), .A2(n236), .B1(n212), .B2(n235), .ZN(n164) );
  INV_X1 U35 ( .A(wr_en_y), .ZN(n16) );
  INV_X1 U36 ( .A(n18), .ZN(n17) );
  INV_X1 U37 ( .A(m_ready), .ZN(n19) );
  NAND2_X1 U38 ( .A1(m_valid), .A2(n19), .ZN(n38) );
  OAI21_X1 U39 ( .B1(sel[4]), .B2(n69), .A(n38), .ZN(n85) );
  MUX2_X1 U40 ( .A(n20), .B(N44), .S(n1), .Z(n218) );
  MUX2_X1 U41 ( .A(n20), .B(N44), .S(n234), .Z(n196) );
  MUX2_X1 U42 ( .A(n21), .B(N43), .S(n1), .Z(n219) );
  MUX2_X1 U43 ( .A(n22), .B(N42), .S(n1), .Z(n220) );
  MUX2_X1 U44 ( .A(n23), .B(N41), .S(n1), .Z(n221) );
  MUX2_X1 U45 ( .A(n24), .B(N40), .S(n1), .Z(n222) );
  MUX2_X1 U46 ( .A(n25), .B(N39), .S(n1), .Z(n223) );
  MUX2_X1 U47 ( .A(n26), .B(N38), .S(n1), .Z(n224) );
  MUX2_X1 U48 ( .A(n27), .B(N37), .S(n1), .Z(n225) );
  MUX2_X1 U49 ( .A(n28), .B(N36), .S(n1), .Z(n226) );
  MUX2_X1 U50 ( .A(n28), .B(N36), .S(n234), .Z(n203) );
  MUX2_X1 U51 ( .A(n29), .B(N35), .S(n1), .Z(n227) );
  MUX2_X1 U52 ( .A(n29), .B(N35), .S(n234), .Z(n202) );
  MUX2_X1 U53 ( .A(n32), .B(N34), .S(n1), .Z(n228) );
  MUX2_X1 U54 ( .A(n32), .B(N34), .S(n234), .Z(n201) );
  MUX2_X1 U55 ( .A(n33), .B(N33), .S(n1), .Z(n229) );
  MUX2_X1 U56 ( .A(n33), .B(N33), .S(n234), .Z(n200) );
  MUX2_X1 U57 ( .A(n34), .B(N32), .S(n1), .Z(n230) );
  MUX2_X1 U58 ( .A(n34), .B(N32), .S(n234), .Z(n199) );
  MUX2_X1 U59 ( .A(n35), .B(N31), .S(n1), .Z(n231) );
  MUX2_X1 U60 ( .A(n35), .B(N31), .S(n234), .Z(n198) );
  MUX2_X1 U61 ( .A(n36), .B(N30), .S(n1), .Z(n232) );
  MUX2_X1 U62 ( .A(n36), .B(N30), .S(n234), .Z(n197) );
  MUX2_X1 U63 ( .A(n37), .B(N29), .S(n1), .Z(n233) );
  MUX2_X1 U64 ( .A(n37), .B(N29), .S(n234), .Z(n190) );
  INV_X1 U65 ( .A(n38), .ZN(n39) );
  OAI21_X1 U66 ( .B1(n39), .B2(n14), .A(n18), .ZN(n40) );
  AOI222_X1 U67 ( .A1(data_out_b[13]), .A2(n17), .B1(adder[13]), .B2(n15), 
        .C1(n58), .C2(n42), .ZN(n43) );
  INV_X1 U68 ( .A(n43), .ZN(n71) );
  AOI222_X1 U69 ( .A1(data_out_b[11]), .A2(n17), .B1(adder[11]), .B2(n15), 
        .C1(n58), .C2(n45), .ZN(n46) );
  INV_X1 U70 ( .A(n46), .ZN(n72) );
  AOI222_X1 U71 ( .A1(data_out_b[10]), .A2(n17), .B1(adder[10]), .B2(n15), 
        .C1(n58), .C2(n47), .ZN(n48) );
  INV_X1 U72 ( .A(n48), .ZN(n73) );
  AOI222_X1 U73 ( .A1(data_out_b[8]), .A2(n17), .B1(adder[8]), .B2(n15), .C1(
        n58), .C2(f[8]), .ZN(n49) );
  INV_X1 U74 ( .A(n49), .ZN(n75) );
  AOI222_X1 U75 ( .A1(data_out_b[7]), .A2(n17), .B1(adder[7]), .B2(n15), .C1(
        n58), .C2(f[7]), .ZN(n50) );
  INV_X1 U76 ( .A(n50), .ZN(n76) );
  AOI222_X1 U77 ( .A1(data_out_b[6]), .A2(n17), .B1(adder[6]), .B2(n15), .C1(
        n58), .C2(f[6]), .ZN(n51) );
  INV_X1 U78 ( .A(n51), .ZN(n77) );
  AOI222_X1 U79 ( .A1(data_out_b[5]), .A2(n17), .B1(adder[5]), .B2(n15), .C1(
        n58), .C2(f[5]), .ZN(n52) );
  INV_X1 U80 ( .A(n52), .ZN(n78) );
  AOI222_X1 U81 ( .A1(data_out_b[4]), .A2(n17), .B1(adder[4]), .B2(n15), .C1(
        n58), .C2(f[4]), .ZN(n53) );
  INV_X1 U82 ( .A(n53), .ZN(n79) );
  AOI222_X1 U83 ( .A1(data_out_b[3]), .A2(n17), .B1(adder[3]), .B2(n15), .C1(
        n58), .C2(f[3]), .ZN(n54) );
  INV_X1 U84 ( .A(n54), .ZN(n80) );
  AOI222_X1 U85 ( .A1(data_out_b[2]), .A2(n17), .B1(adder[2]), .B2(n15), .C1(
        n58), .C2(f[2]), .ZN(n55) );
  INV_X1 U86 ( .A(n55), .ZN(n81) );
  AOI222_X1 U87 ( .A1(data_out_b[1]), .A2(n17), .B1(adder[1]), .B2(n15), .C1(
        n58), .C2(f[1]), .ZN(n56) );
  INV_X1 U88 ( .A(n56), .ZN(n82) );
  AOI222_X1 U89 ( .A1(data_out_b[0]), .A2(n17), .B1(adder[0]), .B2(n15), .C1(
        n58), .C2(f[0]), .ZN(n57) );
  INV_X1 U90 ( .A(n57), .ZN(n83) );
  AOI222_X1 U91 ( .A1(data_out_b[9]), .A2(n17), .B1(adder[9]), .B2(n15), .C1(
        n58), .C2(f[9]), .ZN(n59) );
  INV_X1 U92 ( .A(n59), .ZN(n74) );
  NOR4_X1 U93 ( .A1(n45), .A2(n44), .A3(n42), .A4(n41), .ZN(n66) );
  NOR4_X1 U94 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n47), .ZN(n65) );
  NAND4_X1 U95 ( .A1(n62), .A2(n61), .A3(n60), .A4(n209), .ZN(n63) );
  NOR4_X1 U96 ( .A1(n63), .A2(f[0]), .A3(f[1]), .A4(f[2]), .ZN(n64) );
  NAND3_X1 U97 ( .A1(n66), .A2(n65), .A3(n64), .ZN(n68) );
  NAND3_X1 U98 ( .A1(wr_en_y), .A2(n68), .A3(n67), .ZN(n235) );
  OAI22_X1 U99 ( .A1(n174), .A2(n236), .B1(n206), .B2(n235), .ZN(n173) );
  OAI22_X1 U100 ( .A1(n175), .A2(n236), .B1(n207), .B2(n235), .ZN(n172) );
  OAI22_X1 U101 ( .A1(n176), .A2(n236), .B1(n208), .B2(n235), .ZN(n171) );
  OAI22_X1 U102 ( .A1(n184), .A2(n236), .B1(n213), .B2(n235), .ZN(n163) );
  OAI22_X1 U103 ( .A1(n185), .A2(n236), .B1(n214), .B2(n235), .ZN(n162) );
  OAI22_X1 U104 ( .A1(n186), .A2(n236), .B1(n215), .B2(n235), .ZN(n113) );
  OAI22_X1 U105 ( .A1(n187), .A2(n236), .B1(n216), .B2(n235), .ZN(n112) );
  OAI22_X1 U106 ( .A1(n188), .A2(n236), .B1(n217), .B2(n235), .ZN(n111) );
  OAI22_X1 U107 ( .A1(n189), .A2(n236), .B1(n67), .B2(n235), .ZN(n102) );
  AND4_X1 U108 ( .A1(sel[3]), .A2(sel[2]), .A3(sel[1]), .A4(sel[0]), .ZN(n69)
         );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_9_DW_mult_tc_1 ( a, b, 
        product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n9, n12, n13, n16, n18, n19, n21, n23, n25, n27, n29, n31,
         n32, n34, n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n50,
         n53, n54, n55, n56, n57, n58, n59, n62, n63, n64, n65, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n93, n95, n96, n97, n98, n99, n101,
         n103, n104, n105, n106, n107, n111, n112, n113, n114, n115, n117,
         n119, n120, n122, n125, n131, n135, n139, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n245, n247, n249, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n418, n419,
         n420, n421, n422, n423, n424, n426, n427, n429, n431, n432, n433,
         n490, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U148 ( .A(n265), .B(n144), .Z(n145) );
  XOR2_X1 U150 ( .A(n271), .B(n146), .Z(n147) );
  XOR2_X1 U152 ( .A(n301), .B(n148), .Z(n149) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U162 ( .A(n170), .B(n172), .CI(n179), .CO(n165), .S(n166) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n263), .CI(n291), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n317), .B(n252), .CO(n173), .S(n174) );
  FA_X1 U167 ( .A(n180), .B(n187), .CI(n178), .CO(n175), .S(n176) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U169 ( .A(n193), .B(n282), .CI(n191), .CO(n179), .S(n180) );
  FA_X1 U170 ( .A(n268), .B(n292), .CI(n274), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U172 ( .A(n197), .B(n190), .CI(n188), .CO(n185), .S(n186) );
  FA_X1 U173 ( .A(n199), .B(n201), .CI(n192), .CO(n187), .S(n188) );
  FA_X1 U174 ( .A(n275), .B(n293), .CI(n194), .CO(n189), .S(n190) );
  FA_X1 U175 ( .A(n305), .B(n253), .CI(n283), .CO(n191), .S(n192) );
  HA_X1 U176 ( .A(n269), .B(n319), .CO(n193), .S(n194) );
  FA_X1 U177 ( .A(n205), .B(n200), .CI(n198), .CO(n195), .S(n196) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U179 ( .A(n276), .B(n284), .CI(n294), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n320), .B(n270), .CI(n306), .CO(n201), .S(n202) );
  FA_X1 U181 ( .A(n208), .B(n213), .CI(n206), .CO(n203), .S(n204) );
  FA_X1 U182 ( .A(n215), .B(n307), .CI(n210), .CO(n205), .S(n206) );
  FA_X1 U183 ( .A(n295), .B(n285), .CI(n254), .CO(n207), .S(n208) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U185 ( .A(n216), .B(n219), .CI(n214), .CO(n211), .S(n212) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n322), .B(n278), .CI(n308), .CO(n215), .S(n216) );
  FA_X1 U188 ( .A(n225), .B(n222), .CI(n220), .CO(n217), .S(n218) );
  FA_X1 U189 ( .A(n255), .B(n309), .CI(n297), .CO(n219), .S(n220) );
  HA_X1 U190 ( .A(n287), .B(n323), .CO(n221), .S(n222) );
  FA_X1 U192 ( .A(n324), .B(n288), .CI(n310), .CO(n225), .S(n226) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  HA_X1 U194 ( .A(n311), .B(n325), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n326), .B(n300), .CI(n312), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  BUF_X1 U414 ( .A(n95), .Z(n490) );
  INV_X1 U415 ( .A(n502), .ZN(n41) );
  BUF_X1 U416 ( .A(n16), .Z(n567) );
  INV_X1 U417 ( .A(n499), .ZN(n516) );
  AND2_X1 U418 ( .A1(n492), .A2(n122), .ZN(product[1]) );
  OR2_X1 U419 ( .A1(n329), .A2(n258), .ZN(n492) );
  XNOR2_X1 U420 ( .A(n581), .B(a[6]), .ZN(n493) );
  OR2_X2 U421 ( .A1(n545), .A2(n557), .ZN(n494) );
  CLKBUF_X1 U422 ( .A(n532), .Z(n495) );
  XNOR2_X2 U423 ( .A(n501), .B(a[2]), .ZN(n432) );
  OAI21_X1 U424 ( .B1(n113), .B2(n115), .A(n114), .ZN(n112) );
  AND2_X1 U425 ( .A1(n232), .A2(n233), .ZN(n496) );
  OR2_X1 U426 ( .A1(n196), .A2(n203), .ZN(n497) );
  XNOR2_X1 U427 ( .A(n226), .B(n498), .ZN(n224) );
  XNOR2_X1 U428 ( .A(n229), .B(n298), .ZN(n498) );
  NOR2_X1 U429 ( .A1(n196), .A2(n203), .ZN(n85) );
  XNOR2_X1 U430 ( .A(a[8]), .B(n583), .ZN(n499) );
  INV_X1 U431 ( .A(n19), .ZN(n583) );
  INV_X1 U432 ( .A(n575), .ZN(n574) );
  INV_X1 U433 ( .A(n575), .ZN(n500) );
  INV_X1 U434 ( .A(n7), .ZN(n501) );
  INV_X1 U435 ( .A(n520), .ZN(n37) );
  XNOR2_X1 U436 ( .A(n589), .B(a[14]), .ZN(n502) );
  BUF_X1 U437 ( .A(n581), .Z(n503) );
  INV_X1 U438 ( .A(n517), .ZN(n504) );
  INV_X1 U439 ( .A(n584), .ZN(n505) );
  AND2_X1 U440 ( .A1(n535), .A2(n536), .ZN(n506) );
  AND2_X1 U441 ( .A1(n535), .A2(n536), .ZN(n556) );
  XNOR2_X1 U442 ( .A(n585), .B(a[8]), .ZN(n429) );
  INV_X1 U443 ( .A(n575), .ZN(n569) );
  NOR2_X1 U444 ( .A1(n575), .A2(n507), .ZN(n539) );
  INV_X1 U445 ( .A(a[2]), .ZN(n507) );
  AOI21_X1 U446 ( .B1(n96), .B2(n559), .A(n93), .ZN(n508) );
  AOI21_X1 U447 ( .B1(n96), .B2(n559), .A(n93), .ZN(n91) );
  XNOR2_X1 U448 ( .A(n45), .B(n509), .ZN(product[12]) );
  AND2_X1 U449 ( .A1(n531), .A2(n79), .ZN(n509) );
  XNOR2_X1 U450 ( .A(n513), .B(n510), .ZN(product[9]) );
  AND2_X1 U451 ( .A1(n528), .A2(n90), .ZN(n510) );
  INV_X1 U452 ( .A(n585), .ZN(n511) );
  CLKBUF_X1 U453 ( .A(n186), .Z(n512) );
  CLKBUF_X1 U454 ( .A(n508), .Z(n513) );
  CLKBUF_X1 U455 ( .A(n21), .Z(n514) );
  INV_X1 U456 ( .A(n577), .ZN(n515) );
  INV_X2 U457 ( .A(n501), .ZN(n577) );
  XOR2_X1 U458 ( .A(a[8]), .B(n583), .Z(n27) );
  INV_X1 U459 ( .A(n587), .ZN(n517) );
  INV_X1 U460 ( .A(n585), .ZN(n518) );
  INV_X1 U461 ( .A(n585), .ZN(n584) );
  CLKBUF_X1 U462 ( .A(n104), .Z(n519) );
  XNOR2_X1 U463 ( .A(n587), .B(a[12]), .ZN(n520) );
  INV_X1 U464 ( .A(n587), .ZN(n586) );
  OR2_X2 U465 ( .A1(n521), .A2(n549), .ZN(n34) );
  XNOR2_X1 U466 ( .A(n31), .B(a[10]), .ZN(n521) );
  INV_X1 U467 ( .A(n549), .ZN(n32) );
  NAND2_X1 U468 ( .A1(n9), .A2(n432), .ZN(n522) );
  NAND2_X1 U469 ( .A1(n432), .A2(n9), .ZN(n523) );
  OR2_X2 U470 ( .A1(n540), .A2(n539), .ZN(n9) );
  XNOR2_X1 U471 ( .A(n503), .B(a[4]), .ZN(n431) );
  INV_X1 U472 ( .A(n581), .ZN(n579) );
  INV_X1 U473 ( .A(n247), .ZN(n524) );
  CLKBUF_X1 U474 ( .A(n107), .Z(n525) );
  AOI21_X1 U475 ( .B1(n562), .B2(n112), .A(n496), .ZN(n107) );
  XOR2_X1 U476 ( .A(n583), .B(a[6]), .Z(n545) );
  CLKBUF_X3 U477 ( .A(n16), .Z(n568) );
  NAND2_X1 U478 ( .A1(n431), .A2(n567), .ZN(n526) );
  NAND2_X1 U479 ( .A1(n431), .A2(n567), .ZN(n527) );
  NAND2_X1 U480 ( .A1(n431), .A2(n567), .ZN(n18) );
  OR2_X1 U481 ( .A1(n204), .A2(n211), .ZN(n528) );
  XNOR2_X1 U482 ( .A(n166), .B(n529), .ZN(n164) );
  XNOR2_X1 U483 ( .A(n177), .B(n168), .ZN(n529) );
  NOR2_X1 U484 ( .A1(n195), .A2(n186), .ZN(n530) );
  OR2_X1 U485 ( .A1(n176), .A2(n185), .ZN(n531) );
  OR2_X2 U486 ( .A1(n539), .A2(n540), .ZN(n532) );
  OR2_X1 U487 ( .A1(n228), .A2(n231), .ZN(n533) );
  XNOR2_X1 U488 ( .A(n88), .B(n534), .ZN(product[10]) );
  NAND2_X1 U489 ( .A1(n497), .A2(n86), .ZN(n534) );
  NAND2_X1 U490 ( .A1(n537), .A2(n80), .ZN(n535) );
  INV_X1 U491 ( .A(n81), .ZN(n536) );
  OAI21_X1 U492 ( .B1(n91), .B2(n89), .A(n90), .ZN(n537) );
  CLKBUF_X1 U493 ( .A(n96), .Z(n538) );
  AND2_X1 U494 ( .A1(n575), .A2(n553), .ZN(n540) );
  OR2_X1 U495 ( .A1(n512), .A2(n195), .ZN(n541) );
  NAND2_X1 U496 ( .A1(n166), .A2(n177), .ZN(n542) );
  NAND2_X1 U497 ( .A1(n166), .A2(n168), .ZN(n543) );
  NAND2_X1 U498 ( .A1(n177), .A2(n168), .ZN(n544) );
  NAND3_X1 U499 ( .A1(n542), .A2(n543), .A3(n544), .ZN(n163) );
  INV_X1 U500 ( .A(n578), .ZN(n576) );
  XNOR2_X1 U501 ( .A(n575), .B(n249), .ZN(n433) );
  XOR2_X1 U502 ( .A(n578), .B(a[4]), .Z(n16) );
  OR2_X2 U503 ( .A1(n545), .A2(n557), .ZN(n23) );
  INV_X1 U504 ( .A(n493), .ZN(n21) );
  OAI22_X1 U505 ( .A1(n527), .A2(n375), .B1(n374), .B2(n568), .ZN(n298) );
  NAND2_X2 U506 ( .A1(n429), .A2(n27), .ZN(n29) );
  CLKBUF_X1 U507 ( .A(n99), .Z(n546) );
  NAND2_X1 U508 ( .A1(n432), .A2(n9), .ZN(n547) );
  NAND2_X1 U509 ( .A1(n9), .A2(n432), .ZN(n548) );
  NAND2_X1 U510 ( .A1(n432), .A2(n9), .ZN(n12) );
  NOR2_X2 U511 ( .A1(n164), .A2(n175), .ZN(n75) );
  XNOR2_X1 U512 ( .A(n585), .B(a[10]), .ZN(n549) );
  INV_X2 U513 ( .A(n249), .ZN(n573) );
  NAND2_X1 U514 ( .A1(n226), .A2(n229), .ZN(n550) );
  NAND2_X1 U515 ( .A1(n226), .A2(n298), .ZN(n551) );
  NAND2_X1 U516 ( .A1(n229), .A2(n298), .ZN(n552) );
  NAND3_X1 U517 ( .A1(n550), .A2(n551), .A3(n552), .ZN(n223) );
  INV_X2 U518 ( .A(n583), .ZN(n582) );
  INV_X1 U519 ( .A(a[2]), .ZN(n553) );
  NAND2_X1 U520 ( .A1(n433), .A2(n573), .ZN(n554) );
  NAND2_X1 U521 ( .A1(n433), .A2(n573), .ZN(n555) );
  BUF_X1 U522 ( .A(n43), .Z(n571) );
  XNOR2_X1 U523 ( .A(n581), .B(a[6]), .ZN(n557) );
  NAND2_X1 U524 ( .A1(n558), .A2(n69), .ZN(n47) );
  INV_X1 U525 ( .A(n73), .ZN(n71) );
  AOI21_X1 U526 ( .B1(n74), .B2(n558), .A(n67), .ZN(n65) );
  INV_X1 U527 ( .A(n69), .ZN(n67) );
  INV_X1 U528 ( .A(n74), .ZN(n72) );
  NAND2_X1 U529 ( .A1(n73), .A2(n558), .ZN(n64) );
  INV_X1 U530 ( .A(n95), .ZN(n93) );
  AOI21_X1 U531 ( .B1(n80), .B2(n88), .A(n81), .ZN(n45) );
  NOR2_X1 U532 ( .A1(n530), .A2(n85), .ZN(n80) );
  OAI21_X1 U533 ( .B1(n86), .B2(n82), .A(n83), .ZN(n81) );
  OR2_X1 U534 ( .A1(n152), .A2(n163), .ZN(n558) );
  OAI21_X1 U535 ( .B1(n75), .B2(n79), .A(n76), .ZN(n74) );
  NAND2_X1 U536 ( .A1(n541), .A2(n83), .ZN(n50) );
  NAND2_X1 U537 ( .A1(n125), .A2(n76), .ZN(n48) );
  INV_X1 U538 ( .A(n75), .ZN(n125) );
  NOR2_X1 U539 ( .A1(n75), .A2(n78), .ZN(n73) );
  NAND2_X1 U540 ( .A1(n152), .A2(n163), .ZN(n69) );
  NAND2_X1 U541 ( .A1(n559), .A2(n490), .ZN(n53) );
  INV_X1 U542 ( .A(n103), .ZN(n101) );
  INV_X1 U543 ( .A(n113), .ZN(n135) );
  NOR2_X1 U544 ( .A1(n186), .A2(n195), .ZN(n82) );
  NAND2_X1 U545 ( .A1(n131), .A2(n98), .ZN(n54) );
  INV_X1 U546 ( .A(n97), .ZN(n131) );
  NOR2_X1 U547 ( .A1(n176), .A2(n185), .ZN(n78) );
  NAND2_X1 U548 ( .A1(n560), .A2(n103), .ZN(n55) );
  AOI21_X1 U549 ( .B1(n563), .B2(n120), .A(n117), .ZN(n115) );
  INV_X1 U550 ( .A(n119), .ZN(n117) );
  OAI21_X1 U551 ( .B1(n99), .B2(n97), .A(n98), .ZN(n96) );
  INV_X1 U552 ( .A(n122), .ZN(n120) );
  XNOR2_X1 U553 ( .A(n57), .B(n112), .ZN(product[4]) );
  NAND2_X1 U554 ( .A1(n562), .A2(n111), .ZN(n57) );
  NAND2_X1 U555 ( .A1(n176), .A2(n185), .ZN(n79) );
  NAND2_X1 U556 ( .A1(n186), .A2(n195), .ZN(n83) );
  NAND2_X1 U557 ( .A1(n164), .A2(n175), .ZN(n76) );
  NAND2_X1 U558 ( .A1(n196), .A2(n203), .ZN(n86) );
  NAND2_X1 U559 ( .A1(n212), .A2(n217), .ZN(n95) );
  OR2_X1 U560 ( .A1(n212), .A2(n217), .ZN(n559) );
  XNOR2_X1 U561 ( .A(n59), .B(n120), .ZN(product[2]) );
  NAND2_X1 U562 ( .A1(n563), .A2(n119), .ZN(n59) );
  NAND2_X1 U563 ( .A1(n533), .A2(n106), .ZN(n56) );
  OR2_X1 U564 ( .A1(n224), .A2(n227), .ZN(n560) );
  OR2_X1 U565 ( .A1(n151), .A2(n139), .ZN(n561) );
  NAND2_X1 U566 ( .A1(n328), .A2(n314), .ZN(n119) );
  OR2_X1 U567 ( .A1(n232), .A2(n233), .ZN(n562) );
  NOR2_X1 U568 ( .A1(n218), .A2(n223), .ZN(n97) );
  NOR2_X1 U569 ( .A1(n234), .A2(n257), .ZN(n113) );
  XNOR2_X1 U570 ( .A(n63), .B(n46), .ZN(product[15]) );
  NAND2_X1 U571 ( .A1(n561), .A2(n62), .ZN(n46) );
  OR2_X1 U572 ( .A1(n328), .A2(n314), .ZN(n563) );
  NOR2_X1 U573 ( .A1(n228), .A2(n231), .ZN(n105) );
  NAND2_X1 U574 ( .A1(n218), .A2(n223), .ZN(n98) );
  NAND2_X1 U575 ( .A1(n228), .A2(n231), .ZN(n106) );
  NAND2_X1 U576 ( .A1(n224), .A2(n227), .ZN(n103) );
  NAND2_X1 U577 ( .A1(n232), .A2(n233), .ZN(n111) );
  OR2_X1 U578 ( .A1(n571), .A2(n570), .ZN(n409) );
  OR2_X1 U579 ( .A1(n571), .A2(n515), .ZN(n392) );
  NAND2_X1 U580 ( .A1(n433), .A2(n573), .ZN(n6) );
  XNOR2_X1 U581 ( .A(n511), .B(n571), .ZN(n352) );
  AND2_X1 U582 ( .A1(n572), .A2(n245), .ZN(n300) );
  AND2_X1 U583 ( .A1(n572), .A2(n493), .ZN(n288) );
  AND2_X1 U584 ( .A1(n572), .A2(n499), .ZN(n278) );
  AND2_X1 U585 ( .A1(n572), .A2(n549), .ZN(n270) );
  XNOR2_X1 U586 ( .A(n580), .B(n571), .ZN(n376) );
  XNOR2_X1 U587 ( .A(n155), .B(n564), .ZN(n139) );
  XNOR2_X1 U588 ( .A(n153), .B(n141), .ZN(n564) );
  XNOR2_X1 U589 ( .A(n157), .B(n565), .ZN(n141) );
  XNOR2_X1 U590 ( .A(n145), .B(n143), .ZN(n565) );
  OAI22_X1 U591 ( .A1(n39), .A2(n589), .B1(n337), .B2(n37), .ZN(n252) );
  OR2_X1 U592 ( .A1(n571), .A2(n589), .ZN(n337) );
  OAI22_X1 U593 ( .A1(n42), .A2(n591), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U594 ( .A1(n571), .A2(n591), .ZN(n332) );
  XNOR2_X1 U595 ( .A(n586), .B(n571), .ZN(n343) );
  XNOR2_X1 U596 ( .A(n159), .B(n566), .ZN(n142) );
  XNOR2_X1 U597 ( .A(n315), .B(n261), .ZN(n566) );
  XNOR2_X1 U598 ( .A(n588), .B(n571), .ZN(n336) );
  AND2_X1 U599 ( .A1(n572), .A2(n247), .ZN(n314) );
  NAND2_X1 U600 ( .A1(n427), .A2(n37), .ZN(n39) );
  XOR2_X1 U601 ( .A(n588), .B(a[12]), .Z(n427) );
  OAI22_X1 U602 ( .A1(n39), .A2(n336), .B1(n37), .B2(n335), .ZN(n263) );
  AND2_X1 U603 ( .A1(n572), .A2(n520), .ZN(n264) );
  AND2_X1 U604 ( .A1(n572), .A2(n502), .ZN(n260) );
  OAI22_X1 U605 ( .A1(n39), .A2(n335), .B1(n37), .B2(n334), .ZN(n262) );
  INV_X1 U606 ( .A(n25), .ZN(n585) );
  NAND2_X1 U607 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U608 ( .A(n590), .B(a[14]), .Z(n426) );
  INV_X1 U609 ( .A(n7), .ZN(n578) );
  XNOR2_X1 U610 ( .A(n582), .B(n571), .ZN(n363) );
  AND2_X1 U611 ( .A1(n572), .A2(n249), .ZN(product[0]) );
  OR2_X1 U612 ( .A1(n571), .A2(n583), .ZN(n364) );
  OR2_X1 U613 ( .A1(n571), .A2(n504), .ZN(n344) );
  OR2_X1 U614 ( .A1(n571), .A2(n505), .ZN(n353) );
  OR2_X1 U615 ( .A1(n571), .A2(n503), .ZN(n377) );
  XNOR2_X1 U616 ( .A(n582), .B(b[9]), .ZN(n354) );
  OAI22_X1 U617 ( .A1(n39), .A2(n334), .B1(n37), .B2(n333), .ZN(n261) );
  XNOR2_X1 U618 ( .A(n588), .B(n422), .ZN(n333) );
  XNOR2_X1 U619 ( .A(n580), .B(b[11]), .ZN(n365) );
  XNOR2_X1 U620 ( .A(n588), .B(n423), .ZN(n334) );
  XNOR2_X1 U621 ( .A(n588), .B(n424), .ZN(n335) );
  OAI22_X1 U622 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U623 ( .A(n590), .B(n424), .ZN(n330) );
  XNOR2_X1 U624 ( .A(n590), .B(n571), .ZN(n331) );
  XNOR2_X1 U625 ( .A(n518), .B(n418), .ZN(n345) );
  XNOR2_X1 U626 ( .A(n517), .B(n420), .ZN(n338) );
  XNOR2_X1 U627 ( .A(n577), .B(b[13]), .ZN(n378) );
  XNOR2_X1 U628 ( .A(n586), .B(n424), .ZN(n342) );
  XNOR2_X1 U629 ( .A(n582), .B(n424), .ZN(n362) );
  XNOR2_X1 U630 ( .A(n584), .B(n424), .ZN(n351) );
  XNOR2_X1 U631 ( .A(n586), .B(n423), .ZN(n341) );
  XNOR2_X1 U632 ( .A(n517), .B(n422), .ZN(n340) );
  XNOR2_X1 U633 ( .A(n517), .B(n421), .ZN(n339) );
  XNOR2_X1 U634 ( .A(n577), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U635 ( .A(n577), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U636 ( .A(n577), .B(n418), .ZN(n384) );
  XNOR2_X1 U637 ( .A(n577), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U638 ( .A(n577), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U639 ( .A(n577), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U640 ( .A(n577), .B(n419), .ZN(n385) );
  XNOR2_X1 U641 ( .A(n582), .B(n423), .ZN(n361) );
  XNOR2_X1 U642 ( .A(n511), .B(n423), .ZN(n350) );
  XNOR2_X1 U643 ( .A(n580), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U644 ( .A(n580), .B(n418), .ZN(n369) );
  XNOR2_X1 U645 ( .A(n580), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U646 ( .A(n580), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U647 ( .A(n582), .B(n422), .ZN(n360) );
  XNOR2_X1 U648 ( .A(n518), .B(n422), .ZN(n349) );
  XNOR2_X1 U649 ( .A(n582), .B(n421), .ZN(n359) );
  XNOR2_X1 U650 ( .A(n584), .B(n421), .ZN(n348) );
  XNOR2_X1 U651 ( .A(n582), .B(n420), .ZN(n358) );
  XNOR2_X1 U652 ( .A(n518), .B(n420), .ZN(n347) );
  XNOR2_X1 U653 ( .A(n582), .B(n418), .ZN(n356) );
  XNOR2_X1 U654 ( .A(n582), .B(n419), .ZN(n357) );
  XNOR2_X1 U655 ( .A(n518), .B(n419), .ZN(n346) );
  XNOR2_X1 U656 ( .A(n582), .B(b[8]), .ZN(n355) );
  XNOR2_X1 U657 ( .A(n500), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U658 ( .A(n500), .B(b[14]), .ZN(n394) );
  XNOR2_X1 U659 ( .A(n500), .B(b[11]), .ZN(n397) );
  XNOR2_X1 U660 ( .A(n574), .B(b[13]), .ZN(n395) );
  BUF_X1 U661 ( .A(n43), .Z(n572) );
  XNOR2_X1 U662 ( .A(n500), .B(b[15]), .ZN(n393) );
  OAI22_X1 U663 ( .A1(n34), .A2(n339), .B1(n338), .B2(n32), .ZN(n265) );
  OAI22_X1 U664 ( .A1(n34), .A2(n340), .B1(n339), .B2(n32), .ZN(n266) );
  OAI22_X1 U665 ( .A1(n34), .A2(n341), .B1(n340), .B2(n32), .ZN(n267) );
  OAI22_X1 U666 ( .A1(n34), .A2(n342), .B1(n341), .B2(n32), .ZN(n268) );
  OAI22_X1 U667 ( .A1(n34), .A2(n343), .B1(n342), .B2(n32), .ZN(n269) );
  OAI22_X1 U668 ( .A1(n34), .A2(n504), .B1(n344), .B2(n32), .ZN(n253) );
  OAI22_X1 U669 ( .A1(n6), .A2(n395), .B1(n394), .B2(n573), .ZN(n316) );
  OAI22_X1 U670 ( .A1(n6), .A2(n394), .B1(n393), .B2(n573), .ZN(n315) );
  OAI22_X1 U671 ( .A1(n6), .A2(n400), .B1(n399), .B2(n573), .ZN(n321) );
  OAI22_X1 U672 ( .A1(n554), .A2(n401), .B1(n400), .B2(n573), .ZN(n322) );
  OAI22_X1 U673 ( .A1(n6), .A2(n397), .B1(n396), .B2(n573), .ZN(n318) );
  OAI22_X1 U674 ( .A1(n554), .A2(n396), .B1(n395), .B2(n573), .ZN(n317) );
  OAI22_X1 U675 ( .A1(n555), .A2(n398), .B1(n397), .B2(n573), .ZN(n319) );
  OAI22_X1 U676 ( .A1(n555), .A2(n399), .B1(n398), .B2(n573), .ZN(n320) );
  OAI22_X1 U677 ( .A1(n555), .A2(n402), .B1(n401), .B2(n573), .ZN(n323) );
  OAI22_X1 U678 ( .A1(n6), .A2(n406), .B1(n405), .B2(n573), .ZN(n327) );
  OAI22_X1 U679 ( .A1(n554), .A2(n404), .B1(n403), .B2(n573), .ZN(n325) );
  OAI22_X1 U680 ( .A1(n555), .A2(n405), .B1(n404), .B2(n573), .ZN(n326) );
  OAI22_X1 U681 ( .A1(n6), .A2(n403), .B1(n402), .B2(n573), .ZN(n324) );
  OAI22_X1 U682 ( .A1(n555), .A2(n408), .B1(n407), .B2(n573), .ZN(n329) );
  OAI22_X1 U683 ( .A1(n554), .A2(n407), .B1(n406), .B2(n573), .ZN(n328) );
  INV_X1 U684 ( .A(n13), .ZN(n581) );
  INV_X1 U685 ( .A(n569), .ZN(n570) );
  INV_X1 U686 ( .A(n1), .ZN(n575) );
  XNOR2_X1 U687 ( .A(n84), .B(n50), .ZN(product[11]) );
  XNOR2_X1 U688 ( .A(n70), .B(n47), .ZN(product[14]) );
  NAND2_X1 U689 ( .A1(n204), .A2(n211), .ZN(n90) );
  NOR2_X1 U690 ( .A1(n204), .A2(n211), .ZN(n89) );
  OAI22_X1 U691 ( .A1(n29), .A2(n346), .B1(n345), .B2(n516), .ZN(n271) );
  OAI22_X1 U692 ( .A1(n29), .A2(n350), .B1(n349), .B2(n516), .ZN(n275) );
  OAI22_X1 U693 ( .A1(n29), .A2(n347), .B1(n346), .B2(n516), .ZN(n272) );
  OAI22_X1 U694 ( .A1(n29), .A2(n348), .B1(n347), .B2(n516), .ZN(n273) );
  OAI22_X1 U695 ( .A1(n29), .A2(n349), .B1(n348), .B2(n516), .ZN(n274) );
  OAI22_X1 U696 ( .A1(n29), .A2(n505), .B1(n353), .B2(n516), .ZN(n254) );
  OAI22_X1 U697 ( .A1(n29), .A2(n351), .B1(n350), .B2(n516), .ZN(n276) );
  OAI22_X1 U698 ( .A1(n29), .A2(n352), .B1(n351), .B2(n516), .ZN(n277) );
  XNOR2_X1 U699 ( .A(n538), .B(n53), .ZN(product[8]) );
  NAND2_X1 U700 ( .A1(n151), .A2(n139), .ZN(n62) );
  NAND2_X1 U701 ( .A1(n135), .A2(n114), .ZN(n58) );
  XNOR2_X1 U702 ( .A(n579), .B(n424), .ZN(n375) );
  XNOR2_X1 U703 ( .A(n579), .B(n419), .ZN(n370) );
  XNOR2_X1 U704 ( .A(n579), .B(n420), .ZN(n371) );
  XNOR2_X1 U705 ( .A(n579), .B(n423), .ZN(n374) );
  XNOR2_X1 U706 ( .A(n579), .B(n422), .ZN(n373) );
  XNOR2_X1 U707 ( .A(n579), .B(n421), .ZN(n372) );
  XOR2_X1 U708 ( .A(n546), .B(n54), .Z(product[7]) );
  XOR2_X1 U709 ( .A(n58), .B(n115), .Z(product[3]) );
  OAI21_X1 U710 ( .B1(n105), .B2(n107), .A(n106), .ZN(n104) );
  AOI21_X1 U711 ( .B1(n104), .B2(n560), .A(n101), .ZN(n99) );
  XNOR2_X1 U712 ( .A(n55), .B(n519), .ZN(product[6]) );
  XNOR2_X1 U713 ( .A(n77), .B(n48), .ZN(product[13]) );
  XNOR2_X1 U714 ( .A(n569), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U715 ( .A(n574), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U716 ( .A(n569), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U717 ( .A(n574), .B(n418), .ZN(n401) );
  XNOR2_X1 U718 ( .A(n500), .B(n419), .ZN(n402) );
  XNOR2_X1 U719 ( .A(n569), .B(n420), .ZN(n403) );
  XNOR2_X1 U720 ( .A(n574), .B(n571), .ZN(n408) );
  XNOR2_X1 U721 ( .A(n569), .B(n421), .ZN(n404) );
  XNOR2_X1 U722 ( .A(n574), .B(n422), .ZN(n405) );
  XNOR2_X1 U723 ( .A(n500), .B(n424), .ZN(n407) );
  XNOR2_X1 U724 ( .A(n574), .B(n423), .ZN(n406) );
  OAI22_X1 U725 ( .A1(n23), .A2(n356), .B1(n355), .B2(n514), .ZN(n280) );
  OAI22_X1 U726 ( .A1(n494), .A2(n358), .B1(n357), .B2(n514), .ZN(n282) );
  OAI22_X1 U727 ( .A1(n23), .A2(n362), .B1(n361), .B2(n21), .ZN(n286) );
  OAI22_X1 U728 ( .A1(n23), .A2(n360), .B1(n359), .B2(n21), .ZN(n284) );
  OAI22_X1 U729 ( .A1(n23), .A2(n361), .B1(n360), .B2(n21), .ZN(n285) );
  OAI22_X1 U730 ( .A1(n494), .A2(n583), .B1(n364), .B2(n21), .ZN(n255) );
  OAI22_X1 U731 ( .A1(n494), .A2(n357), .B1(n356), .B2(n21), .ZN(n281) );
  OAI22_X1 U732 ( .A1(n494), .A2(n355), .B1(n354), .B2(n21), .ZN(n279) );
  OAI22_X1 U733 ( .A1(n23), .A2(n363), .B1(n362), .B2(n21), .ZN(n287) );
  OAI22_X1 U734 ( .A1(n494), .A2(n359), .B1(n358), .B2(n21), .ZN(n283) );
  OAI22_X1 U735 ( .A1(n527), .A2(n370), .B1(n369), .B2(n568), .ZN(n293) );
  OAI22_X1 U736 ( .A1(n526), .A2(n367), .B1(n366), .B2(n568), .ZN(n290) );
  OAI22_X1 U737 ( .A1(n18), .A2(n372), .B1(n371), .B2(n568), .ZN(n295) );
  OAI22_X1 U738 ( .A1(n526), .A2(n503), .B1(n377), .B2(n568), .ZN(n256) );
  OAI22_X1 U739 ( .A1(n526), .A2(n373), .B1(n372), .B2(n568), .ZN(n296) );
  OAI22_X1 U740 ( .A1(n18), .A2(n374), .B1(n373), .B2(n568), .ZN(n297) );
  OAI22_X1 U741 ( .A1(n527), .A2(n376), .B1(n375), .B2(n568), .ZN(n299) );
  OAI22_X1 U742 ( .A1(n526), .A2(n368), .B1(n367), .B2(n568), .ZN(n291) );
  OAI22_X1 U743 ( .A1(n526), .A2(n371), .B1(n370), .B2(n568), .ZN(n294) );
  OAI22_X1 U744 ( .A1(n527), .A2(n369), .B1(n368), .B2(n568), .ZN(n292) );
  XNOR2_X1 U745 ( .A(n576), .B(n420), .ZN(n386) );
  OAI22_X1 U746 ( .A1(n18), .A2(n366), .B1(n365), .B2(n568), .ZN(n289) );
  INV_X1 U747 ( .A(n567), .ZN(n245) );
  XNOR2_X1 U748 ( .A(n576), .B(n571), .ZN(n391) );
  XNOR2_X1 U749 ( .A(n576), .B(n423), .ZN(n389) );
  XNOR2_X1 U750 ( .A(n576), .B(n424), .ZN(n390) );
  XNOR2_X1 U751 ( .A(n576), .B(n422), .ZN(n388) );
  XNOR2_X1 U752 ( .A(n576), .B(n421), .ZN(n387) );
  OAI21_X1 U753 ( .B1(n87), .B2(n85), .A(n86), .ZN(n84) );
  XOR2_X1 U754 ( .A(n56), .B(n525), .Z(product[5]) );
  OAI21_X1 U755 ( .B1(n64), .B2(n506), .A(n65), .ZN(n63) );
  OAI21_X1 U756 ( .B1(n556), .B2(n78), .A(n79), .ZN(n77) );
  OAI21_X1 U757 ( .B1(n506), .B2(n71), .A(n72), .ZN(n70) );
  INV_X1 U758 ( .A(n537), .ZN(n87) );
  OAI21_X1 U759 ( .B1(n508), .B2(n89), .A(n90), .ZN(n88) );
  NAND2_X1 U760 ( .A1(n329), .A2(n258), .ZN(n122) );
  OAI22_X1 U761 ( .A1(n554), .A2(n570), .B1(n409), .B2(n573), .ZN(n258) );
  OAI22_X1 U762 ( .A1(n547), .A2(n379), .B1(n378), .B2(n524), .ZN(n301) );
  OAI22_X1 U763 ( .A1(n522), .A2(n380), .B1(n379), .B2(n524), .ZN(n302) );
  OAI22_X1 U764 ( .A1(n522), .A2(n385), .B1(n384), .B2(n524), .ZN(n307) );
  OAI22_X1 U765 ( .A1(n547), .A2(n382), .B1(n381), .B2(n532), .ZN(n304) );
  OAI22_X1 U766 ( .A1(n523), .A2(n381), .B1(n380), .B2(n495), .ZN(n303) );
  NAND2_X1 U767 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U768 ( .A1(n548), .A2(n383), .B1(n532), .B2(n382), .ZN(n305) );
  OAI22_X1 U769 ( .A1(n548), .A2(n384), .B1(n383), .B2(n532), .ZN(n306) );
  OAI22_X1 U770 ( .A1(n522), .A2(n386), .B1(n385), .B2(n532), .ZN(n308) );
  OAI22_X1 U771 ( .A1(n523), .A2(n387), .B1(n386), .B2(n532), .ZN(n309) );
  OAI22_X1 U772 ( .A1(n523), .A2(n515), .B1(n392), .B2(n495), .ZN(n257) );
  OAI22_X1 U773 ( .A1(n12), .A2(n389), .B1(n532), .B2(n388), .ZN(n311) );
  OAI22_X1 U774 ( .A1(n547), .A2(n388), .B1(n387), .B2(n532), .ZN(n310) );
  OAI22_X1 U775 ( .A1(n12), .A2(n390), .B1(n532), .B2(n389), .ZN(n312) );
  INV_X1 U776 ( .A(n532), .ZN(n247) );
  OAI22_X1 U777 ( .A1(n522), .A2(n391), .B1(n390), .B2(n532), .ZN(n313) );
  INV_X1 U778 ( .A(n581), .ZN(n580) );
  INV_X1 U779 ( .A(n31), .ZN(n587) );
  INV_X1 U780 ( .A(n589), .ZN(n588) );
  INV_X1 U781 ( .A(n36), .ZN(n589) );
  INV_X1 U782 ( .A(n591), .ZN(n590) );
  INV_X1 U783 ( .A(n40), .ZN(n591) );
  XOR2_X1 U784 ( .A(n259), .B(n251), .Z(n148) );
  XOR2_X1 U785 ( .A(n289), .B(n279), .Z(n146) );
  XOR2_X1 U786 ( .A(n149), .B(n147), .Z(n144) );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_9_DW01_add_2 ( A, B, CI, 
        SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n8, n9, n10, n11, n12, n13, n14, n15, n16, n19,
         n20, n22, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n44, n45, n47, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n65, n67, n68, n69, n70,
         n71, n73, n75, n76, n77, n78, n79, n81, n83, n84, n86, n88, n90, n91,
         n94, n95, n96, n98, n100, n157, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175;

  AOI21_X1 U122 ( .B1(n52), .B2(n60), .A(n53), .ZN(n157) );
  AND2_X1 U123 ( .A1(n169), .A2(n86), .ZN(SUM[0]) );
  OR2_X1 U124 ( .A1(A[15]), .A2(B[15]), .ZN(n159) );
  XNOR2_X1 U125 ( .A(n45), .B(n160), .ZN(SUM[10]) );
  AND2_X1 U126 ( .A1(n166), .A2(n44), .ZN(n160) );
  NOR2_X1 U127 ( .A1(A[11]), .A2(B[11]), .ZN(n35) );
  OR2_X1 U128 ( .A1(A[13]), .A2(B[13]), .ZN(n161) );
  CLKBUF_X1 U129 ( .A(n29), .Z(n162) );
  NOR2_X1 U130 ( .A1(A[8]), .A2(B[8]), .ZN(n163) );
  NOR2_X1 U131 ( .A1(A[12]), .A2(B[12]), .ZN(n164) );
  NOR2_X1 U132 ( .A1(A[12]), .A2(B[12]), .ZN(n32) );
  NOR2_X1 U133 ( .A1(A[14]), .A2(B[14]), .ZN(n165) );
  NOR2_X1 U134 ( .A1(A[14]), .A2(B[14]), .ZN(n25) );
  OR2_X1 U135 ( .A1(A[10]), .A2(B[10]), .ZN(n166) );
  INV_X1 U136 ( .A(n167), .ZN(n44) );
  AND2_X1 U137 ( .A1(A[10]), .A2(B[10]), .ZN(n167) );
  AOI21_X1 U138 ( .B1(n38), .B2(n30), .A(n31), .ZN(n168) );
  OR2_X1 U139 ( .A1(A[0]), .A2(B[0]), .ZN(n169) );
  INV_X1 U140 ( .A(n157), .ZN(n50) );
  INV_X1 U141 ( .A(n38), .ZN(n37) );
  INV_X1 U142 ( .A(n67), .ZN(n65) );
  AOI21_X1 U143 ( .B1(n171), .B2(n76), .A(n73), .ZN(n71) );
  INV_X1 U144 ( .A(n75), .ZN(n73) );
  OR2_X1 U145 ( .A1(n165), .A2(n28), .ZN(n170) );
  OAI21_X1 U146 ( .B1(n79), .B2(n77), .A(n78), .ZN(n76) );
  AOI21_X1 U147 ( .B1(n50), .B2(n172), .A(n47), .ZN(n45) );
  NAND2_X1 U148 ( .A1(n94), .A2(n55), .ZN(n9) );
  INV_X1 U149 ( .A(n86), .ZN(n84) );
  OAI21_X1 U150 ( .B1(n59), .B2(n57), .A(n58), .ZN(n56) );
  INV_X1 U151 ( .A(n49), .ZN(n47) );
  AOI21_X1 U152 ( .B1(n173), .B2(n84), .A(n81), .ZN(n79) );
  INV_X1 U153 ( .A(n83), .ZN(n81) );
  INV_X1 U154 ( .A(n164), .ZN(n90) );
  NAND2_X1 U155 ( .A1(n172), .A2(n49), .ZN(n8) );
  NAND2_X1 U156 ( .A1(n95), .A2(n58), .ZN(n10) );
  INV_X1 U157 ( .A(n57), .ZN(n95) );
  NAND2_X1 U158 ( .A1(n100), .A2(n78), .ZN(n15) );
  INV_X1 U159 ( .A(n77), .ZN(n100) );
  NAND2_X1 U160 ( .A1(n98), .A2(n70), .ZN(n13) );
  INV_X1 U161 ( .A(n69), .ZN(n98) );
  NAND2_X1 U162 ( .A1(n171), .A2(n75), .ZN(n14) );
  NAND2_X1 U163 ( .A1(n175), .A2(n67), .ZN(n12) );
  NAND2_X1 U164 ( .A1(n173), .A2(n83), .ZN(n16) );
  NAND2_X1 U165 ( .A1(n96), .A2(n62), .ZN(n11) );
  INV_X1 U166 ( .A(n61), .ZN(n96) );
  NAND2_X1 U167 ( .A1(n88), .A2(n26), .ZN(n3) );
  NAND2_X1 U168 ( .A1(n90), .A2(n33), .ZN(n5) );
  XOR2_X1 U169 ( .A(n37), .B(n6), .Z(SUM[11]) );
  NAND2_X1 U170 ( .A1(n91), .A2(n36), .ZN(n6) );
  XOR2_X1 U171 ( .A(n59), .B(n10), .Z(SUM[7]) );
  XNOR2_X1 U172 ( .A(n12), .B(n68), .ZN(SUM[5]) );
  XNOR2_X1 U173 ( .A(n14), .B(n76), .ZN(SUM[3]) );
  XOR2_X1 U174 ( .A(n15), .B(n79), .Z(SUM[2]) );
  NOR2_X1 U175 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  OR2_X1 U176 ( .A1(A[3]), .A2(B[3]), .ZN(n171) );
  NOR2_X1 U177 ( .A1(A[7]), .A2(B[7]), .ZN(n57) );
  NOR2_X1 U178 ( .A1(A[8]), .A2(B[8]), .ZN(n54) );
  OR2_X1 U179 ( .A1(A[9]), .A2(B[9]), .ZN(n172) );
  NOR2_X1 U180 ( .A1(A[2]), .A2(B[2]), .ZN(n77) );
  NAND2_X1 U181 ( .A1(A[11]), .A2(B[11]), .ZN(n36) );
  OR2_X1 U182 ( .A1(A[1]), .A2(B[1]), .ZN(n173) );
  OR2_X1 U183 ( .A1(A[10]), .A2(B[10]), .ZN(n174) );
  NAND2_X1 U184 ( .A1(n159), .A2(n19), .ZN(n2) );
  NAND2_X1 U185 ( .A1(A[14]), .A2(B[14]), .ZN(n26) );
  XNOR2_X1 U186 ( .A(n50), .B(n8), .ZN(SUM[9]) );
  XNOR2_X1 U187 ( .A(n56), .B(n9), .ZN(SUM[8]) );
  NOR2_X1 U188 ( .A1(A[4]), .A2(B[4]), .ZN(n69) );
  NOR2_X1 U189 ( .A1(A[6]), .A2(B[6]), .ZN(n61) );
  NAND2_X1 U190 ( .A1(A[7]), .A2(B[7]), .ZN(n58) );
  NAND2_X1 U191 ( .A1(A[2]), .A2(B[2]), .ZN(n78) );
  NAND2_X1 U192 ( .A1(A[5]), .A2(B[5]), .ZN(n67) );
  NAND2_X1 U193 ( .A1(A[1]), .A2(B[1]), .ZN(n83) );
  NAND2_X1 U194 ( .A1(A[0]), .A2(B[0]), .ZN(n86) );
  NAND2_X1 U195 ( .A1(A[6]), .A2(B[6]), .ZN(n62) );
  NAND2_X1 U196 ( .A1(A[4]), .A2(B[4]), .ZN(n70) );
  NAND2_X1 U197 ( .A1(A[3]), .A2(B[3]), .ZN(n75) );
  OR2_X1 U198 ( .A1(A[5]), .A2(B[5]), .ZN(n175) );
  XOR2_X1 U199 ( .A(n13), .B(n71), .Z(SUM[4]) );
  XNOR2_X1 U200 ( .A(n16), .B(n84), .ZN(SUM[1]) );
  NAND2_X1 U201 ( .A1(n161), .A2(n29), .ZN(n4) );
  NAND2_X1 U202 ( .A1(A[12]), .A2(B[12]), .ZN(n33) );
  INV_X1 U203 ( .A(n24), .ZN(n22) );
  XOR2_X1 U204 ( .A(n168), .B(n4), .Z(SUM[13]) );
  NAND2_X1 U205 ( .A1(A[13]), .A2(B[13]), .ZN(n29) );
  OAI21_X1 U206 ( .B1(n37), .B2(n35), .A(n36), .ZN(n34) );
  INV_X1 U207 ( .A(n35), .ZN(n91) );
  NAND2_X1 U208 ( .A1(A[9]), .A2(B[9]), .ZN(n49) );
  OAI21_X1 U209 ( .B1(n71), .B2(n69), .A(n70), .ZN(n68) );
  INV_X1 U210 ( .A(n163), .ZN(n94) );
  NOR2_X1 U211 ( .A1(n163), .A2(n57), .ZN(n52) );
  OAI21_X1 U212 ( .B1(n54), .B2(n58), .A(n55), .ZN(n53) );
  NAND2_X1 U213 ( .A1(A[8]), .A2(B[8]), .ZN(n55) );
  AOI21_X1 U214 ( .B1(n175), .B2(n68), .A(n65), .ZN(n63) );
  XOR2_X1 U215 ( .A(n11), .B(n63), .Z(SUM[6]) );
  INV_X1 U216 ( .A(n60), .ZN(n59) );
  AOI21_X1 U217 ( .B1(n52), .B2(n60), .A(n53), .ZN(n51) );
  OAI21_X1 U218 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  INV_X1 U219 ( .A(n165), .ZN(n88) );
  OAI21_X1 U220 ( .B1(n29), .B2(n25), .A(n26), .ZN(n24) );
  NAND2_X1 U221 ( .A1(A[15]), .A2(B[15]), .ZN(n19) );
  XNOR2_X1 U222 ( .A(n27), .B(n3), .ZN(SUM[14]) );
  NAND2_X1 U223 ( .A1(n166), .A2(n172), .ZN(n39) );
  AOI21_X1 U224 ( .B1(n174), .B2(n47), .A(n167), .ZN(n40) );
  XNOR2_X1 U225 ( .A(n34), .B(n5), .ZN(SUM[12]) );
  XNOR2_X1 U226 ( .A(n20), .B(n2), .ZN(SUM[15]) );
  OAI21_X1 U227 ( .B1(n168), .B2(n28), .A(n162), .ZN(n27) );
  OAI21_X1 U228 ( .B1(n32), .B2(n36), .A(n33), .ZN(n31) );
  NOR2_X1 U229 ( .A1(n164), .A2(n35), .ZN(n30) );
  OAI21_X1 U230 ( .B1(n168), .B2(n170), .A(n22), .ZN(n20) );
  OAI21_X1 U231 ( .B1(n39), .B2(n51), .A(n40), .ZN(n38) );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_9 ( clk, clear_acc, 
        data_out_x, data_out, data_out_w, data_out_b, wr_en_y, m_valid, 
        m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [4:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
         N39, N40, N41, N42, N43, N44, n1, n2, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n85, n102, n111, n112, n113, n114, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n18), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n221), .CK(clk), .Q(n22) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n222), .CK(clk), .Q(n23) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n223), .CK(clk), .Q(n24) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n224), .CK(clk), .Q(n25) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n225), .CK(clk), .Q(n26) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n226), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n227), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n228), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n229), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n230), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n231), .CK(clk), .Q(n34) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n232), .CK(clk), .Q(n35) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n233), .CK(clk), .Q(n36) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n234), .CK(clk), .Q(n37) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n235), .CK(clk), .Q(n38) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n236), .CK(clk), .Q(n40) );
  DFF_X1 \f_reg[0]  ( .D(n111), .CK(clk), .Q(f[0]), .QN(n210) );
  DFF_X1 \f_reg[1]  ( .D(n102), .CK(clk), .Q(f[1]), .QN(n211) );
  DFF_X1 \f_reg[2]  ( .D(n85), .CK(clk), .Q(f[2]), .QN(n212) );
  DFF_X1 \f_reg[8]  ( .D(n78), .CK(clk), .Q(f[8]), .QN(n214) );
  DFF_X1 \f_reg[9]  ( .D(n77), .CK(clk), .Q(f[9]), .QN(n215) );
  DFF_X1 \f_reg[10]  ( .D(n76), .CK(clk), .Q(n50), .QN(n216) );
  DFF_X1 \f_reg[11]  ( .D(n75), .CK(clk), .Q(n48), .QN(n217) );
  DFF_X1 \f_reg[12]  ( .D(n1), .CK(clk), .Q(n47), .QN(n218) );
  DFF_X1 \f_reg[13]  ( .D(n74), .CK(clk), .Q(n45), .QN(n219) );
  DFF_X1 \f_reg[14]  ( .D(n7), .CK(clk), .Q(n44), .QN(n220) );
  DFF_X1 \f_reg[15]  ( .D(n8), .CK(clk), .Q(f[15]), .QN(n71) );
  DFF_X1 \data_out_reg[15]  ( .D(n113), .CK(clk), .Q(data_out[15]), .QN(n193)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n114), .CK(clk), .Q(data_out[14]), .QN(n192)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n164), .CK(clk), .Q(data_out[13]), .QN(n191)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n165), .CK(clk), .Q(data_out[12]), .QN(n190)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n166), .CK(clk), .Q(data_out[11]), .QN(n189)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n167), .CK(clk), .Q(data_out[10]), .QN(n188)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n168), .CK(clk), .Q(data_out[9]), .QN(n187) );
  DFF_X1 \data_out_reg[8]  ( .D(n169), .CK(clk), .Q(data_out[8]), .QN(n186) );
  DFF_X1 \data_out_reg[7]  ( .D(n170), .CK(clk), .Q(data_out[7]), .QN(n185) );
  DFF_X1 \data_out_reg[6]  ( .D(n171), .CK(clk), .Q(data_out[6]), .QN(n184) );
  DFF_X1 \data_out_reg[5]  ( .D(n172), .CK(clk), .Q(data_out[5]), .QN(n183) );
  DFF_X1 \data_out_reg[4]  ( .D(n173), .CK(clk), .Q(data_out[4]), .QN(n182) );
  DFF_X1 \data_out_reg[3]  ( .D(n174), .CK(clk), .Q(data_out[3]), .QN(n181) );
  DFF_X1 \data_out_reg[2]  ( .D(n175), .CK(clk), .Q(data_out[2]), .QN(n180) );
  DFF_X1 \data_out_reg[1]  ( .D(n176), .CK(clk), .Q(data_out[1]), .QN(n179) );
  DFF_X1 \data_out_reg[0]  ( .D(n177), .CK(clk), .Q(data_out[0]), .QN(n178) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_9_DW_mult_tc_1 mult_2021 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_9_DW01_add_2 add_2022 ( .A({n200, 
        n199, n198, n197, n196, n195, n209, n208, n207, n206, n205, n204, n203, 
        n202, n201, n194}), .B({f[15], n44, n45, n47, n48, n50, f[9:0]}), .CI(
        1'b0), .SUM(adder) );
  DFF_X1 \f_reg[3]  ( .D(n83), .CK(clk), .Q(f[3]), .QN(n63) );
  DFF_X1 \f_reg[4]  ( .D(n82), .CK(clk), .Q(f[4]), .QN(n64) );
  DFF_X1 \f_reg[5]  ( .D(n81), .CK(clk), .Q(f[5]), .QN(n65) );
  DFF_X1 \f_reg[6]  ( .D(n80), .CK(clk), .Q(f[6]), .QN(n66) );
  DFF_X1 \f_reg[7]  ( .D(n79), .CK(clk), .Q(f[7]), .QN(n213) );
  DFF_X2 delay_reg ( .D(n112), .CK(clk), .Q(n2), .QN(n237) );
  AND2_X1 U3 ( .A1(n43), .A2(n19), .ZN(n15) );
  NAND3_X1 U4 ( .A1(n5), .A2(n4), .A3(n6), .ZN(n1) );
  MUX2_X2 U5 ( .A(N39), .B(n27), .S(n2), .Z(n195) );
  NAND2_X1 U6 ( .A1(data_out_b[12]), .A2(n17), .ZN(n4) );
  NAND2_X1 U8 ( .A1(adder[12]), .A2(n15), .ZN(n5) );
  NAND2_X1 U9 ( .A1(n61), .A2(n47), .ZN(n6) );
  INV_X1 U10 ( .A(n43), .ZN(n61) );
  NAND3_X1 U11 ( .A1(n13), .A2(n12), .A3(n14), .ZN(n7) );
  NAND3_X1 U12 ( .A1(n10), .A2(n9), .A3(n11), .ZN(n8) );
  MUX2_X2 U13 ( .A(n24), .B(N42), .S(n237), .Z(n198) );
  MUX2_X2 U14 ( .A(n26), .B(N40), .S(n237), .Z(n196) );
  MUX2_X2 U15 ( .A(n29), .B(N37), .S(n237), .Z(n208) );
  NAND2_X1 U16 ( .A1(data_out_b[15]), .A2(n17), .ZN(n9) );
  NAND2_X1 U17 ( .A1(adder[15]), .A2(n15), .ZN(n10) );
  NAND2_X1 U18 ( .A1(n61), .A2(f[15]), .ZN(n11) );
  MUX2_X2 U19 ( .A(n23), .B(N43), .S(n237), .Z(n199) );
  MUX2_X2 U20 ( .A(n25), .B(N41), .S(n237), .Z(n197) );
  NAND2_X1 U21 ( .A1(data_out_b[14]), .A2(n17), .ZN(n12) );
  NAND2_X1 U22 ( .A1(adder[14]), .A2(n15), .ZN(n13) );
  NAND2_X1 U23 ( .A1(n61), .A2(n44), .ZN(n14) );
  INV_X1 U24 ( .A(n19), .ZN(n17) );
  NAND2_X1 U25 ( .A1(n112), .A2(n16), .ZN(n239) );
  INV_X1 U26 ( .A(clear_acc), .ZN(n19) );
  OAI22_X1 U27 ( .A1(n181), .A2(n239), .B1(n63), .B2(n238), .ZN(n174) );
  OAI22_X1 U28 ( .A1(n182), .A2(n239), .B1(n64), .B2(n238), .ZN(n173) );
  OAI22_X1 U29 ( .A1(n183), .A2(n239), .B1(n65), .B2(n238), .ZN(n172) );
  OAI22_X1 U30 ( .A1(n184), .A2(n239), .B1(n66), .B2(n238), .ZN(n171) );
  OAI22_X1 U31 ( .A1(n185), .A2(n239), .B1(n213), .B2(n238), .ZN(n170) );
  OAI22_X1 U32 ( .A1(n186), .A2(n239), .B1(n214), .B2(n238), .ZN(n169) );
  OAI22_X1 U33 ( .A1(n187), .A2(n239), .B1(n215), .B2(n238), .ZN(n168) );
  MUX2_X1 U34 ( .A(n36), .B(N32), .S(n237), .Z(n203) );
  INV_X1 U35 ( .A(n21), .ZN(n39) );
  INV_X1 U36 ( .A(wr_en_y), .ZN(n16) );
  INV_X1 U37 ( .A(n19), .ZN(n18) );
  INV_X1 U38 ( .A(m_ready), .ZN(n20) );
  NAND2_X1 U39 ( .A1(m_valid), .A2(n20), .ZN(n41) );
  OAI21_X1 U40 ( .B1(sel[4]), .B2(n73), .A(n41), .ZN(n112) );
  NAND2_X1 U41 ( .A1(clear_acc_delay), .A2(n237), .ZN(n21) );
  MUX2_X1 U42 ( .A(n22), .B(N44), .S(n39), .Z(n221) );
  MUX2_X1 U43 ( .A(n22), .B(N44), .S(n237), .Z(n200) );
  MUX2_X1 U44 ( .A(n23), .B(N43), .S(n39), .Z(n222) );
  MUX2_X1 U45 ( .A(n24), .B(N42), .S(n39), .Z(n223) );
  MUX2_X1 U46 ( .A(n25), .B(N41), .S(n39), .Z(n224) );
  MUX2_X1 U47 ( .A(n26), .B(N40), .S(n39), .Z(n225) );
  MUX2_X1 U48 ( .A(n27), .B(N39), .S(n39), .Z(n226) );
  MUX2_X1 U49 ( .A(n28), .B(N38), .S(n39), .Z(n227) );
  MUX2_X1 U50 ( .A(n28), .B(N38), .S(n237), .Z(n209) );
  MUX2_X1 U51 ( .A(n29), .B(N37), .S(n39), .Z(n228) );
  MUX2_X1 U52 ( .A(n32), .B(N36), .S(n39), .Z(n229) );
  MUX2_X1 U53 ( .A(n32), .B(N36), .S(n237), .Z(n207) );
  MUX2_X1 U54 ( .A(n33), .B(N35), .S(n39), .Z(n230) );
  MUX2_X1 U55 ( .A(n33), .B(N35), .S(n237), .Z(n206) );
  MUX2_X1 U56 ( .A(n34), .B(N34), .S(n39), .Z(n231) );
  MUX2_X1 U57 ( .A(n34), .B(N34), .S(n237), .Z(n205) );
  MUX2_X1 U58 ( .A(n35), .B(N33), .S(n39), .Z(n232) );
  MUX2_X1 U59 ( .A(n35), .B(N33), .S(n237), .Z(n204) );
  MUX2_X1 U60 ( .A(n36), .B(N32), .S(n39), .Z(n233) );
  MUX2_X1 U61 ( .A(n37), .B(N31), .S(n39), .Z(n234) );
  MUX2_X1 U62 ( .A(n37), .B(N31), .S(n237), .Z(n202) );
  MUX2_X1 U63 ( .A(n38), .B(N30), .S(n39), .Z(n235) );
  MUX2_X1 U64 ( .A(n38), .B(N30), .S(n237), .Z(n201) );
  MUX2_X1 U65 ( .A(n40), .B(N29), .S(n39), .Z(n236) );
  MUX2_X1 U66 ( .A(n40), .B(N29), .S(n237), .Z(n194) );
  INV_X1 U67 ( .A(n41), .ZN(n42) );
  OAI21_X1 U68 ( .B1(n42), .B2(n2), .A(n19), .ZN(n43) );
  AOI222_X1 U69 ( .A1(data_out_b[13]), .A2(n17), .B1(adder[13]), .B2(n15), 
        .C1(n61), .C2(n45), .ZN(n46) );
  INV_X1 U70 ( .A(n46), .ZN(n74) );
  AOI222_X1 U71 ( .A1(data_out_b[11]), .A2(n17), .B1(adder[11]), .B2(n15), 
        .C1(n61), .C2(n48), .ZN(n49) );
  INV_X1 U72 ( .A(n49), .ZN(n75) );
  AOI222_X1 U73 ( .A1(data_out_b[10]), .A2(n17), .B1(adder[10]), .B2(n15), 
        .C1(n61), .C2(n50), .ZN(n51) );
  INV_X1 U74 ( .A(n51), .ZN(n76) );
  AOI222_X1 U75 ( .A1(data_out_b[8]), .A2(n17), .B1(adder[8]), .B2(n15), .C1(
        n61), .C2(f[8]), .ZN(n52) );
  INV_X1 U76 ( .A(n52), .ZN(n78) );
  AOI222_X1 U77 ( .A1(data_out_b[7]), .A2(n17), .B1(adder[7]), .B2(n15), .C1(
        n61), .C2(f[7]), .ZN(n53) );
  INV_X1 U78 ( .A(n53), .ZN(n79) );
  AOI222_X1 U79 ( .A1(data_out_b[6]), .A2(n17), .B1(adder[6]), .B2(n15), .C1(
        n61), .C2(f[6]), .ZN(n54) );
  INV_X1 U80 ( .A(n54), .ZN(n80) );
  AOI222_X1 U81 ( .A1(data_out_b[5]), .A2(n17), .B1(adder[5]), .B2(n15), .C1(
        n61), .C2(f[5]), .ZN(n55) );
  INV_X1 U82 ( .A(n55), .ZN(n81) );
  AOI222_X1 U83 ( .A1(data_out_b[4]), .A2(n17), .B1(adder[4]), .B2(n15), .C1(
        n61), .C2(f[4]), .ZN(n56) );
  INV_X1 U84 ( .A(n56), .ZN(n82) );
  AOI222_X1 U85 ( .A1(data_out_b[3]), .A2(n17), .B1(adder[3]), .B2(n15), .C1(
        n61), .C2(f[3]), .ZN(n57) );
  INV_X1 U86 ( .A(n57), .ZN(n83) );
  AOI222_X1 U87 ( .A1(data_out_b[2]), .A2(n18), .B1(adder[2]), .B2(n15), .C1(
        n61), .C2(f[2]), .ZN(n58) );
  INV_X1 U88 ( .A(n58), .ZN(n85) );
  AOI222_X1 U89 ( .A1(data_out_b[1]), .A2(n18), .B1(adder[1]), .B2(n15), .C1(
        n61), .C2(f[1]), .ZN(n59) );
  INV_X1 U90 ( .A(n59), .ZN(n102) );
  AOI222_X1 U91 ( .A1(data_out_b[0]), .A2(n18), .B1(adder[0]), .B2(n15), .C1(
        n61), .C2(f[0]), .ZN(n60) );
  INV_X1 U92 ( .A(n60), .ZN(n111) );
  AOI222_X1 U93 ( .A1(data_out_b[9]), .A2(n18), .B1(adder[9]), .B2(n15), .C1(
        n61), .C2(f[9]), .ZN(n62) );
  INV_X1 U94 ( .A(n62), .ZN(n77) );
  NOR4_X1 U95 ( .A1(n48), .A2(n47), .A3(n45), .A4(n44), .ZN(n70) );
  NOR4_X1 U96 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n50), .ZN(n69) );
  NAND4_X1 U97 ( .A1(n66), .A2(n65), .A3(n64), .A4(n63), .ZN(n67) );
  NOR4_X1 U98 ( .A1(n67), .A2(f[0]), .A3(f[1]), .A4(f[2]), .ZN(n68) );
  NAND3_X1 U99 ( .A1(n70), .A2(n69), .A3(n68), .ZN(n72) );
  NAND3_X1 U100 ( .A1(wr_en_y), .A2(n72), .A3(n71), .ZN(n238) );
  OAI22_X1 U101 ( .A1(n178), .A2(n239), .B1(n210), .B2(n238), .ZN(n177) );
  OAI22_X1 U102 ( .A1(n179), .A2(n239), .B1(n211), .B2(n238), .ZN(n176) );
  OAI22_X1 U103 ( .A1(n180), .A2(n239), .B1(n212), .B2(n238), .ZN(n175) );
  OAI22_X1 U104 ( .A1(n188), .A2(n239), .B1(n216), .B2(n238), .ZN(n167) );
  OAI22_X1 U105 ( .A1(n189), .A2(n239), .B1(n217), .B2(n238), .ZN(n166) );
  OAI22_X1 U106 ( .A1(n190), .A2(n239), .B1(n218), .B2(n238), .ZN(n165) );
  OAI22_X1 U107 ( .A1(n191), .A2(n239), .B1(n219), .B2(n238), .ZN(n164) );
  OAI22_X1 U108 ( .A1(n192), .A2(n239), .B1(n220), .B2(n238), .ZN(n114) );
  OAI22_X1 U109 ( .A1(n193), .A2(n239), .B1(n71), .B2(n238), .ZN(n113) );
  AND4_X1 U110 ( .A1(sel[3]), .A2(sel[2]), .A3(sel[1]), .A4(sel[0]), .ZN(n73)
         );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_8_DW_mult_tc_1 ( a, b, 
        product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n9, n12, n13, n16, n18, n19, n21, n23, n25, n27, n29, n31,
         n32, n34, n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n50,
         n52, n53, n54, n55, n56, n57, n58, n59, n62, n63, n64, n65, n67, n69,
         n70, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n93, n95, n96, n97, n98, n99, n101,
         n103, n104, n105, n106, n107, n111, n112, n113, n114, n115, n117,
         n119, n120, n122, n127, n129, n131, n135, n139, n141, n142, n143,
         n144, n145, n146, n148, n149, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n237, n245, n247, n249, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n418, n419, n420, n421, n422, n423, n424, n426, n427, n433, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U148 ( .A(n265), .B(n144), .Z(n145) );
  XOR2_X1 U152 ( .A(n301), .B(n148), .Z(n149) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U162 ( .A(n170), .B(n172), .CI(n179), .CO(n165), .S(n166) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n263), .CI(n291), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n252), .B(n317), .CO(n173), .S(n174) );
  FA_X1 U167 ( .A(n180), .B(n187), .CI(n178), .CO(n175), .S(n176) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U169 ( .A(n193), .B(n282), .CI(n191), .CO(n179), .S(n180) );
  FA_X1 U170 ( .A(n268), .B(n292), .CI(n274), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U172 ( .A(n197), .B(n190), .CI(n188), .CO(n185), .S(n186) );
  FA_X1 U173 ( .A(n199), .B(n201), .CI(n192), .CO(n187), .S(n188) );
  FA_X1 U174 ( .A(n275), .B(n293), .CI(n194), .CO(n189), .S(n190) );
  FA_X1 U175 ( .A(n305), .B(n253), .CI(n283), .CO(n191), .S(n192) );
  HA_X1 U176 ( .A(n319), .B(n269), .CO(n193), .S(n194) );
  FA_X1 U177 ( .A(n205), .B(n200), .CI(n198), .CO(n195), .S(n196) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U179 ( .A(n276), .B(n294), .CI(n284), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n320), .B(n270), .CI(n306), .CO(n201), .S(n202) );
  FA_X1 U181 ( .A(n208), .B(n213), .CI(n206), .CO(n203), .S(n204) );
  FA_X1 U182 ( .A(n210), .B(n307), .CI(n215), .CO(n205), .S(n206) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n322), .B(n278), .CI(n308), .CO(n215), .S(n216) );
  FA_X1 U188 ( .A(n225), .B(n222), .CI(n220), .CO(n217), .S(n218) );
  FA_X1 U189 ( .A(n309), .B(n297), .CI(n255), .CO(n219), .S(n220) );
  HA_X1 U190 ( .A(n287), .B(n323), .CO(n221), .S(n222) );
  FA_X1 U192 ( .A(n324), .B(n288), .CI(n310), .CO(n225), .S(n226) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  HA_X1 U194 ( .A(n311), .B(n325), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n326), .B(n300), .CI(n312), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  XOR2_X1 U414 ( .A(n594), .B(a[10]), .Z(n522) );
  BUF_X1 U415 ( .A(n514), .Z(n490) );
  CLKBUF_X1 U416 ( .A(n19), .Z(n514) );
  CLKBUF_X1 U417 ( .A(n19), .Z(n513) );
  AND2_X1 U418 ( .A1(n232), .A2(n233), .ZN(n549) );
  BUF_X1 U419 ( .A(n37), .Z(n519) );
  BUF_X1 U420 ( .A(n12), .Z(n555) );
  BUF_X2 U421 ( .A(n16), .Z(n575) );
  INV_X1 U422 ( .A(n549), .ZN(n111) );
  OR2_X1 U423 ( .A1(n164), .A2(n175), .ZN(n491) );
  OR2_X1 U424 ( .A1(n329), .A2(n258), .ZN(n492) );
  BUF_X1 U425 ( .A(n91), .Z(n552) );
  XOR2_X1 U426 ( .A(n589), .B(a[6]), .Z(n493) );
  NAND2_X1 U427 ( .A1(n196), .A2(n203), .ZN(n494) );
  INV_X1 U428 ( .A(n502), .ZN(n495) );
  XNOR2_X1 U429 ( .A(n513), .B(a[6]), .ZN(n496) );
  BUF_X1 U430 ( .A(n12), .Z(n554) );
  INV_X1 U431 ( .A(n596), .ZN(n497) );
  OR2_X1 U432 ( .A1(n75), .A2(n78), .ZN(n498) );
  CLKBUF_X1 U433 ( .A(n228), .Z(n499) );
  XOR2_X1 U434 ( .A(n586), .B(a[4]), .Z(n500) );
  OR2_X2 U435 ( .A1(n496), .A2(n563), .ZN(n542) );
  INV_X1 U436 ( .A(n593), .ZN(n501) );
  XOR2_X1 U437 ( .A(n596), .B(a[14]), .Z(n41) );
  INV_X1 U438 ( .A(n596), .ZN(n595) );
  OR2_X1 U439 ( .A1(n196), .A2(n203), .ZN(n502) );
  NOR2_X1 U440 ( .A1(n196), .A2(n203), .ZN(n85) );
  OAI21_X1 U441 ( .B1(n91), .B2(n89), .A(n90), .ZN(n503) );
  OAI21_X1 U442 ( .B1(n91), .B2(n89), .A(n90), .ZN(n88) );
  INV_X1 U443 ( .A(n507), .ZN(n504) );
  INV_X1 U444 ( .A(n587), .ZN(n505) );
  NAND2_X2 U445 ( .A1(n564), .A2(n500), .ZN(n18) );
  BUF_X2 U446 ( .A(n9), .Z(n550) );
  XNOR2_X1 U447 ( .A(n149), .B(n506), .ZN(n144) );
  XNOR2_X1 U448 ( .A(n146), .B(n271), .ZN(n506) );
  XNOR2_X1 U449 ( .A(n590), .B(a[8]), .ZN(n507) );
  BUF_X1 U450 ( .A(n9), .Z(n576) );
  INV_X1 U451 ( .A(n7), .ZN(n508) );
  INV_X1 U452 ( .A(n594), .ZN(n509) );
  INV_X1 U453 ( .A(n592), .ZN(n510) );
  INV_X1 U454 ( .A(n594), .ZN(n511) );
  INV_X1 U455 ( .A(n594), .ZN(n593) );
  CLKBUF_X1 U456 ( .A(n562), .Z(n517) );
  XOR2_X1 U457 ( .A(n583), .B(a[2]), .Z(n512) );
  XNOR2_X1 U458 ( .A(n166), .B(n515), .ZN(n164) );
  XNOR2_X1 U459 ( .A(n177), .B(n168), .ZN(n515) );
  CLKBUF_X1 U460 ( .A(n107), .Z(n516) );
  XNOR2_X1 U461 ( .A(n503), .B(n518), .ZN(product[10]) );
  NAND2_X1 U462 ( .A1(n502), .A2(n494), .ZN(n518) );
  INV_X1 U463 ( .A(n582), .ZN(n520) );
  INV_X1 U464 ( .A(n592), .ZN(n521) );
  INV_X1 U465 ( .A(n592), .ZN(n591) );
  OR2_X2 U466 ( .A1(n522), .A2(n551), .ZN(n34) );
  XOR2_X1 U467 ( .A(n216), .B(n219), .Z(n523) );
  XOR2_X1 U468 ( .A(n214), .B(n523), .Z(n212) );
  NAND2_X1 U469 ( .A1(n214), .A2(n216), .ZN(n524) );
  NAND2_X1 U470 ( .A1(n214), .A2(n219), .ZN(n525) );
  NAND2_X1 U471 ( .A1(n216), .A2(n219), .ZN(n526) );
  NAND3_X1 U472 ( .A1(n524), .A2(n525), .A3(n526), .ZN(n211) );
  XNOR2_X1 U473 ( .A(n45), .B(n527), .ZN(product[12]) );
  AND2_X1 U474 ( .A1(n536), .A2(n79), .ZN(n527) );
  XOR2_X1 U475 ( .A(n285), .B(n295), .Z(n528) );
  XOR2_X1 U476 ( .A(n254), .B(n528), .Z(n208) );
  NAND2_X1 U477 ( .A1(n254), .A2(n285), .ZN(n529) );
  NAND2_X1 U478 ( .A1(n254), .A2(n295), .ZN(n530) );
  NAND2_X1 U479 ( .A1(n285), .A2(n295), .ZN(n531) );
  NAND3_X1 U480 ( .A1(n529), .A2(n530), .A3(n531), .ZN(n207) );
  OR2_X1 U481 ( .A1(n29), .A2(n592), .ZN(n532) );
  OR2_X1 U482 ( .A1(n353), .A2(n27), .ZN(n533) );
  NAND2_X1 U483 ( .A1(n532), .A2(n533), .ZN(n254) );
  CLKBUF_X1 U484 ( .A(n104), .Z(n534) );
  BUF_X2 U485 ( .A(n580), .Z(n535) );
  INV_X1 U486 ( .A(n249), .ZN(n580) );
  XNOR2_X1 U487 ( .A(n589), .B(a[4]), .ZN(n564) );
  OR2_X1 U488 ( .A1(n176), .A2(n185), .ZN(n536) );
  OR2_X2 U489 ( .A1(n537), .A2(n548), .ZN(n29) );
  XNOR2_X1 U490 ( .A(n591), .B(a[8]), .ZN(n537) );
  NAND2_X1 U491 ( .A1(n166), .A2(n177), .ZN(n538) );
  NAND2_X1 U492 ( .A1(n166), .A2(n168), .ZN(n539) );
  NAND2_X1 U493 ( .A1(n177), .A2(n168), .ZN(n540) );
  NAND3_X1 U494 ( .A1(n538), .A2(n539), .A3(n540), .ZN(n163) );
  OR2_X1 U495 ( .A1(n496), .A2(n563), .ZN(n541) );
  OR2_X1 U496 ( .A1(n547), .A2(n563), .ZN(n23) );
  XNOR2_X1 U497 ( .A(n508), .B(a[2]), .ZN(n565) );
  INV_X2 U498 ( .A(n589), .ZN(n587) );
  CLKBUF_X1 U499 ( .A(n99), .Z(n543) );
  XNOR2_X1 U500 ( .A(n226), .B(n544), .ZN(n224) );
  XNOR2_X1 U501 ( .A(n229), .B(n298), .ZN(n544) );
  NOR2_X1 U502 ( .A1(n164), .A2(n175), .ZN(n75) );
  INV_X1 U503 ( .A(n507), .ZN(n27) );
  NOR2_X1 U504 ( .A1(n186), .A2(n195), .ZN(n545) );
  NOR2_X1 U505 ( .A1(n186), .A2(n195), .ZN(n82) );
  CLKBUF_X1 U506 ( .A(n96), .Z(n546) );
  OAI21_X1 U507 ( .B1(n99), .B2(n97), .A(n98), .ZN(n96) );
  XNOR2_X1 U508 ( .A(n513), .B(a[6]), .ZN(n547) );
  INV_X1 U509 ( .A(n563), .ZN(n21) );
  XOR2_X1 U510 ( .A(a[2]), .B(n583), .Z(n9) );
  XNOR2_X1 U511 ( .A(n590), .B(a[8]), .ZN(n548) );
  INV_X1 U512 ( .A(n551), .ZN(n32) );
  XOR2_X1 U513 ( .A(n586), .B(a[4]), .Z(n16) );
  INV_X1 U514 ( .A(n508), .ZN(n584) );
  XNOR2_X1 U515 ( .A(n592), .B(a[10]), .ZN(n551) );
  XNOR2_X1 U516 ( .A(n583), .B(n249), .ZN(n433) );
  OR2_X1 U517 ( .A1(n499), .A2(n231), .ZN(n553) );
  BUF_X2 U518 ( .A(n12), .Z(n556) );
  NAND2_X1 U519 ( .A1(n512), .A2(n565), .ZN(n12) );
  NAND2_X1 U520 ( .A1(n226), .A2(n229), .ZN(n557) );
  NAND2_X1 U521 ( .A1(n226), .A2(n298), .ZN(n558) );
  NAND2_X1 U522 ( .A1(n229), .A2(n298), .ZN(n559) );
  NAND3_X1 U523 ( .A1(n557), .A2(n558), .A3(n559), .ZN(n223) );
  NAND2_X1 U524 ( .A1(n433), .A2(n580), .ZN(n560) );
  NAND2_X1 U525 ( .A1(n433), .A2(n580), .ZN(n561) );
  AOI21_X1 U526 ( .B1(n80), .B2(n88), .A(n81), .ZN(n562) );
  XNOR2_X1 U527 ( .A(n589), .B(a[6]), .ZN(n563) );
  INV_X2 U528 ( .A(n583), .ZN(n581) );
  BUF_X1 U529 ( .A(n43), .Z(n578) );
  AOI21_X1 U530 ( .B1(n74), .B2(n566), .A(n67), .ZN(n65) );
  INV_X1 U531 ( .A(n69), .ZN(n67) );
  NAND2_X1 U532 ( .A1(n566), .A2(n69), .ZN(n47) );
  NAND2_X1 U533 ( .A1(n73), .A2(n566), .ZN(n64) );
  INV_X1 U534 ( .A(n74), .ZN(n72) );
  INV_X1 U535 ( .A(n95), .ZN(n93) );
  NAND2_X1 U536 ( .A1(n129), .A2(n90), .ZN(n52) );
  INV_X1 U537 ( .A(n89), .ZN(n129) );
  OR2_X1 U538 ( .A1(n152), .A2(n163), .ZN(n566) );
  NAND2_X1 U539 ( .A1(n567), .A2(n95), .ZN(n53) );
  NAND2_X1 U540 ( .A1(n491), .A2(n76), .ZN(n48) );
  OAI21_X1 U541 ( .B1(n75), .B2(n79), .A(n76), .ZN(n74) );
  NOR2_X1 U542 ( .A1(n75), .A2(n78), .ZN(n73) );
  XNOR2_X1 U543 ( .A(n84), .B(n50), .ZN(product[11]) );
  NAND2_X1 U544 ( .A1(n127), .A2(n83), .ZN(n50) );
  NAND2_X1 U545 ( .A1(n152), .A2(n163), .ZN(n69) );
  NAND2_X1 U546 ( .A1(n135), .A2(n114), .ZN(n58) );
  OAI21_X1 U547 ( .B1(n113), .B2(n115), .A(n114), .ZN(n112) );
  NAND2_X1 U548 ( .A1(n553), .A2(n106), .ZN(n56) );
  NAND2_X1 U549 ( .A1(n131), .A2(n98), .ZN(n54) );
  INV_X1 U550 ( .A(n97), .ZN(n131) );
  AOI21_X1 U551 ( .B1(n569), .B2(n112), .A(n549), .ZN(n107) );
  NOR2_X1 U552 ( .A1(n176), .A2(n185), .ZN(n78) );
  NAND2_X1 U553 ( .A1(n569), .A2(n111), .ZN(n57) );
  AOI21_X1 U554 ( .B1(n568), .B2(n120), .A(n117), .ZN(n115) );
  INV_X1 U555 ( .A(n119), .ZN(n117) );
  INV_X1 U556 ( .A(n122), .ZN(n120) );
  XNOR2_X1 U557 ( .A(n59), .B(n120), .ZN(product[2]) );
  NAND2_X1 U558 ( .A1(n568), .A2(n119), .ZN(n59) );
  NAND2_X1 U559 ( .A1(n176), .A2(n185), .ZN(n79) );
  NAND2_X1 U560 ( .A1(n164), .A2(n175), .ZN(n76) );
  NAND2_X1 U561 ( .A1(n212), .A2(n217), .ZN(n95) );
  OR2_X1 U562 ( .A1(n212), .A2(n217), .ZN(n567) );
  NAND2_X1 U563 ( .A1(n204), .A2(n211), .ZN(n90) );
  NAND2_X1 U564 ( .A1(n186), .A2(n195), .ZN(n83) );
  NAND2_X1 U565 ( .A1(n196), .A2(n203), .ZN(n86) );
  XNOR2_X1 U566 ( .A(n63), .B(n46), .ZN(product[15]) );
  NAND2_X1 U567 ( .A1(n570), .A2(n62), .ZN(n46) );
  OR2_X1 U568 ( .A1(n328), .A2(n314), .ZN(n568) );
  NOR2_X1 U569 ( .A1(n218), .A2(n223), .ZN(n97) );
  OR2_X1 U570 ( .A1(n232), .A2(n233), .ZN(n569) );
  NAND2_X1 U571 ( .A1(n218), .A2(n223), .ZN(n98) );
  INV_X1 U572 ( .A(n37), .ZN(n237) );
  NAND2_X1 U573 ( .A1(n228), .A2(n231), .ZN(n106) );
  INV_X1 U574 ( .A(n41), .ZN(n235) );
  OR2_X1 U575 ( .A1(n151), .A2(n139), .ZN(n570) );
  AND2_X1 U576 ( .A1(n492), .A2(n122), .ZN(product[1]) );
  OR2_X1 U577 ( .A1(n224), .A2(n227), .ZN(n577) );
  XNOR2_X1 U578 ( .A(n509), .B(a[12]), .ZN(n37) );
  OR2_X1 U579 ( .A1(n578), .A2(n508), .ZN(n392) );
  AND2_X1 U580 ( .A1(n579), .A2(n563), .ZN(n288) );
  AND2_X1 U581 ( .A1(n579), .A2(n551), .ZN(n270) );
  XNOR2_X1 U582 ( .A(n510), .B(n578), .ZN(n352) );
  XNOR2_X1 U583 ( .A(n155), .B(n572), .ZN(n139) );
  XNOR2_X1 U584 ( .A(n153), .B(n141), .ZN(n572) );
  XNOR2_X1 U585 ( .A(n157), .B(n573), .ZN(n141) );
  XNOR2_X1 U586 ( .A(n145), .B(n143), .ZN(n573) );
  OAI22_X1 U587 ( .A1(n39), .A2(n596), .B1(n337), .B2(n519), .ZN(n252) );
  OR2_X1 U588 ( .A1(n578), .A2(n596), .ZN(n337) );
  OAI22_X1 U589 ( .A1(n42), .A2(n598), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U590 ( .A1(n578), .A2(n598), .ZN(n332) );
  XNOR2_X1 U591 ( .A(n593), .B(n578), .ZN(n343) );
  NAND2_X1 U592 ( .A1(n433), .A2(n580), .ZN(n6) );
  XNOR2_X1 U593 ( .A(n159), .B(n574), .ZN(n142) );
  XNOR2_X1 U594 ( .A(n315), .B(n261), .ZN(n574) );
  XNOR2_X1 U595 ( .A(n588), .B(n578), .ZN(n376) );
  XNOR2_X1 U596 ( .A(n595), .B(n578), .ZN(n336) );
  NAND2_X1 U597 ( .A1(n427), .A2(n37), .ZN(n39) );
  XOR2_X1 U598 ( .A(n595), .B(a[12]), .Z(n427) );
  OAI22_X1 U599 ( .A1(n39), .A2(n336), .B1(n519), .B2(n335), .ZN(n263) );
  AND2_X1 U600 ( .A1(n579), .A2(n237), .ZN(n264) );
  AND2_X1 U601 ( .A1(n579), .A2(n245), .ZN(n300) );
  AND2_X1 U602 ( .A1(n579), .A2(n235), .ZN(n260) );
  OAI22_X1 U603 ( .A1(n39), .A2(n335), .B1(n519), .B2(n334), .ZN(n262) );
  INV_X1 U604 ( .A(n19), .ZN(n590) );
  INV_X1 U605 ( .A(n25), .ZN(n592) );
  AND2_X1 U606 ( .A1(n579), .A2(n507), .ZN(n278) );
  INV_X1 U607 ( .A(n1), .ZN(n583) );
  NAND2_X1 U608 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U609 ( .A(n597), .B(a[14]), .Z(n426) );
  INV_X1 U610 ( .A(n7), .ZN(n586) );
  XNOR2_X1 U611 ( .A(n490), .B(n578), .ZN(n363) );
  AND2_X1 U612 ( .A1(n579), .A2(n247), .ZN(n314) );
  AND2_X1 U613 ( .A1(n579), .A2(n249), .ZN(product[0]) );
  OR2_X1 U614 ( .A1(n578), .A2(n501), .ZN(n344) );
  OR2_X1 U615 ( .A1(n578), .A2(n590), .ZN(n364) );
  OR2_X1 U616 ( .A1(n578), .A2(n592), .ZN(n353) );
  OR2_X1 U617 ( .A1(n578), .A2(n505), .ZN(n377) );
  XNOR2_X1 U618 ( .A(n514), .B(b[9]), .ZN(n354) );
  OAI22_X1 U619 ( .A1(n39), .A2(n334), .B1(n519), .B2(n333), .ZN(n261) );
  XNOR2_X1 U620 ( .A(n595), .B(n422), .ZN(n333) );
  XNOR2_X1 U621 ( .A(n588), .B(b[11]), .ZN(n365) );
  XNOR2_X1 U622 ( .A(n497), .B(n424), .ZN(n335) );
  XNOR2_X1 U623 ( .A(n497), .B(n423), .ZN(n334) );
  OAI22_X1 U624 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U625 ( .A(n597), .B(n424), .ZN(n330) );
  XNOR2_X1 U626 ( .A(n597), .B(n578), .ZN(n331) );
  XNOR2_X1 U627 ( .A(n521), .B(n418), .ZN(n345) );
  XNOR2_X1 U628 ( .A(n593), .B(n420), .ZN(n338) );
  XNOR2_X1 U629 ( .A(n585), .B(b[13]), .ZN(n378) );
  XNOR2_X1 U630 ( .A(n511), .B(n424), .ZN(n342) );
  XNOR2_X1 U631 ( .A(n490), .B(n424), .ZN(n362) );
  XNOR2_X1 U632 ( .A(n591), .B(n424), .ZN(n351) );
  XNOR2_X1 U633 ( .A(n511), .B(n423), .ZN(n341) );
  XNOR2_X1 U634 ( .A(n511), .B(n422), .ZN(n340) );
  XNOR2_X1 U635 ( .A(n593), .B(n421), .ZN(n339) );
  XNOR2_X1 U636 ( .A(n585), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U637 ( .A(n585), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U638 ( .A(n585), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U639 ( .A(n585), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U640 ( .A(n585), .B(n419), .ZN(n385) );
  XNOR2_X1 U641 ( .A(n585), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U642 ( .A(n585), .B(n418), .ZN(n384) );
  XNOR2_X1 U643 ( .A(n514), .B(n423), .ZN(n361) );
  XNOR2_X1 U644 ( .A(n510), .B(n423), .ZN(n350) );
  XNOR2_X1 U645 ( .A(n521), .B(n422), .ZN(n349) );
  XNOR2_X1 U646 ( .A(n514), .B(n422), .ZN(n360) );
  XNOR2_X1 U647 ( .A(n588), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U648 ( .A(n588), .B(n418), .ZN(n369) );
  XNOR2_X1 U649 ( .A(n588), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U650 ( .A(n588), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U651 ( .A(n514), .B(n421), .ZN(n359) );
  XNOR2_X1 U652 ( .A(n510), .B(n421), .ZN(n348) );
  XNOR2_X1 U653 ( .A(n513), .B(n420), .ZN(n358) );
  XNOR2_X1 U654 ( .A(n521), .B(n420), .ZN(n347) );
  XNOR2_X1 U655 ( .A(n490), .B(n418), .ZN(n356) );
  XNOR2_X1 U656 ( .A(n582), .B(b[11]), .ZN(n397) );
  XNOR2_X1 U657 ( .A(n581), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U658 ( .A(n581), .B(b[13]), .ZN(n395) );
  XNOR2_X1 U659 ( .A(n581), .B(b[14]), .ZN(n394) );
  XNOR2_X1 U660 ( .A(n513), .B(n419), .ZN(n357) );
  XNOR2_X1 U661 ( .A(n521), .B(n419), .ZN(n346) );
  XNOR2_X1 U662 ( .A(n490), .B(b[8]), .ZN(n355) );
  CLKBUF_X1 U663 ( .A(n43), .Z(n579) );
  XNOR2_X1 U664 ( .A(n581), .B(b[15]), .ZN(n393) );
  NAND2_X1 U665 ( .A1(n328), .A2(n314), .ZN(n119) );
  OAI22_X1 U666 ( .A1(n34), .A2(n339), .B1(n338), .B2(n32), .ZN(n265) );
  OAI22_X1 U667 ( .A1(n34), .A2(n340), .B1(n339), .B2(n32), .ZN(n266) );
  OAI22_X1 U668 ( .A1(n34), .A2(n342), .B1(n341), .B2(n32), .ZN(n268) );
  OAI22_X1 U669 ( .A1(n34), .A2(n341), .B1(n340), .B2(n32), .ZN(n267) );
  OAI22_X1 U670 ( .A1(n34), .A2(n343), .B1(n342), .B2(n32), .ZN(n269) );
  OAI22_X1 U671 ( .A1(n34), .A2(n501), .B1(n344), .B2(n32), .ZN(n253) );
  INV_X1 U672 ( .A(n113), .ZN(n135) );
  NOR2_X1 U673 ( .A1(n234), .A2(n257), .ZN(n113) );
  NAND2_X1 U674 ( .A1(n577), .A2(n103), .ZN(n55) );
  INV_X1 U675 ( .A(n103), .ZN(n101) );
  INV_X1 U676 ( .A(n13), .ZN(n589) );
  NOR2_X1 U677 ( .A1(n228), .A2(n231), .ZN(n105) );
  XNOR2_X1 U678 ( .A(n77), .B(n48), .ZN(product[13]) );
  XNOR2_X1 U679 ( .A(n70), .B(n47), .ZN(product[14]) );
  INV_X1 U680 ( .A(n545), .ZN(n127) );
  NOR2_X1 U681 ( .A1(n545), .A2(n85), .ZN(n80) );
  OAI21_X1 U682 ( .B1(n86), .B2(n82), .A(n83), .ZN(n81) );
  NOR2_X1 U683 ( .A1(n204), .A2(n211), .ZN(n89) );
  OAI22_X1 U684 ( .A1(n29), .A2(n346), .B1(n345), .B2(n504), .ZN(n271) );
  OAI22_X1 U685 ( .A1(n29), .A2(n350), .B1(n349), .B2(n504), .ZN(n275) );
  OAI22_X1 U686 ( .A1(n29), .A2(n347), .B1(n346), .B2(n504), .ZN(n272) );
  OAI22_X1 U687 ( .A1(n29), .A2(n348), .B1(n347), .B2(n504), .ZN(n273) );
  OAI22_X1 U688 ( .A1(n29), .A2(n349), .B1(n348), .B2(n27), .ZN(n274) );
  OAI22_X1 U689 ( .A1(n29), .A2(n351), .B1(n350), .B2(n504), .ZN(n276) );
  OAI22_X1 U690 ( .A1(n29), .A2(n352), .B1(n351), .B2(n27), .ZN(n277) );
  OR2_X1 U691 ( .A1(n578), .A2(n520), .ZN(n409) );
  INV_X1 U692 ( .A(n583), .ZN(n582) );
  OAI21_X1 U693 ( .B1(n87), .B2(n495), .A(n494), .ZN(n84) );
  NAND2_X1 U694 ( .A1(n224), .A2(n227), .ZN(n103) );
  XNOR2_X1 U695 ( .A(n581), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U696 ( .A(n581), .B(n578), .ZN(n408) );
  XNOR2_X1 U697 ( .A(n582), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U698 ( .A(n582), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U699 ( .A(n581), .B(n418), .ZN(n401) );
  XNOR2_X1 U700 ( .A(n582), .B(n421), .ZN(n404) );
  XNOR2_X1 U701 ( .A(n581), .B(n422), .ZN(n405) );
  XNOR2_X1 U702 ( .A(n581), .B(n424), .ZN(n407) );
  XNOR2_X1 U703 ( .A(n582), .B(n420), .ZN(n403) );
  XNOR2_X1 U704 ( .A(n581), .B(n423), .ZN(n406) );
  XNOR2_X1 U705 ( .A(n581), .B(n419), .ZN(n402) );
  OAI22_X1 U706 ( .A1(n541), .A2(n358), .B1(n357), .B2(n493), .ZN(n282) );
  OAI22_X1 U707 ( .A1(n542), .A2(n356), .B1(n355), .B2(n493), .ZN(n280) );
  OAI22_X1 U708 ( .A1(n542), .A2(n355), .B1(n354), .B2(n493), .ZN(n279) );
  OAI22_X1 U709 ( .A1(n542), .A2(n362), .B1(n361), .B2(n493), .ZN(n286) );
  OAI22_X1 U710 ( .A1(n542), .A2(n590), .B1(n364), .B2(n21), .ZN(n255) );
  OAI22_X1 U711 ( .A1(n541), .A2(n357), .B1(n356), .B2(n493), .ZN(n281) );
  OAI22_X1 U712 ( .A1(n541), .A2(n360), .B1(n359), .B2(n493), .ZN(n284) );
  OAI22_X1 U713 ( .A1(n541), .A2(n361), .B1(n360), .B2(n21), .ZN(n285) );
  XNOR2_X1 U714 ( .A(n587), .B(n424), .ZN(n375) );
  OAI22_X1 U715 ( .A1(n23), .A2(n363), .B1(n362), .B2(n21), .ZN(n287) );
  XNOR2_X1 U716 ( .A(n587), .B(n423), .ZN(n374) );
  OAI22_X1 U717 ( .A1(n23), .A2(n359), .B1(n358), .B2(n21), .ZN(n283) );
  XNOR2_X1 U718 ( .A(n587), .B(n421), .ZN(n372) );
  XNOR2_X1 U719 ( .A(n587), .B(n422), .ZN(n373) );
  XNOR2_X1 U720 ( .A(n587), .B(n419), .ZN(n370) );
  XNOR2_X1 U721 ( .A(n587), .B(n420), .ZN(n371) );
  NAND2_X1 U722 ( .A1(n151), .A2(n139), .ZN(n62) );
  OAI22_X1 U723 ( .A1(n18), .A2(n370), .B1(n369), .B2(n575), .ZN(n293) );
  OAI22_X1 U724 ( .A1(n18), .A2(n367), .B1(n366), .B2(n575), .ZN(n290) );
  OAI22_X1 U725 ( .A1(n18), .A2(n375), .B1(n374), .B2(n575), .ZN(n298) );
  OAI22_X1 U726 ( .A1(n18), .A2(n376), .B1(n375), .B2(n575), .ZN(n299) );
  OAI22_X1 U727 ( .A1(n18), .A2(n505), .B1(n377), .B2(n575), .ZN(n256) );
  OAI22_X1 U728 ( .A1(n18), .A2(n373), .B1(n372), .B2(n575), .ZN(n296) );
  OAI22_X1 U729 ( .A1(n18), .A2(n374), .B1(n373), .B2(n575), .ZN(n297) );
  OAI22_X1 U730 ( .A1(n18), .A2(n372), .B1(n371), .B2(n575), .ZN(n295) );
  OAI22_X1 U731 ( .A1(n18), .A2(n368), .B1(n367), .B2(n575), .ZN(n291) );
  OAI22_X1 U732 ( .A1(n18), .A2(n369), .B1(n368), .B2(n575), .ZN(n292) );
  OAI22_X1 U733 ( .A1(n18), .A2(n371), .B1(n370), .B2(n575), .ZN(n294) );
  XNOR2_X1 U734 ( .A(n584), .B(n420), .ZN(n386) );
  OAI22_X1 U735 ( .A1(n18), .A2(n366), .B1(n365), .B2(n575), .ZN(n289) );
  INV_X1 U736 ( .A(n575), .ZN(n245) );
  XNOR2_X1 U737 ( .A(n584), .B(n578), .ZN(n391) );
  XNOR2_X1 U738 ( .A(n584), .B(n423), .ZN(n389) );
  XNOR2_X1 U739 ( .A(n584), .B(n422), .ZN(n388) );
  XNOR2_X1 U740 ( .A(n584), .B(n424), .ZN(n390) );
  XNOR2_X1 U741 ( .A(n584), .B(n421), .ZN(n387) );
  XNOR2_X1 U742 ( .A(n534), .B(n55), .ZN(product[6]) );
  AOI21_X1 U743 ( .B1(n104), .B2(n577), .A(n101), .ZN(n99) );
  XOR2_X1 U744 ( .A(n56), .B(n516), .Z(product[5]) );
  OAI21_X1 U745 ( .B1(n107), .B2(n105), .A(n106), .ZN(n104) );
  XNOR2_X1 U746 ( .A(n57), .B(n112), .ZN(product[4]) );
  INV_X1 U747 ( .A(n88), .ZN(n87) );
  AOI21_X1 U748 ( .B1(n80), .B2(n503), .A(n81), .ZN(n45) );
  OAI21_X1 U749 ( .B1(n64), .B2(n517), .A(n65), .ZN(n63) );
  OAI21_X1 U750 ( .B1(n562), .B2(n498), .A(n72), .ZN(n70) );
  OAI21_X1 U751 ( .B1(n45), .B2(n78), .A(n79), .ZN(n77) );
  XOR2_X1 U752 ( .A(n552), .B(n52), .Z(product[9]) );
  XNOR2_X1 U753 ( .A(n546), .B(n53), .ZN(product[8]) );
  AOI21_X1 U754 ( .B1(n96), .B2(n567), .A(n93), .ZN(n91) );
  XOR2_X1 U755 ( .A(n58), .B(n115), .Z(product[3]) );
  OAI22_X1 U756 ( .A1(n561), .A2(n395), .B1(n394), .B2(n535), .ZN(n316) );
  OAI22_X1 U757 ( .A1(n6), .A2(n394), .B1(n393), .B2(n535), .ZN(n315) );
  OAI22_X1 U758 ( .A1(n560), .A2(n396), .B1(n395), .B2(n535), .ZN(n317) );
  OAI22_X1 U759 ( .A1(n6), .A2(n397), .B1(n396), .B2(n535), .ZN(n318) );
  OAI22_X1 U760 ( .A1(n560), .A2(n398), .B1(n397), .B2(n535), .ZN(n319) );
  OAI22_X1 U761 ( .A1(n6), .A2(n400), .B1(n399), .B2(n535), .ZN(n321) );
  OAI22_X1 U762 ( .A1(n561), .A2(n399), .B1(n398), .B2(n535), .ZN(n320) );
  OAI22_X1 U763 ( .A1(n561), .A2(n401), .B1(n400), .B2(n535), .ZN(n322) );
  OAI22_X1 U764 ( .A1(n6), .A2(n402), .B1(n401), .B2(n535), .ZN(n323) );
  NAND2_X1 U765 ( .A1(n329), .A2(n258), .ZN(n122) );
  OAI22_X1 U766 ( .A1(n404), .A2(n561), .B1(n403), .B2(n535), .ZN(n325) );
  OAI22_X1 U767 ( .A1(n6), .A2(n403), .B1(n402), .B2(n535), .ZN(n324) );
  OAI22_X1 U768 ( .A1(n6), .A2(n406), .B1(n405), .B2(n535), .ZN(n327) );
  OAI22_X1 U769 ( .A1(n560), .A2(n405), .B1(n404), .B2(n580), .ZN(n326) );
  OAI22_X1 U770 ( .A1(n560), .A2(n407), .B1(n406), .B2(n535), .ZN(n328) );
  OAI22_X1 U771 ( .A1(n560), .A2(n408), .B1(n407), .B2(n535), .ZN(n329) );
  OAI22_X1 U772 ( .A1(n561), .A2(n520), .B1(n409), .B2(n535), .ZN(n258) );
  XOR2_X1 U773 ( .A(n543), .B(n54), .Z(product[7]) );
  OAI22_X1 U774 ( .A1(n555), .A2(n379), .B1(n378), .B2(n550), .ZN(n301) );
  OAI22_X1 U775 ( .A1(n556), .A2(n380), .B1(n379), .B2(n550), .ZN(n302) );
  OAI22_X1 U776 ( .A1(n555), .A2(n385), .B1(n384), .B2(n550), .ZN(n307) );
  OAI22_X1 U777 ( .A1(n556), .A2(n382), .B1(n381), .B2(n550), .ZN(n304) );
  OAI22_X1 U778 ( .A1(n555), .A2(n381), .B1(n380), .B2(n550), .ZN(n303) );
  NAND2_X1 U779 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U780 ( .A1(n554), .A2(n383), .B1(n382), .B2(n576), .ZN(n305) );
  OAI22_X1 U781 ( .A1(n556), .A2(n384), .B1(n383), .B2(n550), .ZN(n306) );
  OAI22_X1 U782 ( .A1(n555), .A2(n386), .B1(n385), .B2(n550), .ZN(n308) );
  OAI22_X1 U783 ( .A1(n555), .A2(n387), .B1(n386), .B2(n550), .ZN(n309) );
  OAI22_X1 U784 ( .A1(n556), .A2(n508), .B1(n392), .B2(n550), .ZN(n257) );
  OAI22_X1 U785 ( .A1(n554), .A2(n389), .B1(n388), .B2(n576), .ZN(n311) );
  OAI22_X1 U786 ( .A1(n555), .A2(n388), .B1(n387), .B2(n550), .ZN(n310) );
  OAI22_X1 U787 ( .A1(n556), .A2(n390), .B1(n389), .B2(n576), .ZN(n312) );
  INV_X1 U788 ( .A(n550), .ZN(n247) );
  OAI22_X1 U789 ( .A1(n556), .A2(n391), .B1(n390), .B2(n576), .ZN(n313) );
  INV_X1 U790 ( .A(n586), .ZN(n585) );
  INV_X1 U791 ( .A(n589), .ZN(n588) );
  INV_X1 U792 ( .A(n31), .ZN(n594) );
  INV_X1 U793 ( .A(n36), .ZN(n596) );
  INV_X1 U794 ( .A(n598), .ZN(n597) );
  INV_X1 U795 ( .A(n40), .ZN(n598) );
  XOR2_X1 U796 ( .A(n259), .B(n251), .Z(n148) );
  XOR2_X1 U797 ( .A(n279), .B(n289), .Z(n146) );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_8_DW01_add_2 ( A, B, CI, 
        SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n8, n9, n10, n11, n12, n13, n14, n15, n16, n19,
         n20, n22, n24, n25, n26, n27, n29, n30, n31, n32, n33, n34, n35, n36,
         n38, n39, n40, n44, n45, n47, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n65, n67, n68, n69, n70, n71, n73,
         n75, n76, n77, n78, n79, n81, n83, n84, n86, n90, n91, n95, n96, n98,
         n100, n157, n158, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184;

  XNOR2_X1 U122 ( .A(n38), .B(n6), .ZN(SUM[11]) );
  BUF_X1 U123 ( .A(n36), .Z(n157) );
  OR2_X2 U124 ( .A1(A[13]), .A2(B[13]), .ZN(n164) );
  OR2_X1 U125 ( .A1(A[8]), .A2(B[8]), .ZN(n158) );
  AND2_X1 U126 ( .A1(n177), .A2(n86), .ZN(SUM[0]) );
  NOR2_X1 U127 ( .A1(A[8]), .A2(B[8]), .ZN(n160) );
  NOR2_X1 U128 ( .A1(A[8]), .A2(B[8]), .ZN(n54) );
  XNOR2_X1 U129 ( .A(n45), .B(n161), .ZN(SUM[10]) );
  AND2_X1 U130 ( .A1(n44), .A2(n174), .ZN(n161) );
  NAND2_X1 U131 ( .A1(n163), .A2(n164), .ZN(n162) );
  OR2_X1 U132 ( .A1(A[14]), .A2(B[14]), .ZN(n163) );
  INV_X1 U133 ( .A(n91), .ZN(n165) );
  NOR2_X1 U134 ( .A1(A[11]), .A2(B[11]), .ZN(n35) );
  AOI21_X1 U135 ( .B1(n183), .B2(n47), .A(n184), .ZN(n166) );
  INV_X1 U136 ( .A(n38), .ZN(n167) );
  OR2_X1 U137 ( .A1(A[15]), .A2(B[15]), .ZN(n168) );
  OAI21_X1 U138 ( .B1(n39), .B2(n51), .A(n40), .ZN(n169) );
  AND2_X1 U139 ( .A1(A[9]), .A2(B[9]), .ZN(n47) );
  NOR2_X1 U140 ( .A1(A[12]), .A2(B[12]), .ZN(n170) );
  NOR2_X1 U141 ( .A1(B[12]), .A2(A[12]), .ZN(n32) );
  INV_X1 U142 ( .A(n164), .ZN(n171) );
  BUF_X1 U143 ( .A(n29), .Z(n172) );
  OAI21_X1 U144 ( .B1(n32), .B2(n36), .A(n33), .ZN(n173) );
  NOR2_X1 U145 ( .A1(A[14]), .A2(B[14]), .ZN(n25) );
  OR2_X1 U146 ( .A1(A[10]), .A2(B[10]), .ZN(n174) );
  OR2_X1 U147 ( .A1(A[10]), .A2(B[10]), .ZN(n183) );
  AOI21_X1 U148 ( .B1(n169), .B2(n30), .A(n31), .ZN(n175) );
  AOI21_X1 U149 ( .B1(n169), .B2(n30), .A(n173), .ZN(n176) );
  OR2_X1 U150 ( .A1(A[0]), .A2(B[0]), .ZN(n177) );
  AOI21_X1 U151 ( .B1(n180), .B2(n76), .A(n73), .ZN(n71) );
  INV_X1 U152 ( .A(n75), .ZN(n73) );
  OAI21_X1 U153 ( .B1(n79), .B2(n77), .A(n78), .ZN(n76) );
  AOI21_X1 U154 ( .B1(n181), .B2(n68), .A(n65), .ZN(n63) );
  INV_X1 U155 ( .A(n67), .ZN(n65) );
  INV_X1 U156 ( .A(n24), .ZN(n22) );
  OAI21_X1 U157 ( .B1(n71), .B2(n69), .A(n70), .ZN(n68) );
  AOI21_X1 U158 ( .B1(n50), .B2(n178), .A(n47), .ZN(n45) );
  INV_X1 U159 ( .A(n86), .ZN(n84) );
  OAI21_X1 U160 ( .B1(n59), .B2(n57), .A(n58), .ZN(n56) );
  AOI21_X1 U161 ( .B1(n179), .B2(n84), .A(n81), .ZN(n79) );
  INV_X1 U162 ( .A(n83), .ZN(n81) );
  NAND2_X1 U163 ( .A1(n98), .A2(n70), .ZN(n13) );
  INV_X1 U164 ( .A(n69), .ZN(n98) );
  NAND2_X1 U165 ( .A1(n158), .A2(n55), .ZN(n9) );
  NAND2_X1 U166 ( .A1(n164), .A2(n172), .ZN(n4) );
  NAND2_X1 U167 ( .A1(n180), .A2(n75), .ZN(n14) );
  NAND2_X1 U168 ( .A1(n95), .A2(n58), .ZN(n10) );
  INV_X1 U169 ( .A(n57), .ZN(n95) );
  NAND2_X1 U170 ( .A1(n178), .A2(n49), .ZN(n8) );
  NAND2_X1 U171 ( .A1(n100), .A2(n78), .ZN(n15) );
  INV_X1 U172 ( .A(n77), .ZN(n100) );
  NAND2_X1 U173 ( .A1(n181), .A2(n67), .ZN(n12) );
  NAND2_X1 U174 ( .A1(n179), .A2(n83), .ZN(n16) );
  NAND2_X1 U175 ( .A1(n96), .A2(n62), .ZN(n11) );
  INV_X1 U176 ( .A(n61), .ZN(n96) );
  NAND2_X1 U177 ( .A1(n163), .A2(n26), .ZN(n3) );
  XNOR2_X1 U178 ( .A(n34), .B(n5), .ZN(SUM[12]) );
  NAND2_X1 U179 ( .A1(n90), .A2(n33), .ZN(n5) );
  NAND2_X1 U180 ( .A1(n91), .A2(n36), .ZN(n6) );
  XNOR2_X1 U181 ( .A(n50), .B(n8), .ZN(SUM[9]) );
  XOR2_X1 U182 ( .A(n59), .B(n10), .Z(SUM[7]) );
  XNOR2_X1 U183 ( .A(n14), .B(n76), .ZN(SUM[3]) );
  XOR2_X1 U184 ( .A(n15), .B(n79), .Z(SUM[2]) );
  NOR2_X1 U185 ( .A1(A[7]), .A2(B[7]), .ZN(n57) );
  OR2_X1 U186 ( .A1(A[9]), .A2(B[9]), .ZN(n178) );
  NOR2_X1 U187 ( .A1(A[2]), .A2(B[2]), .ZN(n77) );
  NOR2_X1 U188 ( .A1(A[4]), .A2(B[4]), .ZN(n69) );
  NAND2_X1 U189 ( .A1(A[13]), .A2(B[13]), .ZN(n29) );
  NAND2_X1 U190 ( .A1(A[11]), .A2(B[11]), .ZN(n36) );
  OR2_X1 U191 ( .A1(A[1]), .A2(B[1]), .ZN(n179) );
  OR2_X1 U192 ( .A1(A[3]), .A2(B[3]), .ZN(n180) );
  NAND2_X1 U193 ( .A1(A[14]), .A2(B[14]), .ZN(n26) );
  NAND2_X1 U194 ( .A1(A[12]), .A2(B[12]), .ZN(n33) );
  XNOR2_X1 U195 ( .A(n56), .B(n9), .ZN(SUM[8]) );
  XNOR2_X1 U196 ( .A(n16), .B(n84), .ZN(SUM[1]) );
  NOR2_X1 U197 ( .A1(A[6]), .A2(B[6]), .ZN(n61) );
  NAND2_X1 U198 ( .A1(A[7]), .A2(B[7]), .ZN(n58) );
  OR2_X1 U199 ( .A1(A[5]), .A2(B[5]), .ZN(n181) );
  NAND2_X1 U200 ( .A1(A[2]), .A2(B[2]), .ZN(n78) );
  NAND2_X1 U201 ( .A1(A[4]), .A2(B[4]), .ZN(n70) );
  NAND2_X1 U202 ( .A1(A[1]), .A2(B[1]), .ZN(n83) );
  NAND2_X1 U203 ( .A1(A[5]), .A2(B[5]), .ZN(n67) );
  NAND2_X1 U204 ( .A1(A[0]), .A2(B[0]), .ZN(n86) );
  NAND2_X1 U205 ( .A1(A[9]), .A2(B[9]), .ZN(n49) );
  NAND2_X1 U206 ( .A1(A[6]), .A2(B[6]), .ZN(n62) );
  NAND2_X1 U207 ( .A1(A[8]), .A2(B[8]), .ZN(n55) );
  XNOR2_X1 U208 ( .A(n12), .B(n68), .ZN(SUM[5]) );
  XOR2_X1 U209 ( .A(n13), .B(n71), .Z(SUM[4]) );
  NAND2_X1 U210 ( .A1(n168), .A2(n19), .ZN(n2) );
  AOI21_X1 U211 ( .B1(n52), .B2(n60), .A(n53), .ZN(n182) );
  INV_X1 U212 ( .A(n182), .ZN(n50) );
  AOI21_X1 U213 ( .B1(n52), .B2(n60), .A(n53), .ZN(n51) );
  INV_X1 U214 ( .A(n60), .ZN(n59) );
  INV_X1 U215 ( .A(n184), .ZN(n44) );
  NOR2_X1 U216 ( .A1(n160), .A2(n57), .ZN(n52) );
  OAI21_X1 U217 ( .B1(n54), .B2(n58), .A(n55), .ZN(n53) );
  AOI21_X1 U218 ( .B1(n183), .B2(n47), .A(n184), .ZN(n40) );
  AND2_X1 U219 ( .A1(A[10]), .A2(B[10]), .ZN(n184) );
  INV_X1 U220 ( .A(n170), .ZN(n90) );
  OAI21_X1 U221 ( .B1(n170), .B2(n36), .A(n33), .ZN(n31) );
  XOR2_X1 U222 ( .A(n11), .B(n63), .Z(SUM[6]) );
  OAI21_X1 U223 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  NAND2_X1 U224 ( .A1(A[3]), .A2(B[3]), .ZN(n75) );
  OAI21_X1 U225 ( .B1(n167), .B2(n165), .A(n157), .ZN(n34) );
  INV_X1 U226 ( .A(n35), .ZN(n91) );
  NOR2_X1 U227 ( .A1(n32), .A2(n35), .ZN(n30) );
  OAI21_X1 U228 ( .B1(n25), .B2(n29), .A(n26), .ZN(n24) );
  NAND2_X1 U229 ( .A1(A[15]), .A2(B[15]), .ZN(n19) );
  OAI21_X1 U230 ( .B1(n39), .B2(n51), .A(n166), .ZN(n38) );
  NAND2_X1 U231 ( .A1(n174), .A2(n178), .ZN(n39) );
  XNOR2_X1 U232 ( .A(n20), .B(n2), .ZN(SUM[15]) );
  XNOR2_X1 U233 ( .A(n27), .B(n3), .ZN(SUM[14]) );
  XOR2_X1 U234 ( .A(n4), .B(n175), .Z(SUM[13]) );
  OAI21_X1 U235 ( .B1(n175), .B2(n171), .A(n172), .ZN(n27) );
  OAI21_X1 U236 ( .B1(n176), .B2(n162), .A(n22), .ZN(n20) );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_8 ( clk, clear_acc, 
        data_out_x, data_out, data_out_w, data_out_b, wr_en_y, m_valid, 
        m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [4:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
         N39, N40, N41, N42, N43, N44, n1, n2, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n85, n102, n111, n112, n113, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n22), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n227), .CK(clk), .Q(n26) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n228), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n229), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n230), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n231), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n232), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n233), .CK(clk), .Q(n34) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n234), .CK(clk), .Q(n35) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n235), .CK(clk), .Q(n36) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n236), .CK(clk), .Q(n37) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n237), .CK(clk), .Q(n38) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n238), .CK(clk), .Q(n39) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n239), .CK(clk), .Q(n40) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n240), .CK(clk), .Q(n41) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n241), .CK(clk), .Q(n42) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n242), .CK(clk), .Q(n44) );
  DFF_X1 \f_reg[0]  ( .D(n113), .CK(clk), .Q(f[0]), .QN(n215) );
  DFF_X1 \f_reg[1]  ( .D(n112), .CK(clk), .Q(f[1]), .QN(n216) );
  DFF_X1 \f_reg[2]  ( .D(n111), .CK(clk), .Q(f[2]), .QN(n217) );
  DFF_X1 \f_reg[3]  ( .D(n102), .CK(clk), .Q(f[3]), .QN(n218) );
  DFF_X1 \f_reg[7]  ( .D(n81), .CK(clk), .Q(f[7]), .QN(n219) );
  DFF_X1 \f_reg[8]  ( .D(n80), .CK(clk), .Q(f[8]), .QN(n220) );
  DFF_X1 \f_reg[9]  ( .D(n79), .CK(clk), .Q(f[9]), .QN(n221) );
  DFF_X1 \f_reg[10]  ( .D(n78), .CK(clk), .Q(n53), .QN(n222) );
  DFF_X1 \f_reg[11]  ( .D(n77), .CK(clk), .Q(n51), .QN(n223) );
  DFF_X1 \f_reg[12]  ( .D(n2), .CK(clk), .Q(n50), .QN(n224) );
  DFF_X1 \f_reg[13]  ( .D(n16), .CK(clk), .Q(n49), .QN(n225) );
  DFF_X1 \f_reg[14]  ( .D(n7), .CK(clk), .Q(n48), .QN(n226) );
  DFF_X1 \data_out_reg[15]  ( .D(n167), .CK(clk), .Q(data_out[15]), .QN(n198)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n168), .CK(clk), .Q(data_out[14]), .QN(n197)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n169), .CK(clk), .Q(data_out[13]), .QN(n196)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n170), .CK(clk), .Q(data_out[12]), .QN(n195)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n171), .CK(clk), .Q(data_out[11]), .QN(n194)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n172), .CK(clk), .Q(data_out[10]), .QN(n193)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n173), .CK(clk), .Q(data_out[9]), .QN(n192) );
  DFF_X1 \data_out_reg[8]  ( .D(n174), .CK(clk), .Q(data_out[8]), .QN(n191) );
  DFF_X1 \data_out_reg[7]  ( .D(n175), .CK(clk), .Q(data_out[7]), .QN(n190) );
  DFF_X1 \data_out_reg[6]  ( .D(n176), .CK(clk), .Q(data_out[6]), .QN(n189) );
  DFF_X1 \data_out_reg[5]  ( .D(n177), .CK(clk), .Q(data_out[5]), .QN(n188) );
  DFF_X1 \data_out_reg[4]  ( .D(n178), .CK(clk), .Q(data_out[4]), .QN(n187) );
  DFF_X1 \data_out_reg[3]  ( .D(n179), .CK(clk), .Q(data_out[3]), .QN(n186) );
  DFF_X1 \data_out_reg[2]  ( .D(n180), .CK(clk), .Q(data_out[2]), .QN(n185) );
  DFF_X1 \data_out_reg[1]  ( .D(n181), .CK(clk), .Q(data_out[1]), .QN(n184) );
  DFF_X1 \data_out_reg[0]  ( .D(n182), .CK(clk), .Q(data_out[0]), .QN(n183) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_8_DW_mult_tc_1 mult_2021 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_8_DW01_add_2 add_2022 ( .A({n205, 
        n204, n203, n202, n201, n200, n214, n213, n212, n211, n210, n209, n208, 
        n207, n206, n199}), .B({f[15], n48, n49, n50, n51, n53, f[9:0]}), .CI(
        1'b0), .SUM(adder) );
  DFF_X1 delay_reg ( .D(n166), .CK(clk), .Q(n14), .QN(n243) );
  DFF_X1 \f_reg[4]  ( .D(n85), .CK(clk), .Q(f[4]), .QN(n66) );
  DFF_X1 \f_reg[5]  ( .D(n83), .CK(clk), .Q(f[5]), .QN(n67) );
  DFF_X1 \f_reg[6]  ( .D(n82), .CK(clk), .Q(f[6]), .QN(n68) );
  DFF_X1 \f_reg[15]  ( .D(n76), .CK(clk), .Q(f[15]), .QN(n73) );
  CLKBUF_X1 U3 ( .A(N41), .Z(n1) );
  MUX2_X2 U4 ( .A(N40), .B(n32), .S(n14), .Z(n201) );
  AND2_X1 U5 ( .A1(n47), .A2(n23), .ZN(n15) );
  NAND3_X1 U6 ( .A1(n5), .A2(n4), .A3(n6), .ZN(n2) );
  MUX2_X2 U8 ( .A(n35), .B(N37), .S(n243), .Z(n213) );
  NAND2_X1 U9 ( .A1(data_out_b[12]), .A2(n21), .ZN(n4) );
  NAND2_X1 U10 ( .A1(adder[12]), .A2(n15), .ZN(n5) );
  NAND2_X1 U11 ( .A1(n64), .A2(n50), .ZN(n6) );
  INV_X1 U12 ( .A(n47), .ZN(n64) );
  NAND3_X1 U13 ( .A1(n12), .A2(n11), .A3(n13), .ZN(n7) );
  OAI222_X1 U14 ( .A1(n47), .A2(n73), .B1(n8), .B2(n23), .C1(n9), .C2(n10), 
        .ZN(n76) );
  INV_X1 U15 ( .A(data_out_b[15]), .ZN(n8) );
  INV_X1 U16 ( .A(adder[15]), .ZN(n9) );
  INV_X1 U17 ( .A(n15), .ZN(n10) );
  NAND2_X1 U18 ( .A1(data_out_b[14]), .A2(n21), .ZN(n11) );
  NAND2_X1 U19 ( .A1(adder[14]), .A2(n15), .ZN(n12) );
  NAND2_X1 U20 ( .A1(n64), .A2(n48), .ZN(n13) );
  MUX2_X2 U21 ( .A(n29), .B(N41), .S(n243), .Z(n202) );
  MUX2_X2 U22 ( .A(n28), .B(N42), .S(n243), .Z(n203) );
  MUX2_X2 U23 ( .A(N39), .B(n33), .S(n14), .Z(n200) );
  MUX2_X2 U24 ( .A(n27), .B(N43), .S(n243), .Z(n204) );
  NAND2_X1 U25 ( .A1(n166), .A2(n20), .ZN(n245) );
  INV_X1 U26 ( .A(clear_acc), .ZN(n23) );
  INV_X1 U27 ( .A(n25), .ZN(n43) );
  OAI22_X1 U28 ( .A1(n186), .A2(n245), .B1(n218), .B2(n244), .ZN(n179) );
  OAI22_X1 U29 ( .A1(n187), .A2(n245), .B1(n66), .B2(n244), .ZN(n178) );
  OAI22_X1 U30 ( .A1(n188), .A2(n245), .B1(n67), .B2(n244), .ZN(n177) );
  OAI22_X1 U31 ( .A1(n189), .A2(n245), .B1(n68), .B2(n244), .ZN(n176) );
  OAI22_X1 U32 ( .A1(n190), .A2(n245), .B1(n219), .B2(n244), .ZN(n175) );
  OAI22_X1 U33 ( .A1(n191), .A2(n245), .B1(n220), .B2(n244), .ZN(n174) );
  OAI22_X1 U34 ( .A1(n192), .A2(n245), .B1(n221), .B2(n244), .ZN(n173) );
  NAND3_X1 U35 ( .A1(n18), .A2(n17), .A3(n19), .ZN(n16) );
  MUX2_X1 U36 ( .A(n40), .B(N32), .S(n243), .Z(n208) );
  NAND2_X1 U37 ( .A1(data_out_b[13]), .A2(n21), .ZN(n17) );
  NAND2_X1 U38 ( .A1(adder[13]), .A2(n15), .ZN(n18) );
  NAND2_X1 U39 ( .A1(n64), .A2(n49), .ZN(n19) );
  INV_X1 U40 ( .A(n23), .ZN(n21) );
  INV_X1 U41 ( .A(wr_en_y), .ZN(n20) );
  INV_X1 U42 ( .A(n23), .ZN(n22) );
  INV_X1 U43 ( .A(m_ready), .ZN(n24) );
  NAND2_X1 U44 ( .A1(m_valid), .A2(n24), .ZN(n45) );
  OAI21_X1 U45 ( .B1(sel[4]), .B2(n75), .A(n45), .ZN(n166) );
  NAND2_X1 U46 ( .A1(clear_acc_delay), .A2(n243), .ZN(n25) );
  MUX2_X1 U47 ( .A(n26), .B(N44), .S(n43), .Z(n227) );
  MUX2_X1 U48 ( .A(n26), .B(N44), .S(n243), .Z(n205) );
  MUX2_X1 U49 ( .A(n27), .B(N43), .S(n43), .Z(n228) );
  MUX2_X1 U50 ( .A(n28), .B(N42), .S(n43), .Z(n229) );
  MUX2_X1 U51 ( .A(n29), .B(n1), .S(n43), .Z(n230) );
  MUX2_X1 U52 ( .A(n32), .B(N40), .S(n43), .Z(n231) );
  MUX2_X1 U53 ( .A(n33), .B(N39), .S(n43), .Z(n232) );
  MUX2_X1 U54 ( .A(n34), .B(N38), .S(n43), .Z(n233) );
  MUX2_X1 U55 ( .A(n34), .B(N38), .S(n243), .Z(n214) );
  MUX2_X1 U56 ( .A(n35), .B(N37), .S(n43), .Z(n234) );
  MUX2_X1 U57 ( .A(n36), .B(N36), .S(n43), .Z(n235) );
  MUX2_X1 U58 ( .A(n36), .B(N36), .S(n243), .Z(n212) );
  MUX2_X1 U59 ( .A(n37), .B(N35), .S(n43), .Z(n236) );
  MUX2_X1 U60 ( .A(n37), .B(N35), .S(n243), .Z(n211) );
  MUX2_X1 U61 ( .A(n38), .B(N34), .S(n43), .Z(n237) );
  MUX2_X1 U62 ( .A(n38), .B(N34), .S(n243), .Z(n210) );
  MUX2_X1 U63 ( .A(n39), .B(N33), .S(n43), .Z(n238) );
  MUX2_X1 U64 ( .A(n39), .B(N33), .S(n243), .Z(n209) );
  MUX2_X1 U65 ( .A(n40), .B(N32), .S(n43), .Z(n239) );
  MUX2_X1 U66 ( .A(n41), .B(N31), .S(n43), .Z(n240) );
  MUX2_X1 U67 ( .A(n41), .B(N31), .S(n243), .Z(n207) );
  MUX2_X1 U68 ( .A(n42), .B(N30), .S(n43), .Z(n241) );
  MUX2_X1 U69 ( .A(n42), .B(N30), .S(n243), .Z(n206) );
  MUX2_X1 U70 ( .A(n44), .B(N29), .S(n43), .Z(n242) );
  MUX2_X1 U71 ( .A(n44), .B(N29), .S(n243), .Z(n199) );
  INV_X1 U72 ( .A(n45), .ZN(n46) );
  OAI21_X1 U73 ( .B1(n46), .B2(n14), .A(n23), .ZN(n47) );
  AOI222_X1 U74 ( .A1(data_out_b[11]), .A2(n21), .B1(adder[11]), .B2(n15), 
        .C1(n64), .C2(n51), .ZN(n52) );
  INV_X1 U75 ( .A(n52), .ZN(n77) );
  AOI222_X1 U76 ( .A1(data_out_b[10]), .A2(n21), .B1(adder[10]), .B2(n15), 
        .C1(n64), .C2(n53), .ZN(n54) );
  INV_X1 U77 ( .A(n54), .ZN(n78) );
  AOI222_X1 U78 ( .A1(data_out_b[8]), .A2(n21), .B1(adder[8]), .B2(n15), .C1(
        n64), .C2(f[8]), .ZN(n55) );
  INV_X1 U79 ( .A(n55), .ZN(n80) );
  AOI222_X1 U80 ( .A1(data_out_b[7]), .A2(n21), .B1(adder[7]), .B2(n15), .C1(
        n64), .C2(f[7]), .ZN(n56) );
  INV_X1 U81 ( .A(n56), .ZN(n81) );
  AOI222_X1 U82 ( .A1(data_out_b[6]), .A2(n21), .B1(adder[6]), .B2(n15), .C1(
        n64), .C2(f[6]), .ZN(n57) );
  INV_X1 U83 ( .A(n57), .ZN(n82) );
  AOI222_X1 U84 ( .A1(data_out_b[5]), .A2(n21), .B1(adder[5]), .B2(n15), .C1(
        n64), .C2(f[5]), .ZN(n58) );
  INV_X1 U85 ( .A(n58), .ZN(n83) );
  AOI222_X1 U86 ( .A1(data_out_b[4]), .A2(n21), .B1(adder[4]), .B2(n15), .C1(
        n64), .C2(f[4]), .ZN(n59) );
  INV_X1 U87 ( .A(n59), .ZN(n85) );
  AOI222_X1 U88 ( .A1(data_out_b[3]), .A2(n21), .B1(adder[3]), .B2(n15), .C1(
        n64), .C2(f[3]), .ZN(n60) );
  INV_X1 U89 ( .A(n60), .ZN(n102) );
  AOI222_X1 U90 ( .A1(data_out_b[2]), .A2(n22), .B1(adder[2]), .B2(n15), .C1(
        n64), .C2(f[2]), .ZN(n61) );
  INV_X1 U91 ( .A(n61), .ZN(n111) );
  AOI222_X1 U92 ( .A1(data_out_b[1]), .A2(n22), .B1(adder[1]), .B2(n15), .C1(
        n64), .C2(f[1]), .ZN(n62) );
  INV_X1 U93 ( .A(n62), .ZN(n112) );
  AOI222_X1 U94 ( .A1(data_out_b[0]), .A2(n22), .B1(adder[0]), .B2(n15), .C1(
        n64), .C2(f[0]), .ZN(n63) );
  INV_X1 U95 ( .A(n63), .ZN(n113) );
  AOI222_X1 U96 ( .A1(data_out_b[9]), .A2(n22), .B1(adder[9]), .B2(n15), .C1(
        n64), .C2(f[9]), .ZN(n65) );
  INV_X1 U97 ( .A(n65), .ZN(n79) );
  NOR4_X1 U98 ( .A1(n51), .A2(n50), .A3(n49), .A4(n48), .ZN(n72) );
  NOR4_X1 U99 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n53), .ZN(n71) );
  NAND4_X1 U100 ( .A1(n68), .A2(n67), .A3(n66), .A4(n218), .ZN(n69) );
  NOR4_X1 U101 ( .A1(n69), .A2(f[0]), .A3(f[1]), .A4(f[2]), .ZN(n70) );
  NAND3_X1 U102 ( .A1(n72), .A2(n71), .A3(n70), .ZN(n74) );
  NAND3_X1 U103 ( .A1(wr_en_y), .A2(n74), .A3(n73), .ZN(n244) );
  OAI22_X1 U104 ( .A1(n183), .A2(n245), .B1(n215), .B2(n244), .ZN(n182) );
  OAI22_X1 U105 ( .A1(n184), .A2(n245), .B1(n216), .B2(n244), .ZN(n181) );
  OAI22_X1 U106 ( .A1(n185), .A2(n245), .B1(n217), .B2(n244), .ZN(n180) );
  OAI22_X1 U107 ( .A1(n193), .A2(n245), .B1(n222), .B2(n244), .ZN(n172) );
  OAI22_X1 U108 ( .A1(n194), .A2(n245), .B1(n223), .B2(n244), .ZN(n171) );
  OAI22_X1 U109 ( .A1(n195), .A2(n245), .B1(n224), .B2(n244), .ZN(n170) );
  OAI22_X1 U110 ( .A1(n196), .A2(n245), .B1(n225), .B2(n244), .ZN(n169) );
  OAI22_X1 U111 ( .A1(n197), .A2(n245), .B1(n226), .B2(n244), .ZN(n168) );
  OAI22_X1 U112 ( .A1(n198), .A2(n245), .B1(n73), .B2(n244), .ZN(n167) );
  AND4_X1 U113 ( .A1(sel[3]), .A2(sel[2]), .A3(sel[1]), .A4(sel[0]), .ZN(n75)
         );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_7_DW_mult_tc_1 ( a, b, 
        product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n9, n12, n13, n16, n18, n19, n21, n23, n25, n27, n29, n31,
         n32, n34, n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n50,
         n53, n54, n55, n56, n57, n58, n59, n62, n63, n64, n65, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n93, n95, n96, n97, n98, n99, n103,
         n104, n105, n106, n107, n111, n112, n113, n114, n115, n117, n119,
         n120, n122, n127, n128, n133, n135, n139, n141, n142, n143, n144,
         n145, n146, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n245, n249, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n418, n419, n420,
         n421, n422, n423, n424, n426, n427, n429, n432, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U148 ( .A(n265), .B(n144), .Z(n145) );
  XOR2_X1 U152 ( .A(n301), .B(n148), .Z(n149) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n263), .CI(n291), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n317), .B(n252), .CO(n173), .S(n174) );
  FA_X1 U167 ( .A(n180), .B(n187), .CI(n178), .CO(n175), .S(n176) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U170 ( .A(n268), .B(n292), .CI(n274), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U173 ( .A(n199), .B(n201), .CI(n192), .CO(n187), .S(n188) );
  FA_X1 U174 ( .A(n275), .B(n293), .CI(n194), .CO(n189), .S(n190) );
  HA_X1 U176 ( .A(n319), .B(n269), .CO(n193), .S(n194) );
  FA_X1 U179 ( .A(n276), .B(n294), .CI(n284), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n320), .B(n270), .CI(n306), .CO(n201), .S(n202) );
  FA_X1 U182 ( .A(n215), .B(n307), .CI(n210), .CO(n205), .S(n206) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U185 ( .A(n216), .B(n219), .CI(n214), .CO(n211), .S(n212) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n322), .B(n278), .CI(n308), .CO(n215), .S(n216) );
  FA_X1 U188 ( .A(n225), .B(n222), .CI(n220), .CO(n217), .S(n218) );
  FA_X1 U189 ( .A(n297), .B(n255), .CI(n309), .CO(n219), .S(n220) );
  HA_X1 U190 ( .A(n287), .B(n323), .CO(n221), .S(n222) );
  FA_X1 U192 ( .A(n324), .B(n288), .CI(n310), .CO(n225), .S(n226) );
  HA_X1 U194 ( .A(n311), .B(n325), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n326), .B(n300), .CI(n312), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  XOR2_X1 U414 ( .A(n616), .B(a[4]), .Z(n490) );
  AND2_X1 U415 ( .A1(n224), .A2(n227), .ZN(n491) );
  XNOR2_X1 U416 ( .A(n590), .B(n492), .ZN(product[9]) );
  AND2_X1 U417 ( .A1(n576), .A2(n90), .ZN(n492) );
  OR2_X1 U418 ( .A1(n218), .A2(n223), .ZN(n493) );
  XOR2_X1 U419 ( .A(n624), .B(a[10]), .Z(n552) );
  BUF_X1 U420 ( .A(n112), .Z(n494) );
  XNOR2_X1 U421 ( .A(n45), .B(n495), .ZN(product[12]) );
  AND2_X1 U422 ( .A1(n527), .A2(n79), .ZN(n495) );
  OR2_X1 U423 ( .A1(n577), .A2(n587), .ZN(n6) );
  CLKBUF_X3 U424 ( .A(n9), .Z(n605) );
  NOR2_X1 U425 ( .A1(n218), .A2(n223), .ZN(n97) );
  OR2_X1 U426 ( .A1(n164), .A2(n175), .ZN(n496) );
  OR2_X1 U427 ( .A1(n329), .A2(n258), .ZN(n497) );
  OR2_X1 U428 ( .A1(n232), .A2(n233), .ZN(n498) );
  BUF_X2 U429 ( .A(n16), .Z(n603) );
  XOR2_X1 U430 ( .A(n626), .B(a[14]), .Z(n41) );
  CLKBUF_X1 U431 ( .A(n95), .Z(n499) );
  XNOR2_X1 U432 ( .A(n500), .B(n166), .ZN(n164) );
  XNOR2_X1 U433 ( .A(n177), .B(n168), .ZN(n500) );
  BUF_X1 U434 ( .A(n9), .Z(n604) );
  BUF_X1 U435 ( .A(n543), .Z(n590) );
  XNOR2_X1 U436 ( .A(n226), .B(n501), .ZN(n224) );
  XNOR2_X1 U437 ( .A(n229), .B(n298), .ZN(n501) );
  OR2_X2 U438 ( .A1(n577), .A2(n587), .ZN(n524) );
  OAI21_X1 U439 ( .B1(n91), .B2(n89), .A(n90), .ZN(n502) );
  AOI21_X1 U440 ( .B1(n498), .B2(n112), .A(n579), .ZN(n503) );
  INV_X1 U441 ( .A(n535), .ZN(n504) );
  NAND2_X1 U442 ( .A1(n427), .A2(n37), .ZN(n505) );
  XOR2_X1 U443 ( .A(n625), .B(a[14]), .Z(n506) );
  XOR2_X1 U444 ( .A(n170), .B(n172), .Z(n507) );
  XOR2_X1 U445 ( .A(n507), .B(n179), .Z(n166) );
  NAND2_X1 U446 ( .A1(n170), .A2(n172), .ZN(n508) );
  NAND2_X1 U447 ( .A1(n170), .A2(n179), .ZN(n509) );
  NAND2_X1 U448 ( .A1(n172), .A2(n179), .ZN(n510) );
  NAND3_X1 U449 ( .A1(n508), .A2(n509), .A3(n510), .ZN(n165) );
  NAND2_X1 U450 ( .A1(n177), .A2(n168), .ZN(n511) );
  NAND2_X1 U451 ( .A1(n177), .A2(n166), .ZN(n512) );
  NAND2_X1 U452 ( .A1(n168), .A2(n166), .ZN(n513) );
  NAND3_X1 U453 ( .A1(n511), .A2(n512), .A3(n513), .ZN(n163) );
  OR3_X2 U454 ( .A1(n514), .A2(n515), .A3(n516), .ZN(n191) );
  AND2_X1 U455 ( .A1(n253), .A2(n283), .ZN(n514) );
  AND2_X1 U456 ( .A1(n253), .A2(n305), .ZN(n515) );
  AND2_X1 U457 ( .A1(n305), .A2(n283), .ZN(n516) );
  INV_X1 U458 ( .A(n605), .ZN(n517) );
  XOR2_X1 U459 ( .A(n256), .B(n299), .Z(n518) );
  XOR2_X1 U460 ( .A(n230), .B(n518), .Z(n228) );
  NAND2_X1 U461 ( .A1(n230), .A2(n256), .ZN(n519) );
  NAND2_X1 U462 ( .A1(n230), .A2(n299), .ZN(n520) );
  NAND2_X1 U463 ( .A1(n256), .A2(n299), .ZN(n521) );
  NAND3_X1 U464 ( .A1(n519), .A2(n520), .A3(n521), .ZN(n227) );
  XNOR2_X1 U465 ( .A(n502), .B(n522), .ZN(product[10]) );
  NAND2_X1 U466 ( .A1(n128), .A2(n86), .ZN(n522) );
  INV_X1 U467 ( .A(n617), .ZN(n523) );
  XNOR2_X1 U468 ( .A(n525), .B(n198), .ZN(n196) );
  XNOR2_X1 U469 ( .A(n205), .B(n200), .ZN(n525) );
  XNOR2_X1 U470 ( .A(n622), .B(a[8]), .ZN(n429) );
  XNOR2_X1 U471 ( .A(n526), .B(n202), .ZN(n198) );
  XNOR2_X1 U472 ( .A(n207), .B(n209), .ZN(n526) );
  INV_X2 U473 ( .A(n626), .ZN(n625) );
  CLKBUF_X1 U474 ( .A(n254), .Z(n546) );
  OR2_X1 U475 ( .A1(n176), .A2(n185), .ZN(n527) );
  OAI21_X1 U476 ( .B1(n105), .B2(n503), .A(n106), .ZN(n528) );
  AOI21_X1 U477 ( .B1(n598), .B2(n528), .A(n491), .ZN(n529) );
  OAI21_X1 U478 ( .B1(n529), .B2(n97), .A(n98), .ZN(n530) );
  INV_X1 U479 ( .A(n544), .ZN(n37) );
  CLKBUF_X1 U480 ( .A(n529), .Z(n531) );
  INV_X1 U481 ( .A(n620), .ZN(n532) );
  INV_X1 U482 ( .A(n620), .ZN(n533) );
  INV_X1 U483 ( .A(n624), .ZN(n534) );
  INV_X1 U484 ( .A(n624), .ZN(n535) );
  XNOR2_X1 U485 ( .A(n188), .B(n536), .ZN(n186) );
  XNOR2_X1 U486 ( .A(n197), .B(n190), .ZN(n536) );
  INV_X1 U487 ( .A(n614), .ZN(n537) );
  CLKBUF_X1 U488 ( .A(n18), .Z(n538) );
  BUF_X1 U489 ( .A(n18), .Z(n539) );
  BUF_X1 U490 ( .A(n18), .Z(n540) );
  NAND2_X1 U491 ( .A1(n429), .A2(n27), .ZN(n541) );
  INV_X1 U492 ( .A(n612), .ZN(n542) );
  NAND2_X1 U493 ( .A1(n593), .A2(n490), .ZN(n18) );
  AOI21_X1 U494 ( .B1(n530), .B2(n595), .A(n93), .ZN(n543) );
  XNOR2_X1 U495 ( .A(n624), .B(a[12]), .ZN(n544) );
  INV_X1 U496 ( .A(n624), .ZN(n623) );
  AOI21_X1 U497 ( .B1(n558), .B2(n80), .A(n81), .ZN(n545) );
  XOR2_X1 U498 ( .A(n253), .B(n283), .Z(n547) );
  XOR2_X1 U499 ( .A(n547), .B(n305), .Z(n192) );
  XOR2_X1 U500 ( .A(n193), .B(n282), .Z(n548) );
  XOR2_X1 U501 ( .A(n548), .B(n191), .Z(n180) );
  NAND2_X1 U502 ( .A1(n193), .A2(n282), .ZN(n549) );
  NAND2_X1 U503 ( .A1(n193), .A2(n191), .ZN(n550) );
  NAND2_X1 U504 ( .A1(n282), .A2(n191), .ZN(n551) );
  NAND3_X1 U505 ( .A1(n549), .A2(n550), .A3(n551), .ZN(n179) );
  OR2_X2 U506 ( .A1(n552), .A2(n591), .ZN(n34) );
  INV_X1 U507 ( .A(n591), .ZN(n32) );
  OR2_X2 U508 ( .A1(n553), .A2(n592), .ZN(n23) );
  XNOR2_X1 U509 ( .A(n19), .B(a[6]), .ZN(n553) );
  XOR2_X1 U510 ( .A(n613), .B(a[2]), .Z(n9) );
  XNOR2_X1 U511 ( .A(n619), .B(a[4]), .ZN(n593) );
  XNOR2_X1 U512 ( .A(n149), .B(n554), .ZN(n144) );
  XNOR2_X1 U513 ( .A(n271), .B(n146), .ZN(n554) );
  INV_X1 U514 ( .A(n619), .ZN(n617) );
  NAND2_X1 U515 ( .A1(n188), .A2(n197), .ZN(n555) );
  NAND2_X1 U516 ( .A1(n188), .A2(n190), .ZN(n556) );
  NAND2_X1 U517 ( .A1(n197), .A2(n190), .ZN(n557) );
  NAND3_X1 U518 ( .A1(n555), .A2(n556), .A3(n557), .ZN(n185) );
  OAI21_X1 U519 ( .B1(n543), .B2(n89), .A(n90), .ZN(n558) );
  NOR2_X1 U520 ( .A1(n196), .A2(n203), .ZN(n85) );
  NAND2_X1 U521 ( .A1(n429), .A2(n27), .ZN(n29) );
  INV_X2 U522 ( .A(n567), .ZN(n27) );
  XNOR2_X1 U523 ( .A(n546), .B(n559), .ZN(n208) );
  XNOR2_X1 U524 ( .A(n295), .B(n285), .ZN(n559) );
  XNOR2_X1 U525 ( .A(n206), .B(n560), .ZN(n204) );
  XNOR2_X1 U526 ( .A(n208), .B(n213), .ZN(n560) );
  NAND2_X1 U527 ( .A1(n207), .A2(n209), .ZN(n561) );
  NAND2_X1 U528 ( .A1(n207), .A2(n202), .ZN(n562) );
  NAND2_X1 U529 ( .A1(n209), .A2(n202), .ZN(n563) );
  NAND3_X1 U530 ( .A1(n561), .A2(n562), .A3(n563), .ZN(n197) );
  NAND2_X1 U531 ( .A1(n205), .A2(n200), .ZN(n564) );
  NAND2_X1 U532 ( .A1(n205), .A2(n198), .ZN(n565) );
  NAND2_X1 U533 ( .A1(n200), .A2(n198), .ZN(n566) );
  NAND3_X1 U534 ( .A1(n564), .A2(n565), .A3(n566), .ZN(n195) );
  XNOR2_X1 U535 ( .A(n620), .B(a[8]), .ZN(n567) );
  CLKBUF_X1 U536 ( .A(n104), .Z(n568) );
  CLKBUF_X1 U537 ( .A(n503), .Z(n569) );
  NAND2_X1 U538 ( .A1(n254), .A2(n295), .ZN(n570) );
  NAND2_X1 U539 ( .A1(n254), .A2(n285), .ZN(n571) );
  NAND2_X1 U540 ( .A1(n295), .A2(n285), .ZN(n572) );
  NAND3_X1 U541 ( .A1(n570), .A2(n571), .A3(n572), .ZN(n207) );
  XOR2_X1 U542 ( .A(n616), .B(a[4]), .Z(n16) );
  NAND2_X1 U543 ( .A1(n206), .A2(n208), .ZN(n573) );
  NAND2_X1 U544 ( .A1(n206), .A2(n213), .ZN(n574) );
  NAND2_X1 U545 ( .A1(n208), .A2(n213), .ZN(n575) );
  NAND3_X1 U546 ( .A1(n573), .A2(n574), .A3(n575), .ZN(n203) );
  OR2_X1 U547 ( .A1(n204), .A2(n211), .ZN(n576) );
  XNOR2_X1 U548 ( .A(n616), .B(a[2]), .ZN(n432) );
  XNOR2_X1 U549 ( .A(n611), .B(n249), .ZN(n577) );
  NOR2_X1 U550 ( .A1(n186), .A2(n195), .ZN(n578) );
  NOR2_X1 U551 ( .A1(n186), .A2(n195), .ZN(n82) );
  AND2_X1 U552 ( .A1(n232), .A2(n233), .ZN(n579) );
  NAND2_X1 U553 ( .A1(n604), .A2(n432), .ZN(n580) );
  NAND2_X1 U554 ( .A1(n604), .A2(n432), .ZN(n581) );
  NAND2_X1 U555 ( .A1(n604), .A2(n432), .ZN(n12) );
  NOR2_X1 U556 ( .A1(n164), .A2(n175), .ZN(n582) );
  NOR2_X1 U557 ( .A1(n164), .A2(n175), .ZN(n75) );
  INV_X1 U558 ( .A(n592), .ZN(n21) );
  INV_X1 U559 ( .A(n616), .ZN(n583) );
  INV_X1 U560 ( .A(n616), .ZN(n614) );
  INV_X1 U561 ( .A(n249), .ZN(n610) );
  NAND2_X1 U562 ( .A1(n226), .A2(n229), .ZN(n584) );
  NAND2_X1 U563 ( .A1(n226), .A2(n298), .ZN(n585) );
  NAND2_X1 U564 ( .A1(n229), .A2(n298), .ZN(n586) );
  NAND3_X1 U565 ( .A1(n584), .A2(n585), .A3(n586), .ZN(n223) );
  INV_X1 U566 ( .A(n610), .ZN(n587) );
  INV_X2 U567 ( .A(n587), .ZN(n588) );
  CLKBUF_X1 U568 ( .A(n96), .Z(n589) );
  XNOR2_X1 U569 ( .A(n622), .B(a[10]), .ZN(n591) );
  INV_X2 U570 ( .A(n622), .ZN(n621) );
  AOI21_X1 U571 ( .B1(n558), .B2(n80), .A(n81), .ZN(n45) );
  XNOR2_X1 U572 ( .A(n619), .B(a[6]), .ZN(n592) );
  BUF_X1 U573 ( .A(n43), .Z(n608) );
  NAND2_X1 U574 ( .A1(n594), .A2(n69), .ZN(n47) );
  INV_X1 U575 ( .A(n73), .ZN(n71) );
  AOI21_X1 U576 ( .B1(n594), .B2(n74), .A(n67), .ZN(n65) );
  INV_X1 U577 ( .A(n69), .ZN(n67) );
  NAND2_X1 U578 ( .A1(n73), .A2(n594), .ZN(n64) );
  INV_X1 U579 ( .A(n74), .ZN(n72) );
  INV_X1 U580 ( .A(n95), .ZN(n93) );
  XNOR2_X1 U581 ( .A(n77), .B(n48), .ZN(product[13]) );
  NAND2_X1 U582 ( .A1(n496), .A2(n76), .ZN(n48) );
  INV_X1 U583 ( .A(n85), .ZN(n128) );
  OR2_X1 U584 ( .A1(n152), .A2(n163), .ZN(n594) );
  OAI21_X1 U585 ( .B1(n79), .B2(n75), .A(n76), .ZN(n74) );
  NOR2_X1 U586 ( .A1(n582), .A2(n78), .ZN(n73) );
  XNOR2_X1 U587 ( .A(n84), .B(n50), .ZN(product[11]) );
  NAND2_X1 U588 ( .A1(n127), .A2(n83), .ZN(n50) );
  OAI21_X1 U589 ( .B1(n87), .B2(n85), .A(n86), .ZN(n84) );
  INV_X1 U590 ( .A(n578), .ZN(n127) );
  NAND2_X1 U591 ( .A1(n152), .A2(n163), .ZN(n69) );
  NOR2_X1 U592 ( .A1(n578), .A2(n85), .ZN(n80) );
  OAI21_X1 U593 ( .B1(n82), .B2(n86), .A(n83), .ZN(n81) );
  NAND2_X1 U594 ( .A1(n595), .A2(n499), .ZN(n53) );
  NAND2_X1 U595 ( .A1(n133), .A2(n106), .ZN(n56) );
  INV_X1 U596 ( .A(n105), .ZN(n133) );
  NAND2_X1 U597 ( .A1(n493), .A2(n98), .ZN(n54) );
  NOR2_X1 U598 ( .A1(n176), .A2(n185), .ZN(n78) );
  NAND2_X1 U599 ( .A1(n598), .A2(n103), .ZN(n55) );
  NAND2_X1 U600 ( .A1(n599), .A2(n111), .ZN(n57) );
  NAND2_X1 U601 ( .A1(n186), .A2(n195), .ZN(n83) );
  AOI21_X1 U602 ( .B1(n596), .B2(n120), .A(n117), .ZN(n115) );
  INV_X1 U603 ( .A(n119), .ZN(n117) );
  NAND2_X1 U604 ( .A1(n196), .A2(n203), .ZN(n86) );
  INV_X1 U605 ( .A(n122), .ZN(n120) );
  XNOR2_X1 U606 ( .A(n59), .B(n120), .ZN(product[2]) );
  NAND2_X1 U607 ( .A1(n596), .A2(n119), .ZN(n59) );
  NAND2_X1 U608 ( .A1(n176), .A2(n185), .ZN(n79) );
  NOR2_X1 U609 ( .A1(n204), .A2(n211), .ZN(n89) );
  NAND2_X1 U610 ( .A1(n164), .A2(n175), .ZN(n76) );
  NAND2_X1 U611 ( .A1(n204), .A2(n211), .ZN(n90) );
  NAND2_X1 U612 ( .A1(n212), .A2(n217), .ZN(n95) );
  OR2_X1 U613 ( .A1(n212), .A2(n217), .ZN(n595) );
  NAND2_X1 U614 ( .A1(n328), .A2(n314), .ZN(n119) );
  XNOR2_X1 U615 ( .A(n63), .B(n46), .ZN(product[15]) );
  NAND2_X1 U616 ( .A1(n597), .A2(n62), .ZN(n46) );
  OR2_X1 U617 ( .A1(n328), .A2(n314), .ZN(n596) );
  OR2_X1 U618 ( .A1(n151), .A2(n139), .ZN(n597) );
  NOR2_X1 U619 ( .A1(n228), .A2(n231), .ZN(n105) );
  NOR2_X1 U620 ( .A1(n234), .A2(n257), .ZN(n113) );
  NAND2_X1 U621 ( .A1(n218), .A2(n223), .ZN(n98) );
  NAND2_X1 U622 ( .A1(n228), .A2(n231), .ZN(n106) );
  OR2_X1 U623 ( .A1(n224), .A2(n227), .ZN(n598) );
  OR2_X1 U624 ( .A1(n232), .A2(n233), .ZN(n599) );
  NAND2_X1 U625 ( .A1(n224), .A2(n227), .ZN(n103) );
  NAND2_X1 U626 ( .A1(n232), .A2(n233), .ZN(n111) );
  AND2_X1 U627 ( .A1(n497), .A2(n122), .ZN(product[1]) );
  OR2_X1 U628 ( .A1(n608), .A2(n537), .ZN(n392) );
  AND2_X1 U629 ( .A1(n609), .A2(n592), .ZN(n288) );
  AND2_X1 U630 ( .A1(n609), .A2(n567), .ZN(n278) );
  OR2_X1 U631 ( .A1(n608), .A2(n523), .ZN(n377) );
  XNOR2_X1 U632 ( .A(n621), .B(n608), .ZN(n352) );
  OAI22_X1 U633 ( .A1(n42), .A2(n628), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U634 ( .A1(n608), .A2(n628), .ZN(n332) );
  XNOR2_X1 U635 ( .A(n623), .B(n608), .ZN(n343) );
  XOR2_X1 U636 ( .A(n315), .B(n261), .Z(n150) );
  XNOR2_X1 U637 ( .A(n155), .B(n601), .ZN(n139) );
  XNOR2_X1 U638 ( .A(n153), .B(n141), .ZN(n601) );
  XNOR2_X1 U639 ( .A(n157), .B(n602), .ZN(n141) );
  XNOR2_X1 U640 ( .A(n145), .B(n143), .ZN(n602) );
  AND2_X1 U641 ( .A1(n245), .A2(n609), .ZN(n300) );
  XNOR2_X1 U642 ( .A(n625), .B(n608), .ZN(n336) );
  AND2_X1 U643 ( .A1(n609), .A2(n517), .ZN(n314) );
  NAND2_X1 U644 ( .A1(n427), .A2(n37), .ZN(n39) );
  XOR2_X1 U645 ( .A(n625), .B(a[12]), .Z(n427) );
  XNOR2_X1 U646 ( .A(n618), .B(n608), .ZN(n376) );
  OAI22_X1 U647 ( .A1(n505), .A2(n336), .B1(n37), .B2(n335), .ZN(n263) );
  AND2_X1 U648 ( .A1(n609), .A2(n544), .ZN(n264) );
  AND2_X1 U649 ( .A1(n609), .A2(n591), .ZN(n270) );
  AND2_X1 U650 ( .A1(n609), .A2(n506), .ZN(n260) );
  OAI22_X1 U651 ( .A1(n505), .A2(n335), .B1(n37), .B2(n334), .ZN(n262) );
  INV_X1 U652 ( .A(n19), .ZN(n620) );
  INV_X1 U653 ( .A(n25), .ZN(n622) );
  NAND2_X1 U654 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U655 ( .A(n627), .B(a[14]), .Z(n426) );
  INV_X1 U656 ( .A(n7), .ZN(n616) );
  XNOR2_X1 U657 ( .A(n533), .B(n608), .ZN(n363) );
  OAI22_X1 U658 ( .A1(n39), .A2(n626), .B1(n337), .B2(n37), .ZN(n252) );
  OR2_X1 U659 ( .A1(n608), .A2(n626), .ZN(n337) );
  AND2_X1 U660 ( .A1(n609), .A2(n249), .ZN(product[0]) );
  OR2_X1 U661 ( .A1(n608), .A2(n504), .ZN(n344) );
  OR2_X1 U662 ( .A1(n608), .A2(n620), .ZN(n364) );
  OR2_X1 U663 ( .A1(n608), .A2(n622), .ZN(n353) );
  XNOR2_X1 U664 ( .A(n533), .B(b[9]), .ZN(n354) );
  OAI22_X1 U665 ( .A1(n505), .A2(n334), .B1(n37), .B2(n333), .ZN(n261) );
  XNOR2_X1 U666 ( .A(n625), .B(n422), .ZN(n333) );
  XNOR2_X1 U667 ( .A(n618), .B(b[11]), .ZN(n365) );
  XNOR2_X1 U668 ( .A(n625), .B(n424), .ZN(n335) );
  XNOR2_X1 U669 ( .A(n625), .B(n423), .ZN(n334) );
  OAI22_X1 U670 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U671 ( .A(n627), .B(n424), .ZN(n330) );
  XNOR2_X1 U672 ( .A(n627), .B(n608), .ZN(n331) );
  XNOR2_X1 U673 ( .A(n621), .B(n418), .ZN(n345) );
  XNOR2_X1 U674 ( .A(n623), .B(n420), .ZN(n338) );
  XNOR2_X1 U675 ( .A(n615), .B(b[13]), .ZN(n378) );
  XNOR2_X1 U676 ( .A(n621), .B(n424), .ZN(n351) );
  XNOR2_X1 U677 ( .A(n534), .B(n424), .ZN(n342) );
  XNOR2_X1 U678 ( .A(n533), .B(n424), .ZN(n362) );
  XNOR2_X1 U679 ( .A(n535), .B(n423), .ZN(n341) );
  XNOR2_X1 U680 ( .A(n534), .B(n422), .ZN(n340) );
  XNOR2_X1 U681 ( .A(n535), .B(n421), .ZN(n339) );
  XNOR2_X1 U682 ( .A(n615), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U683 ( .A(n615), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U684 ( .A(n615), .B(n418), .ZN(n384) );
  XNOR2_X1 U685 ( .A(n615), .B(n419), .ZN(n385) );
  XNOR2_X1 U686 ( .A(n615), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U687 ( .A(n615), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U688 ( .A(n615), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U689 ( .A(n532), .B(n423), .ZN(n361) );
  XNOR2_X1 U690 ( .A(n621), .B(n423), .ZN(n350) );
  XNOR2_X1 U691 ( .A(n533), .B(n422), .ZN(n360) );
  XNOR2_X1 U692 ( .A(n621), .B(n422), .ZN(n349) );
  XNOR2_X1 U693 ( .A(n618), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U694 ( .A(n618), .B(n418), .ZN(n369) );
  XNOR2_X1 U695 ( .A(n618), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U696 ( .A(n618), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U697 ( .A(n532), .B(n421), .ZN(n359) );
  XNOR2_X1 U698 ( .A(n621), .B(n421), .ZN(n348) );
  XNOR2_X1 U699 ( .A(n532), .B(n420), .ZN(n358) );
  XNOR2_X1 U700 ( .A(n621), .B(n420), .ZN(n347) );
  XNOR2_X1 U701 ( .A(n533), .B(n418), .ZN(n356) );
  XNOR2_X1 U702 ( .A(n532), .B(n419), .ZN(n357) );
  XNOR2_X1 U703 ( .A(n621), .B(n419), .ZN(n346) );
  XNOR2_X1 U704 ( .A(n612), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U705 ( .A(n532), .B(b[8]), .ZN(n355) );
  XNOR2_X1 U706 ( .A(n612), .B(b[11]), .ZN(n397) );
  XNOR2_X1 U707 ( .A(n607), .B(b[13]), .ZN(n395) );
  XNOR2_X1 U708 ( .A(n607), .B(b[14]), .ZN(n394) );
  BUF_X1 U709 ( .A(n43), .Z(n609) );
  XNOR2_X1 U710 ( .A(n606), .B(b[15]), .ZN(n393) );
  OAI22_X1 U711 ( .A1(n524), .A2(n395), .B1(n394), .B2(n588), .ZN(n316) );
  OAI22_X1 U712 ( .A1(n524), .A2(n394), .B1(n393), .B2(n588), .ZN(n315) );
  OAI22_X1 U713 ( .A1(n6), .A2(n397), .B1(n396), .B2(n588), .ZN(n318) );
  OAI22_X1 U714 ( .A1(n524), .A2(n396), .B1(n395), .B2(n588), .ZN(n317) );
  OAI22_X1 U715 ( .A1(n6), .A2(n402), .B1(n401), .B2(n588), .ZN(n323) );
  OAI22_X1 U716 ( .A1(n524), .A2(n398), .B1(n397), .B2(n588), .ZN(n319) );
  OAI22_X1 U717 ( .A1(n524), .A2(n401), .B1(n400), .B2(n588), .ZN(n322) );
  OAI22_X1 U718 ( .A1(n524), .A2(n406), .B1(n405), .B2(n588), .ZN(n327) );
  OAI22_X1 U719 ( .A1(n524), .A2(n399), .B1(n398), .B2(n588), .ZN(n320) );
  OAI22_X1 U720 ( .A1(n524), .A2(n400), .B1(n399), .B2(n588), .ZN(n321) );
  OAI22_X1 U721 ( .A1(n524), .A2(n405), .B1(n404), .B2(n588), .ZN(n326) );
  OAI22_X1 U722 ( .A1(n6), .A2(n408), .B1(n407), .B2(n588), .ZN(n329) );
  OAI22_X1 U723 ( .A1(n524), .A2(n403), .B1(n402), .B2(n588), .ZN(n324) );
  OAI22_X1 U724 ( .A1(n6), .A2(n407), .B1(n406), .B2(n588), .ZN(n328) );
  OAI22_X1 U725 ( .A1(n6), .A2(n404), .B1(n403), .B2(n588), .ZN(n325) );
  INV_X1 U726 ( .A(n13), .ZN(n619) );
  OAI21_X1 U727 ( .B1(n105), .B2(n107), .A(n106), .ZN(n104) );
  OAI22_X1 U728 ( .A1(n541), .A2(n346), .B1(n345), .B2(n27), .ZN(n271) );
  OAI22_X1 U729 ( .A1(n541), .A2(n347), .B1(n346), .B2(n27), .ZN(n272) );
  OAI22_X1 U730 ( .A1(n541), .A2(n350), .B1(n349), .B2(n27), .ZN(n275) );
  OAI22_X1 U731 ( .A1(n29), .A2(n348), .B1(n347), .B2(n27), .ZN(n273) );
  OAI22_X1 U732 ( .A1(n541), .A2(n352), .B1(n351), .B2(n27), .ZN(n277) );
  OAI22_X1 U733 ( .A1(n29), .A2(n349), .B1(n348), .B2(n27), .ZN(n274) );
  OAI22_X1 U734 ( .A1(n541), .A2(n351), .B1(n350), .B2(n27), .ZN(n276) );
  OAI22_X1 U735 ( .A1(n29), .A2(n622), .B1(n353), .B2(n27), .ZN(n254) );
  AOI21_X1 U736 ( .B1(n598), .B2(n104), .A(n491), .ZN(n99) );
  OAI21_X1 U737 ( .B1(n113), .B2(n115), .A(n114), .ZN(n112) );
  XNOR2_X1 U738 ( .A(n589), .B(n53), .ZN(product[8]) );
  OAI21_X1 U739 ( .B1(n99), .B2(n97), .A(n98), .ZN(n96) );
  AOI21_X1 U740 ( .B1(n599), .B2(n112), .A(n579), .ZN(n107) );
  XNOR2_X1 U741 ( .A(n57), .B(n494), .ZN(product[4]) );
  OAI22_X1 U742 ( .A1(n34), .A2(n339), .B1(n338), .B2(n32), .ZN(n265) );
  OAI22_X1 U743 ( .A1(n34), .A2(n340), .B1(n339), .B2(n32), .ZN(n266) );
  OAI22_X1 U744 ( .A1(n34), .A2(n342), .B1(n341), .B2(n32), .ZN(n268) );
  OAI22_X1 U745 ( .A1(n34), .A2(n341), .B1(n340), .B2(n32), .ZN(n267) );
  OAI22_X1 U746 ( .A1(n34), .A2(n343), .B1(n342), .B2(n32), .ZN(n269) );
  OAI22_X1 U747 ( .A1(n34), .A2(n504), .B1(n344), .B2(n32), .ZN(n253) );
  NAND2_X1 U748 ( .A1(n151), .A2(n139), .ZN(n62) );
  INV_X1 U749 ( .A(n613), .ZN(n606) );
  INV_X1 U750 ( .A(n613), .ZN(n607) );
  INV_X1 U751 ( .A(n613), .ZN(n611) );
  INV_X1 U752 ( .A(n1), .ZN(n613) );
  INV_X1 U753 ( .A(n113), .ZN(n135) );
  OR2_X1 U754 ( .A1(n608), .A2(n542), .ZN(n409) );
  INV_X1 U755 ( .A(n613), .ZN(n612) );
  XOR2_X1 U756 ( .A(n58), .B(n115), .Z(product[3]) );
  NAND2_X1 U757 ( .A1(n135), .A2(n114), .ZN(n58) );
  OAI21_X1 U758 ( .B1(n91), .B2(n89), .A(n90), .ZN(n88) );
  INV_X1 U759 ( .A(n88), .ZN(n87) );
  XNOR2_X1 U760 ( .A(n70), .B(n47), .ZN(product[14]) );
  XOR2_X1 U761 ( .A(n54), .B(n531), .Z(product[7]) );
  OAI22_X1 U762 ( .A1(n23), .A2(n358), .B1(n21), .B2(n357), .ZN(n282) );
  OAI22_X1 U763 ( .A1(n23), .A2(n356), .B1(n355), .B2(n21), .ZN(n280) );
  OAI22_X1 U764 ( .A1(n23), .A2(n360), .B1(n21), .B2(n359), .ZN(n284) );
  OAI22_X1 U765 ( .A1(n23), .A2(n357), .B1(n356), .B2(n21), .ZN(n281) );
  OAI22_X1 U766 ( .A1(n23), .A2(n362), .B1(n361), .B2(n21), .ZN(n286) );
  OAI22_X1 U767 ( .A1(n23), .A2(n361), .B1(n360), .B2(n21), .ZN(n285) );
  OAI22_X1 U768 ( .A1(n23), .A2(n355), .B1(n354), .B2(n21), .ZN(n279) );
  OAI22_X1 U769 ( .A1(n23), .A2(n620), .B1(n364), .B2(n21), .ZN(n255) );
  OAI22_X1 U770 ( .A1(n23), .A2(n359), .B1(n21), .B2(n358), .ZN(n283) );
  OAI22_X1 U771 ( .A1(n23), .A2(n363), .B1(n362), .B2(n21), .ZN(n287) );
  XNOR2_X1 U772 ( .A(n617), .B(n419), .ZN(n370) );
  XNOR2_X1 U773 ( .A(n617), .B(n420), .ZN(n371) );
  XNOR2_X1 U774 ( .A(n617), .B(n424), .ZN(n375) );
  XNOR2_X1 U775 ( .A(n617), .B(n421), .ZN(n372) );
  XNOR2_X1 U776 ( .A(n617), .B(n423), .ZN(n374) );
  XNOR2_X1 U777 ( .A(n617), .B(n422), .ZN(n373) );
  XNOR2_X1 U778 ( .A(n612), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U779 ( .A(n606), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U780 ( .A(n606), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U781 ( .A(n606), .B(n418), .ZN(n401) );
  XNOR2_X1 U782 ( .A(n606), .B(n608), .ZN(n408) );
  XNOR2_X1 U783 ( .A(n612), .B(n419), .ZN(n402) );
  XNOR2_X1 U784 ( .A(n607), .B(n420), .ZN(n403) );
  XNOR2_X1 U785 ( .A(n607), .B(n422), .ZN(n405) );
  XNOR2_X1 U786 ( .A(n606), .B(n424), .ZN(n407) );
  XNOR2_X1 U787 ( .A(n612), .B(n423), .ZN(n406) );
  XNOR2_X1 U788 ( .A(n607), .B(n421), .ZN(n404) );
  OAI21_X1 U789 ( .B1(n64), .B2(n45), .A(n65), .ZN(n63) );
  OAI21_X1 U790 ( .B1(n545), .B2(n78), .A(n79), .ZN(n77) );
  XNOR2_X1 U791 ( .A(n568), .B(n55), .ZN(product[6]) );
  OAI22_X1 U792 ( .A1(n539), .A2(n370), .B1(n369), .B2(n603), .ZN(n293) );
  OAI22_X1 U793 ( .A1(n540), .A2(n367), .B1(n366), .B2(n603), .ZN(n290) );
  OAI22_X1 U794 ( .A1(n539), .A2(n375), .B1(n374), .B2(n603), .ZN(n298) );
  OAI22_X1 U795 ( .A1(n540), .A2(n368), .B1(n367), .B2(n603), .ZN(n291) );
  OAI22_X1 U796 ( .A1(n539), .A2(n373), .B1(n372), .B2(n603), .ZN(n296) );
  OAI22_X1 U797 ( .A1(n540), .A2(n369), .B1(n368), .B2(n603), .ZN(n292) );
  OAI22_X1 U798 ( .A1(n539), .A2(n372), .B1(n371), .B2(n603), .ZN(n295) );
  OAI22_X1 U799 ( .A1(n538), .A2(n374), .B1(n373), .B2(n603), .ZN(n297) );
  OAI22_X1 U800 ( .A1(n540), .A2(n376), .B1(n375), .B2(n603), .ZN(n299) );
  OAI22_X1 U801 ( .A1(n539), .A2(n523), .B1(n377), .B2(n603), .ZN(n256) );
  OAI22_X1 U802 ( .A1(n540), .A2(n371), .B1(n370), .B2(n603), .ZN(n294) );
  OAI22_X1 U803 ( .A1(n538), .A2(n366), .B1(n365), .B2(n603), .ZN(n289) );
  XNOR2_X1 U804 ( .A(n583), .B(n420), .ZN(n386) );
  INV_X1 U805 ( .A(n603), .ZN(n245) );
  XNOR2_X1 U806 ( .A(n583), .B(n608), .ZN(n391) );
  XNOR2_X1 U807 ( .A(n614), .B(n422), .ZN(n388) );
  XNOR2_X1 U808 ( .A(n583), .B(n421), .ZN(n387) );
  XNOR2_X1 U809 ( .A(n583), .B(n424), .ZN(n390) );
  XNOR2_X1 U810 ( .A(n614), .B(n423), .ZN(n389) );
  OAI21_X1 U811 ( .B1(n71), .B2(n545), .A(n72), .ZN(n70) );
  XOR2_X1 U812 ( .A(n56), .B(n569), .Z(product[5]) );
  NAND2_X1 U813 ( .A1(n329), .A2(n258), .ZN(n122) );
  AOI21_X1 U814 ( .B1(n96), .B2(n595), .A(n93), .ZN(n91) );
  OAI22_X1 U815 ( .A1(n524), .A2(n542), .B1(n409), .B2(n588), .ZN(n258) );
  OAI22_X1 U816 ( .A1(n580), .A2(n379), .B1(n378), .B2(n605), .ZN(n301) );
  OAI22_X1 U817 ( .A1(n581), .A2(n380), .B1(n379), .B2(n605), .ZN(n302) );
  OAI22_X1 U818 ( .A1(n580), .A2(n385), .B1(n384), .B2(n605), .ZN(n307) );
  OAI22_X1 U819 ( .A1(n12), .A2(n382), .B1(n381), .B2(n605), .ZN(n304) );
  OAI22_X1 U820 ( .A1(n580), .A2(n381), .B1(n380), .B2(n605), .ZN(n303) );
  NAND2_X1 U821 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U822 ( .A1(n580), .A2(n383), .B1(n382), .B2(n605), .ZN(n305) );
  OAI22_X1 U823 ( .A1(n12), .A2(n384), .B1(n383), .B2(n605), .ZN(n306) );
  OAI22_X1 U824 ( .A1(n581), .A2(n386), .B1(n385), .B2(n605), .ZN(n308) );
  OAI22_X1 U825 ( .A1(n12), .A2(n387), .B1(n386), .B2(n605), .ZN(n309) );
  OAI22_X1 U826 ( .A1(n581), .A2(n537), .B1(n392), .B2(n605), .ZN(n257) );
  OAI22_X1 U827 ( .A1(n581), .A2(n389), .B1(n605), .B2(n388), .ZN(n311) );
  OAI22_X1 U828 ( .A1(n580), .A2(n388), .B1(n387), .B2(n605), .ZN(n310) );
  OAI22_X1 U829 ( .A1(n12), .A2(n390), .B1(n389), .B2(n605), .ZN(n312) );
  OAI22_X1 U830 ( .A1(n581), .A2(n391), .B1(n390), .B2(n605), .ZN(n313) );
  INV_X1 U831 ( .A(n616), .ZN(n615) );
  INV_X1 U832 ( .A(n619), .ZN(n618) );
  INV_X1 U833 ( .A(n31), .ZN(n624) );
  INV_X1 U834 ( .A(n36), .ZN(n626) );
  INV_X1 U835 ( .A(n628), .ZN(n627) );
  INV_X1 U836 ( .A(n40), .ZN(n628) );
  XOR2_X1 U837 ( .A(n259), .B(n251), .Z(n148) );
  XOR2_X1 U838 ( .A(n289), .B(n279), .Z(n146) );
  XOR2_X1 U839 ( .A(n159), .B(n150), .Z(n142) );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_7_DW01_add_2 ( A, B, CI, 
        SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n8, n9, n10, n11, n12, n13, n14, n15, n16, n18, n20,
         n22, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n42, n44, n45, n47, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n65, n67, n68, n69, n70,
         n71, n73, n75, n76, n77, n78, n79, n81, n83, n84, n86, n88, n89, n91,
         n94, n95, n96, n98, n100, n157, n158, n159, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175;

  XNOR2_X1 U122 ( .A(n45), .B(n157), .ZN(SUM[10]) );
  AND2_X1 U123 ( .A1(n174), .A2(n44), .ZN(n157) );
  INV_X1 U124 ( .A(n91), .ZN(n158) );
  XNOR2_X1 U125 ( .A(n37), .B(n159), .ZN(SUM[11]) );
  AND2_X1 U126 ( .A1(n91), .A2(n36), .ZN(n159) );
  AND2_X1 U127 ( .A1(n168), .A2(n86), .ZN(SUM[0]) );
  CLKBUF_X1 U128 ( .A(n55), .Z(n161) );
  NOR2_X1 U129 ( .A1(A[12]), .A2(B[12]), .ZN(n162) );
  OR2_X1 U130 ( .A1(n18), .A2(n173), .ZN(n2) );
  NOR2_X1 U131 ( .A1(A[8]), .A2(B[8]), .ZN(n163) );
  NOR2_X1 U132 ( .A1(A[14]), .A2(B[14]), .ZN(n164) );
  OR2_X1 U133 ( .A1(A[12]), .A2(B[12]), .ZN(n165) );
  AOI21_X1 U134 ( .B1(n38), .B2(n30), .A(n31), .ZN(n166) );
  AOI21_X1 U135 ( .B1(n38), .B2(n30), .A(n31), .ZN(n167) );
  INV_X1 U136 ( .A(n24), .ZN(n22) );
  OR2_X1 U137 ( .A1(A[0]), .A2(B[0]), .ZN(n168) );
  INV_X1 U138 ( .A(n60), .ZN(n59) );
  INV_X1 U139 ( .A(n51), .ZN(n50) );
  AOI21_X1 U140 ( .B1(n171), .B2(n68), .A(n65), .ZN(n63) );
  INV_X1 U141 ( .A(n67), .ZN(n65) );
  AOI21_X1 U142 ( .B1(n172), .B2(n84), .A(n81), .ZN(n79) );
  INV_X1 U143 ( .A(n83), .ZN(n81) );
  AOI21_X1 U144 ( .B1(n170), .B2(n76), .A(n73), .ZN(n71) );
  INV_X1 U145 ( .A(n75), .ZN(n73) );
  OAI21_X1 U146 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  OR2_X1 U147 ( .A1(n25), .A2(n28), .ZN(n169) );
  OAI21_X1 U148 ( .B1(n79), .B2(n77), .A(n78), .ZN(n76) );
  AOI21_X1 U149 ( .B1(n52), .B2(n60), .A(n53), .ZN(n51) );
  AOI21_X1 U150 ( .B1(n50), .B2(n175), .A(n47), .ZN(n45) );
  INV_X1 U151 ( .A(n86), .ZN(n84) );
  OAI21_X1 U152 ( .B1(n59), .B2(n57), .A(n58), .ZN(n56) );
  INV_X1 U153 ( .A(n49), .ZN(n47) );
  NAND2_X1 U154 ( .A1(n96), .A2(n62), .ZN(n11) );
  INV_X1 U155 ( .A(n61), .ZN(n96) );
  NAND2_X1 U156 ( .A1(n94), .A2(n161), .ZN(n9) );
  INV_X1 U157 ( .A(n163), .ZN(n94) );
  INV_X1 U158 ( .A(n28), .ZN(n89) );
  NAND2_X1 U159 ( .A1(n170), .A2(n75), .ZN(n14) );
  NAND2_X1 U160 ( .A1(n95), .A2(n58), .ZN(n10) );
  INV_X1 U161 ( .A(n57), .ZN(n95) );
  NAND2_X1 U162 ( .A1(n175), .A2(n49), .ZN(n8) );
  NAND2_X1 U163 ( .A1(n100), .A2(n78), .ZN(n15) );
  INV_X1 U164 ( .A(n77), .ZN(n100) );
  NAND2_X1 U165 ( .A1(n171), .A2(n67), .ZN(n12) );
  NAND2_X1 U166 ( .A1(n172), .A2(n83), .ZN(n16) );
  NAND2_X1 U167 ( .A1(n98), .A2(n70), .ZN(n13) );
  INV_X1 U168 ( .A(n69), .ZN(n98) );
  XNOR2_X1 U169 ( .A(n12), .B(n68), .ZN(SUM[5]) );
  XNOR2_X1 U170 ( .A(n14), .B(n76), .ZN(SUM[3]) );
  XOR2_X1 U171 ( .A(n15), .B(n79), .Z(SUM[2]) );
  XNOR2_X1 U172 ( .A(n16), .B(n84), .ZN(SUM[1]) );
  NAND2_X1 U173 ( .A1(n88), .A2(n26), .ZN(n3) );
  NAND2_X1 U174 ( .A1(n165), .A2(n33), .ZN(n5) );
  NAND2_X1 U175 ( .A1(n89), .A2(n29), .ZN(n4) );
  NOR2_X1 U176 ( .A1(A[8]), .A2(B[8]), .ZN(n54) );
  NOR2_X1 U177 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  OR2_X1 U178 ( .A1(A[3]), .A2(B[3]), .ZN(n170) );
  NOR2_X1 U179 ( .A1(A[7]), .A2(B[7]), .ZN(n57) );
  NOR2_X1 U180 ( .A1(A[14]), .A2(B[14]), .ZN(n25) );
  NOR2_X1 U181 ( .A1(A[12]), .A2(B[12]), .ZN(n32) );
  NOR2_X1 U182 ( .A1(A[2]), .A2(B[2]), .ZN(n77) );
  NOR2_X1 U183 ( .A1(A[6]), .A2(B[6]), .ZN(n61) );
  NAND2_X1 U184 ( .A1(A[13]), .A2(B[13]), .ZN(n29) );
  NAND2_X1 U185 ( .A1(A[11]), .A2(B[11]), .ZN(n36) );
  OR2_X1 U186 ( .A1(A[5]), .A2(B[5]), .ZN(n171) );
  OR2_X1 U187 ( .A1(A[1]), .A2(B[1]), .ZN(n172) );
  AND2_X1 U188 ( .A1(A[15]), .A2(B[15]), .ZN(n173) );
  OR2_X1 U189 ( .A1(A[10]), .A2(B[10]), .ZN(n174) );
  NAND2_X1 U190 ( .A1(A[12]), .A2(B[12]), .ZN(n33) );
  XNOR2_X1 U191 ( .A(n56), .B(n9), .ZN(SUM[8]) );
  XNOR2_X1 U192 ( .A(n50), .B(n8), .ZN(SUM[9]) );
  NOR2_X1 U193 ( .A1(A[4]), .A2(B[4]), .ZN(n69) );
  NAND2_X1 U194 ( .A1(A[7]), .A2(B[7]), .ZN(n58) );
  NAND2_X1 U195 ( .A1(A[2]), .A2(B[2]), .ZN(n78) );
  NAND2_X1 U196 ( .A1(A[6]), .A2(B[6]), .ZN(n62) );
  OR2_X1 U197 ( .A1(A[9]), .A2(B[9]), .ZN(n175) );
  NAND2_X1 U198 ( .A1(A[9]), .A2(B[9]), .ZN(n49) );
  NAND2_X1 U199 ( .A1(A[5]), .A2(B[5]), .ZN(n67) );
  NAND2_X1 U200 ( .A1(A[1]), .A2(B[1]), .ZN(n83) );
  NAND2_X1 U201 ( .A1(A[0]), .A2(B[0]), .ZN(n86) );
  NAND2_X1 U202 ( .A1(A[4]), .A2(B[4]), .ZN(n70) );
  NAND2_X1 U203 ( .A1(A[14]), .A2(B[14]), .ZN(n26) );
  NAND2_X1 U204 ( .A1(A[8]), .A2(B[8]), .ZN(n55) );
  XOR2_X1 U205 ( .A(n59), .B(n10), .Z(SUM[7]) );
  XOR2_X1 U206 ( .A(n11), .B(n63), .Z(SUM[6]) );
  XOR2_X1 U207 ( .A(n13), .B(n71), .Z(SUM[4]) );
  OAI21_X1 U208 ( .B1(n71), .B2(n69), .A(n70), .ZN(n68) );
  NAND2_X1 U209 ( .A1(A[3]), .A2(B[3]), .ZN(n75) );
  NAND2_X1 U210 ( .A1(A[10]), .A2(B[10]), .ZN(n44) );
  INV_X1 U211 ( .A(n44), .ZN(n42) );
  NOR2_X1 U212 ( .A1(n163), .A2(n57), .ZN(n52) );
  OAI21_X1 U213 ( .B1(n54), .B2(n58), .A(n55), .ZN(n53) );
  OAI21_X1 U214 ( .B1(n32), .B2(n36), .A(n33), .ZN(n31) );
  INV_X1 U215 ( .A(n25), .ZN(n88) );
  OAI21_X1 U216 ( .B1(n164), .B2(n29), .A(n26), .ZN(n24) );
  INV_X1 U217 ( .A(n35), .ZN(n91) );
  NOR2_X1 U218 ( .A1(n162), .A2(n35), .ZN(n30) );
  NOR2_X1 U219 ( .A1(A[11]), .A2(B[11]), .ZN(n35) );
  AOI21_X1 U220 ( .B1(n174), .B2(n47), .A(n42), .ZN(n40) );
  NAND2_X1 U221 ( .A1(n174), .A2(n175), .ZN(n39) );
  OAI21_X1 U222 ( .B1(n37), .B2(n158), .A(n36), .ZN(n34) );
  XNOR2_X1 U223 ( .A(n27), .B(n3), .ZN(SUM[14]) );
  INV_X1 U224 ( .A(n38), .ZN(n37) );
  XNOR2_X1 U225 ( .A(n20), .B(n2), .ZN(SUM[15]) );
  NOR2_X1 U226 ( .A1(A[15]), .A2(B[15]), .ZN(n18) );
  XNOR2_X1 U227 ( .A(n34), .B(n5), .ZN(SUM[12]) );
  XOR2_X1 U228 ( .A(n167), .B(n4), .Z(SUM[13]) );
  OAI21_X1 U229 ( .B1(n166), .B2(n28), .A(n29), .ZN(n27) );
  OAI21_X1 U230 ( .B1(n169), .B2(n167), .A(n22), .ZN(n20) );
  OAI21_X1 U231 ( .B1(n39), .B2(n51), .A(n40), .ZN(n38) );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_7 ( clk, clear_acc, 
        data_out_x, data_out, data_out_w, data_out_b, wr_en_y, m_valid, 
        m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [4:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
         N39, N40, N41, N42, N43, N44, n1, n2, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n85, n102, n111, n112, n113, n114, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n18), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n219), .CK(clk), .Q(n21) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n220), .CK(clk), .Q(n22) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n221), .CK(clk), .Q(n23) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n222), .CK(clk), .Q(n24) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n223), .CK(clk), .Q(n25) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n224), .CK(clk), .Q(n26) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n225), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n226), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n227), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n228), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n229), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n230), .CK(clk), .Q(n34) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n231), .CK(clk), .Q(n35) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n232), .CK(clk), .Q(n36) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n233), .CK(clk), .Q(n37) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n234), .CK(clk), .Q(n38) );
  DFF_X1 \f_reg[0]  ( .D(n102), .CK(clk), .Q(f[0]), .QN(n208) );
  DFF_X1 \f_reg[1]  ( .D(n85), .CK(clk), .Q(f[1]), .QN(n209) );
  DFF_X1 \f_reg[2]  ( .D(n83), .CK(clk), .Q(f[2]), .QN(n210) );
  DFF_X1 \f_reg[7]  ( .D(n78), .CK(clk), .Q(f[7]), .QN(n211) );
  DFF_X1 \f_reg[8]  ( .D(n77), .CK(clk), .Q(f[8]), .QN(n212) );
  DFF_X1 \f_reg[9]  ( .D(n76), .CK(clk), .Q(f[9]), .QN(n213) );
  DFF_X1 \f_reg[10]  ( .D(n75), .CK(clk), .Q(n48), .QN(n214) );
  DFF_X1 \f_reg[11]  ( .D(n74), .CK(clk), .Q(n46), .QN(n215) );
  DFF_X1 \f_reg[12]  ( .D(n2), .CK(clk), .Q(n45), .QN(n216) );
  DFF_X1 \f_reg[13]  ( .D(n73), .CK(clk), .Q(n43), .QN(n217) );
  DFF_X1 \f_reg[14]  ( .D(n5), .CK(clk), .Q(n42), .QN(n218) );
  DFF_X1 \f_reg[15]  ( .D(n72), .CK(clk), .Q(f[15]), .QN(n69) );
  DFF_X1 \data_out_reg[15]  ( .D(n112), .CK(clk), .Q(data_out[15]), .QN(n191)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n113), .CK(clk), .Q(data_out[14]), .QN(n190)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n114), .CK(clk), .Q(data_out[13]), .QN(n189)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n163), .CK(clk), .Q(data_out[12]), .QN(n188)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n164), .CK(clk), .Q(data_out[11]), .QN(n187)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n165), .CK(clk), .Q(data_out[10]), .QN(n186)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n166), .CK(clk), .Q(data_out[9]), .QN(n185) );
  DFF_X1 \data_out_reg[8]  ( .D(n167), .CK(clk), .Q(data_out[8]), .QN(n184) );
  DFF_X1 \data_out_reg[7]  ( .D(n168), .CK(clk), .Q(data_out[7]), .QN(n183) );
  DFF_X1 \data_out_reg[6]  ( .D(n169), .CK(clk), .Q(data_out[6]), .QN(n182) );
  DFF_X1 \data_out_reg[5]  ( .D(n170), .CK(clk), .Q(data_out[5]), .QN(n181) );
  DFF_X1 \data_out_reg[4]  ( .D(n171), .CK(clk), .Q(data_out[4]), .QN(n180) );
  DFF_X1 \data_out_reg[3]  ( .D(n172), .CK(clk), .Q(data_out[3]), .QN(n179) );
  DFF_X1 \data_out_reg[2]  ( .D(n173), .CK(clk), .Q(data_out[2]), .QN(n178) );
  DFF_X1 \data_out_reg[1]  ( .D(n174), .CK(clk), .Q(data_out[1]), .QN(n177) );
  DFF_X1 \data_out_reg[0]  ( .D(n175), .CK(clk), .Q(data_out[0]), .QN(n176) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_7_DW_mult_tc_1 mult_2021 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_7_DW01_add_2 add_2022 ( .A({n198, 
        n197, n196, n195, n194, n193, n207, n206, n205, n204, n203, n202, n201, 
        n200, n199, n192}), .B({f[15], n42, n43, n45, n46, n48, f[9:0]}), .CI(
        1'b0), .SUM(adder) );
  DFF_X1 delay_reg ( .D(n111), .CK(clk), .Q(n6), .QN(n235) );
  DFF_X1 \f_reg[3]  ( .D(n82), .CK(clk), .Q(f[3]), .QN(n61) );
  DFF_X1 \f_reg[4]  ( .D(n81), .CK(clk), .Q(f[4]), .QN(n62) );
  DFF_X1 \f_reg[5]  ( .D(n80), .CK(clk), .Q(f[5]), .QN(n63) );
  DFF_X1 \f_reg[6]  ( .D(n79), .CK(clk), .Q(f[6]), .QN(n64) );
  AND2_X1 U3 ( .A1(clear_acc_delay), .A2(n235), .ZN(n1) );
  AND2_X1 U4 ( .A1(n41), .A2(n19), .ZN(n16) );
  MUX2_X1 U5 ( .A(n27), .B(N38), .S(n235), .Z(n207) );
  NAND3_X1 U6 ( .A1(n8), .A2(n7), .A3(n9), .ZN(n2) );
  AND2_X1 U8 ( .A1(n15), .A2(n13), .ZN(n4) );
  NAND2_X1 U9 ( .A1(n14), .A2(n4), .ZN(n72) );
  MUX2_X2 U10 ( .A(n28), .B(N37), .S(n235), .Z(n206) );
  NAND3_X1 U11 ( .A1(n11), .A2(n10), .A3(n12), .ZN(n5) );
  MUX2_X2 U12 ( .A(N43), .B(n22), .S(n6), .Z(n197) );
  MUX2_X1 U13 ( .A(N44), .B(n21), .S(n6), .Z(n198) );
  MUX2_X2 U14 ( .A(N39), .B(n26), .S(n6), .Z(n193) );
  NAND2_X1 U15 ( .A1(data_out_b[12]), .A2(n18), .ZN(n7) );
  NAND2_X1 U16 ( .A1(adder[12]), .A2(n16), .ZN(n8) );
  NAND2_X1 U17 ( .A1(n59), .A2(n45), .ZN(n9) );
  MUX2_X2 U18 ( .A(n24), .B(N41), .S(n235), .Z(n195) );
  NAND2_X1 U19 ( .A1(data_out_b[14]), .A2(n18), .ZN(n10) );
  NAND2_X1 U20 ( .A1(adder[14]), .A2(n16), .ZN(n11) );
  NAND2_X1 U21 ( .A1(n59), .A2(n42), .ZN(n12) );
  NAND2_X1 U22 ( .A1(data_out_b[15]), .A2(n18), .ZN(n13) );
  NAND2_X1 U23 ( .A1(adder[15]), .A2(n16), .ZN(n14) );
  NAND2_X1 U24 ( .A1(n59), .A2(f[15]), .ZN(n15) );
  INV_X1 U25 ( .A(n19), .ZN(n18) );
  NAND2_X1 U26 ( .A1(n111), .A2(n17), .ZN(n237) );
  INV_X1 U27 ( .A(n41), .ZN(n59) );
  INV_X1 U28 ( .A(clear_acc), .ZN(n19) );
  OAI22_X1 U29 ( .A1(n179), .A2(n237), .B1(n61), .B2(n236), .ZN(n172) );
  OAI22_X1 U30 ( .A1(n180), .A2(n237), .B1(n62), .B2(n236), .ZN(n171) );
  OAI22_X1 U31 ( .A1(n181), .A2(n237), .B1(n63), .B2(n236), .ZN(n170) );
  OAI22_X1 U32 ( .A1(n182), .A2(n237), .B1(n64), .B2(n236), .ZN(n169) );
  OAI22_X1 U33 ( .A1(n183), .A2(n237), .B1(n211), .B2(n236), .ZN(n168) );
  OAI22_X1 U34 ( .A1(n184), .A2(n237), .B1(n212), .B2(n236), .ZN(n167) );
  OAI22_X1 U35 ( .A1(n185), .A2(n237), .B1(n213), .B2(n236), .ZN(n166) );
  MUX2_X1 U36 ( .A(n25), .B(N40), .S(n235), .Z(n194) );
  INV_X1 U37 ( .A(wr_en_y), .ZN(n17) );
  INV_X1 U38 ( .A(m_ready), .ZN(n20) );
  NAND2_X1 U39 ( .A1(m_valid), .A2(n20), .ZN(n39) );
  OAI21_X1 U40 ( .B1(sel[4]), .B2(n71), .A(n39), .ZN(n111) );
  MUX2_X1 U41 ( .A(n21), .B(N44), .S(n1), .Z(n219) );
  MUX2_X1 U42 ( .A(n22), .B(N43), .S(n1), .Z(n220) );
  MUX2_X1 U43 ( .A(n23), .B(N42), .S(n1), .Z(n221) );
  MUX2_X1 U44 ( .A(n23), .B(N42), .S(n235), .Z(n196) );
  MUX2_X1 U45 ( .A(n24), .B(N41), .S(n1), .Z(n222) );
  MUX2_X1 U46 ( .A(n25), .B(N40), .S(n1), .Z(n223) );
  MUX2_X1 U47 ( .A(n26), .B(N39), .S(n1), .Z(n224) );
  MUX2_X1 U48 ( .A(n27), .B(N38), .S(n1), .Z(n225) );
  MUX2_X1 U49 ( .A(n28), .B(N37), .S(n1), .Z(n226) );
  MUX2_X1 U50 ( .A(n29), .B(N36), .S(n1), .Z(n227) );
  MUX2_X1 U51 ( .A(n29), .B(N36), .S(n235), .Z(n205) );
  MUX2_X1 U52 ( .A(n32), .B(N35), .S(n1), .Z(n228) );
  MUX2_X1 U53 ( .A(n32), .B(N35), .S(n235), .Z(n204) );
  MUX2_X1 U54 ( .A(n33), .B(N34), .S(n1), .Z(n229) );
  MUX2_X1 U55 ( .A(n33), .B(N34), .S(n235), .Z(n203) );
  MUX2_X1 U56 ( .A(n34), .B(N33), .S(n1), .Z(n230) );
  MUX2_X1 U57 ( .A(n34), .B(N33), .S(n235), .Z(n202) );
  MUX2_X1 U58 ( .A(n35), .B(N32), .S(n1), .Z(n231) );
  MUX2_X1 U59 ( .A(n35), .B(N32), .S(n235), .Z(n201) );
  MUX2_X1 U60 ( .A(n36), .B(N31), .S(n1), .Z(n232) );
  MUX2_X1 U61 ( .A(n36), .B(N31), .S(n235), .Z(n200) );
  MUX2_X1 U62 ( .A(n37), .B(N30), .S(n1), .Z(n233) );
  MUX2_X1 U63 ( .A(n37), .B(N30), .S(n235), .Z(n199) );
  MUX2_X1 U64 ( .A(n38), .B(N29), .S(n1), .Z(n234) );
  MUX2_X1 U65 ( .A(n38), .B(N29), .S(n235), .Z(n192) );
  INV_X1 U66 ( .A(n39), .ZN(n40) );
  OAI21_X1 U67 ( .B1(n40), .B2(n6), .A(n19), .ZN(n41) );
  AOI222_X1 U68 ( .A1(data_out_b[13]), .A2(n18), .B1(adder[13]), .B2(n16), 
        .C1(n59), .C2(n43), .ZN(n44) );
  INV_X1 U69 ( .A(n44), .ZN(n73) );
  AOI222_X1 U70 ( .A1(data_out_b[11]), .A2(n18), .B1(adder[11]), .B2(n16), 
        .C1(n59), .C2(n46), .ZN(n47) );
  INV_X1 U71 ( .A(n47), .ZN(n74) );
  AOI222_X1 U72 ( .A1(data_out_b[10]), .A2(n18), .B1(adder[10]), .B2(n16), 
        .C1(n59), .C2(n48), .ZN(n49) );
  INV_X1 U73 ( .A(n49), .ZN(n75) );
  AOI222_X1 U74 ( .A1(data_out_b[8]), .A2(n18), .B1(adder[8]), .B2(n16), .C1(
        n59), .C2(f[8]), .ZN(n50) );
  INV_X1 U75 ( .A(n50), .ZN(n77) );
  AOI222_X1 U76 ( .A1(data_out_b[7]), .A2(n18), .B1(adder[7]), .B2(n16), .C1(
        n59), .C2(f[7]), .ZN(n51) );
  INV_X1 U77 ( .A(n51), .ZN(n78) );
  AOI222_X1 U78 ( .A1(data_out_b[6]), .A2(n18), .B1(adder[6]), .B2(n16), .C1(
        n59), .C2(f[6]), .ZN(n52) );
  INV_X1 U79 ( .A(n52), .ZN(n79) );
  AOI222_X1 U80 ( .A1(data_out_b[5]), .A2(n18), .B1(adder[5]), .B2(n16), .C1(
        n59), .C2(f[5]), .ZN(n53) );
  INV_X1 U81 ( .A(n53), .ZN(n80) );
  AOI222_X1 U82 ( .A1(data_out_b[4]), .A2(n18), .B1(adder[4]), .B2(n16), .C1(
        n59), .C2(f[4]), .ZN(n54) );
  INV_X1 U83 ( .A(n54), .ZN(n81) );
  AOI222_X1 U84 ( .A1(data_out_b[3]), .A2(n18), .B1(adder[3]), .B2(n16), .C1(
        n59), .C2(f[3]), .ZN(n55) );
  INV_X1 U85 ( .A(n55), .ZN(n82) );
  AOI222_X1 U86 ( .A1(data_out_b[2]), .A2(n18), .B1(adder[2]), .B2(n16), .C1(
        n59), .C2(f[2]), .ZN(n56) );
  INV_X1 U87 ( .A(n56), .ZN(n83) );
  AOI222_X1 U88 ( .A1(data_out_b[1]), .A2(n18), .B1(adder[1]), .B2(n16), .C1(
        n59), .C2(f[1]), .ZN(n57) );
  INV_X1 U89 ( .A(n57), .ZN(n85) );
  AOI222_X1 U90 ( .A1(data_out_b[0]), .A2(n18), .B1(adder[0]), .B2(n16), .C1(
        n59), .C2(f[0]), .ZN(n58) );
  INV_X1 U91 ( .A(n58), .ZN(n102) );
  AOI222_X1 U92 ( .A1(data_out_b[9]), .A2(n18), .B1(adder[9]), .B2(n16), .C1(
        n59), .C2(f[9]), .ZN(n60) );
  INV_X1 U93 ( .A(n60), .ZN(n76) );
  NOR4_X1 U94 ( .A1(n46), .A2(n45), .A3(n43), .A4(n42), .ZN(n68) );
  NOR4_X1 U95 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n48), .ZN(n67) );
  NAND4_X1 U96 ( .A1(n64), .A2(n63), .A3(n62), .A4(n61), .ZN(n65) );
  NOR4_X1 U97 ( .A1(n65), .A2(f[0]), .A3(f[1]), .A4(f[2]), .ZN(n66) );
  NAND3_X1 U98 ( .A1(n68), .A2(n67), .A3(n66), .ZN(n70) );
  NAND3_X1 U99 ( .A1(wr_en_y), .A2(n70), .A3(n69), .ZN(n236) );
  OAI22_X1 U100 ( .A1(n176), .A2(n237), .B1(n208), .B2(n236), .ZN(n175) );
  OAI22_X1 U101 ( .A1(n177), .A2(n237), .B1(n209), .B2(n236), .ZN(n174) );
  OAI22_X1 U102 ( .A1(n178), .A2(n237), .B1(n210), .B2(n236), .ZN(n173) );
  OAI22_X1 U103 ( .A1(n186), .A2(n237), .B1(n214), .B2(n236), .ZN(n165) );
  OAI22_X1 U104 ( .A1(n187), .A2(n237), .B1(n215), .B2(n236), .ZN(n164) );
  OAI22_X1 U105 ( .A1(n188), .A2(n237), .B1(n216), .B2(n236), .ZN(n163) );
  OAI22_X1 U106 ( .A1(n189), .A2(n237), .B1(n217), .B2(n236), .ZN(n114) );
  OAI22_X1 U107 ( .A1(n190), .A2(n237), .B1(n218), .B2(n236), .ZN(n113) );
  OAI22_X1 U108 ( .A1(n191), .A2(n237), .B1(n69), .B2(n236), .ZN(n112) );
  AND4_X1 U109 ( .A1(sel[3]), .A2(sel[2]), .A3(sel[1]), .A4(sel[0]), .ZN(n71)
         );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_6_DW_mult_tc_1 ( a, b, 
        product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n9, n12, n13, n16, n18, n19, n23, n25, n27, n29, n31, n32,
         n34, n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n50, n51,
         n53, n54, n55, n56, n57, n58, n59, n62, n63, n64, n65, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n89, n90, n91, n93, n95, n96, n97, n98, n99, n103,
         n104, n105, n106, n107, n109, n111, n112, n113, n114, n115, n117,
         n119, n120, n122, n125, n127, n131, n133, n135, n139, n141, n142,
         n143, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n237, n249, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n418,
         n419, n420, n421, n422, n423, n424, n426, n427, n429, n433, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U150 ( .A(n146), .B(n271), .Z(n147) );
  XOR2_X1 U152 ( .A(n301), .B(n148), .Z(n149) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U161 ( .A(n177), .B(n168), .CI(n166), .CO(n163), .S(n164) );
  FA_X1 U162 ( .A(n170), .B(n172), .CI(n179), .CO(n165), .S(n166) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n263), .CI(n291), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n317), .B(n252), .CO(n173), .S(n174) );
  FA_X1 U167 ( .A(n180), .B(n187), .CI(n178), .CO(n175), .S(n176) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U169 ( .A(n193), .B(n282), .CI(n191), .CO(n179), .S(n180) );
  FA_X1 U170 ( .A(n268), .B(n274), .CI(n292), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U172 ( .A(n197), .B(n190), .CI(n188), .CO(n185), .S(n186) );
  FA_X1 U173 ( .A(n199), .B(n201), .CI(n192), .CO(n187), .S(n188) );
  FA_X1 U174 ( .A(n275), .B(n293), .CI(n194), .CO(n189), .S(n190) );
  FA_X1 U175 ( .A(n253), .B(n305), .CI(n283), .CO(n191), .S(n192) );
  HA_X1 U176 ( .A(n269), .B(n319), .CO(n193), .S(n194) );
  FA_X1 U177 ( .A(n205), .B(n200), .CI(n198), .CO(n195), .S(n196) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U179 ( .A(n276), .B(n294), .CI(n284), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n320), .B(n270), .CI(n306), .CO(n201), .S(n202) );
  FA_X1 U181 ( .A(n208), .B(n213), .CI(n206), .CO(n203), .S(n204) );
  FA_X1 U182 ( .A(n215), .B(n307), .CI(n210), .CO(n205), .S(n206) );
  FA_X1 U183 ( .A(n285), .B(n254), .CI(n295), .CO(n207), .S(n208) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U185 ( .A(n216), .B(n219), .CI(n214), .CO(n211), .S(n212) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n322), .B(n278), .CI(n308), .CO(n215), .S(n216) );
  FA_X1 U188 ( .A(n225), .B(n222), .CI(n220), .CO(n217), .S(n218) );
  FA_X1 U189 ( .A(n255), .B(n309), .CI(n297), .CO(n219), .S(n220) );
  HA_X1 U190 ( .A(n287), .B(n323), .CO(n221), .S(n222) );
  FA_X1 U191 ( .A(n229), .B(n298), .CI(n226), .CO(n223), .S(n224) );
  FA_X1 U192 ( .A(n310), .B(n288), .CI(n324), .CO(n225), .S(n226) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  HA_X1 U194 ( .A(n325), .B(n311), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n326), .B(n300), .CI(n312), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  OR2_X2 U414 ( .A1(n224), .A2(n227), .ZN(n548) );
  BUF_X1 U415 ( .A(n115), .Z(n490) );
  OAI21_X1 U416 ( .B1(n113), .B2(n115), .A(n114), .ZN(n491) );
  INV_X1 U417 ( .A(n496), .ZN(n41) );
  OAI21_X1 U418 ( .B1(n113), .B2(n115), .A(n114), .ZN(n112) );
  OR2_X1 U419 ( .A1(n329), .A2(n258), .ZN(n492) );
  OR2_X2 U420 ( .A1(n493), .A2(n543), .ZN(n23) );
  XOR2_X1 U421 ( .A(n567), .B(a[6]), .Z(n493) );
  INV_X1 U422 ( .A(n508), .ZN(n103) );
  NAND2_X2 U423 ( .A1(n433), .A2(n529), .ZN(n541) );
  OR2_X2 U424 ( .A1(n535), .A2(n518), .ZN(n12) );
  XNOR2_X1 U425 ( .A(n265), .B(n494), .ZN(n145) );
  XNOR2_X1 U426 ( .A(n149), .B(n147), .ZN(n494) );
  CLKBUF_X1 U427 ( .A(n107), .Z(n495) );
  AOI21_X1 U428 ( .B1(n549), .B2(n112), .A(n109), .ZN(n107) );
  XNOR2_X1 U429 ( .A(n573), .B(a[14]), .ZN(n496) );
  XNOR2_X1 U430 ( .A(n524), .B(n497), .ZN(product[9]) );
  AND2_X1 U431 ( .A1(n539), .A2(n90), .ZN(n497) );
  INV_X1 U432 ( .A(n569), .ZN(n498) );
  INV_X1 U433 ( .A(n569), .ZN(n499) );
  INV_X1 U434 ( .A(n569), .ZN(n568) );
  INV_X2 U435 ( .A(n553), .ZN(n500) );
  INV_X1 U436 ( .A(n553), .ZN(n9) );
  BUF_X1 U437 ( .A(n37), .Z(n501) );
  INV_X1 U438 ( .A(n562), .ZN(n502) );
  INV_X2 U439 ( .A(n563), .ZN(n562) );
  OR2_X2 U440 ( .A1(n503), .A2(n531), .ZN(n34) );
  XNOR2_X1 U441 ( .A(n570), .B(a[10]), .ZN(n503) );
  INV_X1 U442 ( .A(n531), .ZN(n32) );
  INV_X1 U443 ( .A(n526), .ZN(n504) );
  INV_X1 U444 ( .A(n564), .ZN(n505) );
  XOR2_X1 U445 ( .A(n568), .B(a[8]), .Z(n506) );
  NOR2_X1 U446 ( .A1(n186), .A2(n195), .ZN(n507) );
  NOR2_X1 U447 ( .A1(n186), .A2(n195), .ZN(n82) );
  AND2_X2 U448 ( .A1(n224), .A2(n227), .ZN(n508) );
  OR2_X1 U449 ( .A1(n196), .A2(n203), .ZN(n509) );
  CLKBUF_X1 U450 ( .A(n542), .Z(n510) );
  NOR2_X1 U451 ( .A1(n164), .A2(n175), .ZN(n511) );
  NOR2_X1 U452 ( .A1(n164), .A2(n175), .ZN(n75) );
  INV_X1 U453 ( .A(n559), .ZN(n512) );
  OR2_X1 U454 ( .A1(n513), .A2(n538), .ZN(n18) );
  XNOR2_X1 U455 ( .A(n565), .B(a[4]), .ZN(n513) );
  OR2_X2 U456 ( .A1(n513), .A2(n538), .ZN(n514) );
  OR2_X1 U457 ( .A1(n513), .A2(n538), .ZN(n515) );
  OR2_X1 U458 ( .A1(n176), .A2(n185), .ZN(n516) );
  INV_X1 U459 ( .A(n566), .ZN(n517) );
  XNOR2_X1 U460 ( .A(n560), .B(a[2]), .ZN(n518) );
  NAND2_X1 U461 ( .A1(n506), .A2(n27), .ZN(n519) );
  INV_X1 U462 ( .A(n543), .ZN(n520) );
  INV_X1 U463 ( .A(n571), .ZN(n521) );
  INV_X1 U464 ( .A(n571), .ZN(n522) );
  CLKBUF_X1 U465 ( .A(n27), .Z(n523) );
  AOI21_X1 U466 ( .B1(n96), .B2(n545), .A(n93), .ZN(n524) );
  AOI21_X1 U467 ( .B1(n96), .B2(n545), .A(n93), .ZN(n91) );
  INV_X1 U468 ( .A(n567), .ZN(n525) );
  INV_X1 U469 ( .A(n567), .ZN(n526) );
  INV_X1 U470 ( .A(n538), .ZN(n16) );
  INV_X1 U471 ( .A(n534), .ZN(n27) );
  AOI21_X1 U472 ( .B1(n104), .B2(n548), .A(n508), .ZN(n527) );
  AOI21_X1 U473 ( .B1(n548), .B2(n104), .A(n508), .ZN(n99) );
  XOR2_X1 U474 ( .A(n563), .B(a[2]), .Z(n535) );
  INV_X1 U475 ( .A(n563), .ZN(n561) );
  OR2_X1 U476 ( .A1(n535), .A2(n518), .ZN(n536) );
  INV_X1 U477 ( .A(n557), .ZN(n528) );
  INV_X1 U478 ( .A(n528), .ZN(n529) );
  INV_X2 U479 ( .A(n528), .ZN(n530) );
  XNOR2_X1 U480 ( .A(n569), .B(a[10]), .ZN(n531) );
  OAI21_X1 U481 ( .B1(n524), .B2(n89), .A(n90), .ZN(n532) );
  OAI21_X1 U482 ( .B1(n527), .B2(n97), .A(n98), .ZN(n533) );
  XNOR2_X1 U483 ( .A(n567), .B(a[8]), .ZN(n534) );
  OR2_X1 U484 ( .A1(n535), .A2(n518), .ZN(n537) );
  XNOR2_X1 U485 ( .A(n560), .B(n249), .ZN(n433) );
  XNOR2_X1 U486 ( .A(n563), .B(a[4]), .ZN(n538) );
  OR2_X1 U487 ( .A1(n204), .A2(n211), .ZN(n539) );
  INV_X2 U488 ( .A(n560), .ZN(n558) );
  OAI21_X1 U489 ( .B1(n91), .B2(n89), .A(n90), .ZN(n540) );
  AOI21_X1 U490 ( .B1(n80), .B2(n532), .A(n81), .ZN(n542) );
  XNOR2_X1 U491 ( .A(n566), .B(a[6]), .ZN(n543) );
  BUF_X1 U492 ( .A(n43), .Z(n555) );
  NAND2_X1 U493 ( .A1(n544), .A2(n69), .ZN(n47) );
  INV_X1 U494 ( .A(n73), .ZN(n71) );
  AOI21_X1 U495 ( .B1(n74), .B2(n544), .A(n67), .ZN(n65) );
  INV_X1 U496 ( .A(n69), .ZN(n67) );
  INV_X1 U497 ( .A(n74), .ZN(n72) );
  NAND2_X1 U498 ( .A1(n73), .A2(n544), .ZN(n64) );
  INV_X1 U499 ( .A(n95), .ZN(n93) );
  AOI21_X1 U500 ( .B1(n80), .B2(n532), .A(n81), .ZN(n45) );
  NOR2_X1 U501 ( .A1(n507), .A2(n85), .ZN(n80) );
  OAI21_X1 U502 ( .B1(n86), .B2(n82), .A(n83), .ZN(n81) );
  OR2_X1 U503 ( .A1(n152), .A2(n163), .ZN(n544) );
  OAI21_X1 U504 ( .B1(n75), .B2(n79), .A(n76), .ZN(n74) );
  NAND2_X1 U505 ( .A1(n125), .A2(n76), .ZN(n48) );
  INV_X1 U506 ( .A(n511), .ZN(n125) );
  NAND2_X1 U507 ( .A1(n127), .A2(n83), .ZN(n50) );
  INV_X1 U508 ( .A(n507), .ZN(n127) );
  NAND2_X1 U509 ( .A1(n509), .A2(n86), .ZN(n51) );
  NOR2_X1 U510 ( .A1(n511), .A2(n78), .ZN(n73) );
  NAND2_X1 U511 ( .A1(n152), .A2(n163), .ZN(n69) );
  NAND2_X1 U512 ( .A1(n545), .A2(n95), .ZN(n53) );
  INV_X1 U513 ( .A(n111), .ZN(n109) );
  NAND2_X1 U514 ( .A1(n131), .A2(n98), .ZN(n54) );
  INV_X1 U515 ( .A(n97), .ZN(n131) );
  NOR2_X1 U516 ( .A1(n176), .A2(n185), .ZN(n78) );
  NOR2_X1 U517 ( .A1(n196), .A2(n203), .ZN(n85) );
  AOI21_X1 U518 ( .B1(n546), .B2(n120), .A(n117), .ZN(n115) );
  INV_X1 U519 ( .A(n119), .ZN(n117) );
  XNOR2_X1 U520 ( .A(n55), .B(n104), .ZN(product[6]) );
  NAND2_X1 U521 ( .A1(n548), .A2(n103), .ZN(n55) );
  XNOR2_X1 U522 ( .A(n59), .B(n120), .ZN(product[2]) );
  NAND2_X1 U523 ( .A1(n546), .A2(n119), .ZN(n59) );
  XNOR2_X1 U524 ( .A(n57), .B(n491), .ZN(product[4]) );
  NAND2_X1 U525 ( .A1(n549), .A2(n111), .ZN(n57) );
  NAND2_X1 U526 ( .A1(n196), .A2(n203), .ZN(n86) );
  NAND2_X1 U527 ( .A1(n186), .A2(n195), .ZN(n83) );
  NAND2_X1 U528 ( .A1(n164), .A2(n175), .ZN(n76) );
  NAND2_X1 U529 ( .A1(n176), .A2(n185), .ZN(n79) );
  NAND2_X1 U530 ( .A1(n212), .A2(n217), .ZN(n95) );
  NAND2_X1 U531 ( .A1(n204), .A2(n211), .ZN(n90) );
  OR2_X1 U532 ( .A1(n212), .A2(n217), .ZN(n545) );
  NAND2_X1 U533 ( .A1(n133), .A2(n106), .ZN(n56) );
  INV_X1 U534 ( .A(n105), .ZN(n133) );
  NAND2_X1 U535 ( .A1(n547), .A2(n62), .ZN(n46) );
  NAND2_X1 U536 ( .A1(n328), .A2(n314), .ZN(n119) );
  OR2_X1 U537 ( .A1(n328), .A2(n314), .ZN(n546) );
  OR2_X1 U538 ( .A1(n139), .A2(n151), .ZN(n547) );
  NOR2_X1 U539 ( .A1(n228), .A2(n231), .ZN(n105) );
  NOR2_X1 U540 ( .A1(n218), .A2(n223), .ZN(n97) );
  NOR2_X1 U541 ( .A1(n234), .A2(n257), .ZN(n113) );
  NAND2_X1 U542 ( .A1(n218), .A2(n223), .ZN(n98) );
  NAND2_X1 U543 ( .A1(n228), .A2(n231), .ZN(n106) );
  INV_X1 U544 ( .A(n37), .ZN(n237) );
  OR2_X1 U545 ( .A1(n232), .A2(n233), .ZN(n549) );
  AND2_X1 U546 ( .A1(n492), .A2(n122), .ZN(product[1]) );
  XNOR2_X1 U547 ( .A(n570), .B(a[12]), .ZN(n37) );
  OR2_X1 U548 ( .A1(n555), .A2(n502), .ZN(n392) );
  INV_X1 U549 ( .A(n249), .ZN(n557) );
  XNOR2_X1 U550 ( .A(n562), .B(n555), .ZN(n391) );
  AND2_X1 U551 ( .A1(n556), .A2(n237), .ZN(n264) );
  XNOR2_X1 U552 ( .A(n565), .B(n555), .ZN(n376) );
  XNOR2_X1 U553 ( .A(n498), .B(n555), .ZN(n352) );
  OAI22_X1 U554 ( .A1(n39), .A2(n573), .B1(n337), .B2(n501), .ZN(n252) );
  OR2_X1 U555 ( .A1(n555), .A2(n573), .ZN(n337) );
  NAND2_X1 U556 ( .A1(n429), .A2(n27), .ZN(n29) );
  XOR2_X1 U557 ( .A(n568), .B(a[8]), .Z(n429) );
  OAI22_X1 U558 ( .A1(n42), .A2(n575), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U559 ( .A1(n555), .A2(n575), .ZN(n332) );
  OAI22_X1 U560 ( .A1(n34), .A2(n343), .B1(n342), .B2(n32), .ZN(n269) );
  XNOR2_X1 U561 ( .A(n521), .B(n555), .ZN(n343) );
  NAND2_X1 U562 ( .A1(n529), .A2(n433), .ZN(n6) );
  AND2_X1 U563 ( .A1(n556), .A2(n538), .ZN(n300) );
  XOR2_X1 U564 ( .A(n315), .B(n261), .Z(n150) );
  XNOR2_X1 U565 ( .A(n155), .B(n551), .ZN(n139) );
  XNOR2_X1 U566 ( .A(n153), .B(n141), .ZN(n551) );
  XNOR2_X1 U567 ( .A(n552), .B(n157), .ZN(n141) );
  XNOR2_X1 U568 ( .A(n145), .B(n143), .ZN(n552) );
  XNOR2_X1 U569 ( .A(n572), .B(n555), .ZN(n336) );
  AND2_X1 U570 ( .A1(n556), .A2(n518), .ZN(n314) );
  NAND2_X1 U571 ( .A1(n427), .A2(n37), .ZN(n39) );
  XOR2_X1 U572 ( .A(n572), .B(a[12]), .Z(n427) );
  OAI22_X1 U573 ( .A1(n34), .A2(n342), .B1(n341), .B2(n32), .ZN(n268) );
  OAI22_X1 U574 ( .A1(n34), .A2(n341), .B1(n340), .B2(n32), .ZN(n267) );
  OAI22_X1 U575 ( .A1(n39), .A2(n336), .B1(n501), .B2(n335), .ZN(n263) );
  AND2_X1 U576 ( .A1(n556), .A2(n496), .ZN(n260) );
  OAI22_X1 U577 ( .A1(n39), .A2(n335), .B1(n501), .B2(n334), .ZN(n262) );
  AND2_X1 U578 ( .A1(n556), .A2(n543), .ZN(n288) );
  AND2_X1 U579 ( .A1(n556), .A2(n531), .ZN(n270) );
  INV_X1 U580 ( .A(n19), .ZN(n567) );
  INV_X1 U581 ( .A(n25), .ZN(n569) );
  AND2_X1 U582 ( .A1(n556), .A2(n534), .ZN(n278) );
  OAI22_X1 U583 ( .A1(n34), .A2(n571), .B1(n344), .B2(n32), .ZN(n253) );
  OAI22_X1 U584 ( .A1(n34), .A2(n340), .B1(n339), .B2(n32), .ZN(n266) );
  NAND2_X1 U585 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U586 ( .A(n574), .B(a[14]), .Z(n426) );
  OR2_X1 U587 ( .A1(n555), .A2(n571), .ZN(n344) );
  AND2_X1 U588 ( .A1(n556), .A2(n249), .ZN(product[0]) );
  OR2_X1 U589 ( .A1(n555), .A2(n504), .ZN(n364) );
  OR2_X1 U590 ( .A1(n555), .A2(n569), .ZN(n353) );
  OR2_X1 U591 ( .A1(n555), .A2(n505), .ZN(n377) );
  OAI22_X1 U592 ( .A1(n39), .A2(n334), .B1(n501), .B2(n333), .ZN(n261) );
  XNOR2_X1 U593 ( .A(n572), .B(n422), .ZN(n333) );
  XNOR2_X1 U594 ( .A(n565), .B(b[11]), .ZN(n365) );
  XNOR2_X1 U595 ( .A(n522), .B(n424), .ZN(n342) );
  XNOR2_X1 U596 ( .A(n522), .B(n423), .ZN(n341) );
  XNOR2_X1 U597 ( .A(n521), .B(n422), .ZN(n340) );
  XNOR2_X1 U598 ( .A(n522), .B(n421), .ZN(n339) );
  XNOR2_X1 U599 ( .A(n572), .B(n424), .ZN(n335) );
  XNOR2_X1 U600 ( .A(n572), .B(n423), .ZN(n334) );
  OAI22_X1 U601 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U602 ( .A(n574), .B(n424), .ZN(n330) );
  XNOR2_X1 U603 ( .A(n574), .B(n555), .ZN(n331) );
  XNOR2_X1 U604 ( .A(n498), .B(n418), .ZN(n345) );
  OAI22_X1 U605 ( .A1(n34), .A2(n339), .B1(n338), .B2(n32), .ZN(n265) );
  XNOR2_X1 U606 ( .A(n521), .B(n420), .ZN(n338) );
  XNOR2_X1 U607 ( .A(n562), .B(b[13]), .ZN(n378) );
  XNOR2_X1 U608 ( .A(n561), .B(n424), .ZN(n390) );
  XNOR2_X1 U609 ( .A(n499), .B(n424), .ZN(n351) );
  XNOR2_X1 U610 ( .A(n562), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U611 ( .A(n562), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U612 ( .A(n562), .B(n418), .ZN(n384) );
  XNOR2_X1 U613 ( .A(n562), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U614 ( .A(n562), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U615 ( .A(n562), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U616 ( .A(n562), .B(n419), .ZN(n385) );
  XNOR2_X1 U617 ( .A(n561), .B(n422), .ZN(n388) );
  XNOR2_X1 U618 ( .A(n561), .B(n423), .ZN(n389) );
  XNOR2_X1 U619 ( .A(n498), .B(n423), .ZN(n350) );
  XNOR2_X1 U620 ( .A(n499), .B(n422), .ZN(n349) );
  XNOR2_X1 U621 ( .A(n517), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U622 ( .A(n564), .B(n418), .ZN(n369) );
  XNOR2_X1 U623 ( .A(n565), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U624 ( .A(n564), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U625 ( .A(n558), .B(b[11]), .ZN(n397) );
  XNOR2_X1 U626 ( .A(n558), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U627 ( .A(n558), .B(b[13]), .ZN(n395) );
  XNOR2_X1 U628 ( .A(n558), .B(b[14]), .ZN(n394) );
  XNOR2_X1 U629 ( .A(n562), .B(n420), .ZN(n386) );
  XNOR2_X1 U630 ( .A(n498), .B(n420), .ZN(n347) );
  XNOR2_X1 U631 ( .A(n561), .B(n421), .ZN(n387) );
  XNOR2_X1 U632 ( .A(n499), .B(n421), .ZN(n348) );
  XNOR2_X1 U633 ( .A(n499), .B(n419), .ZN(n346) );
  XNOR2_X1 U634 ( .A(n558), .B(b[15]), .ZN(n393) );
  BUF_X1 U635 ( .A(n43), .Z(n556) );
  XNOR2_X1 U636 ( .A(n560), .B(a[2]), .ZN(n553) );
  INV_X1 U637 ( .A(n1), .ZN(n560) );
  INV_X1 U638 ( .A(n13), .ZN(n566) );
  OAI21_X1 U639 ( .B1(n87), .B2(n85), .A(n86), .ZN(n84) );
  XNOR2_X1 U640 ( .A(n45), .B(n554), .ZN(product[12]) );
  AND2_X1 U641 ( .A1(n516), .A2(n79), .ZN(n554) );
  XNOR2_X1 U642 ( .A(n84), .B(n50), .ZN(product[11]) );
  NOR2_X1 U643 ( .A1(n204), .A2(n211), .ZN(n89) );
  OAI22_X1 U644 ( .A1(n519), .A2(n350), .B1(n349), .B2(n523), .ZN(n275) );
  OAI22_X1 U645 ( .A1(n519), .A2(n346), .B1(n345), .B2(n523), .ZN(n271) );
  OAI22_X1 U646 ( .A1(n519), .A2(n347), .B1(n346), .B2(n523), .ZN(n272) );
  OAI22_X1 U647 ( .A1(n519), .A2(n348), .B1(n347), .B2(n523), .ZN(n273) );
  OAI22_X1 U648 ( .A1(n29), .A2(n349), .B1(n348), .B2(n27), .ZN(n274) );
  OAI22_X1 U649 ( .A1(n29), .A2(n569), .B1(n353), .B2(n27), .ZN(n254) );
  OAI22_X1 U650 ( .A1(n519), .A2(n351), .B1(n350), .B2(n27), .ZN(n276) );
  XNOR2_X1 U651 ( .A(n525), .B(n419), .ZN(n357) );
  XNOR2_X1 U652 ( .A(n525), .B(n418), .ZN(n356) );
  OAI22_X1 U653 ( .A1(n29), .A2(n352), .B1(n351), .B2(n27), .ZN(n277) );
  XNOR2_X1 U654 ( .A(n525), .B(n422), .ZN(n360) );
  XNOR2_X1 U655 ( .A(n526), .B(n423), .ZN(n361) );
  XNOR2_X1 U656 ( .A(n526), .B(b[9]), .ZN(n354) );
  XNOR2_X1 U657 ( .A(n525), .B(n555), .ZN(n363) );
  XNOR2_X1 U658 ( .A(n526), .B(b[8]), .ZN(n355) );
  XNOR2_X1 U659 ( .A(n525), .B(n421), .ZN(n359) );
  XNOR2_X1 U660 ( .A(n526), .B(n424), .ZN(n362) );
  XNOR2_X1 U661 ( .A(n526), .B(n420), .ZN(n358) );
  XOR2_X1 U662 ( .A(n58), .B(n490), .Z(product[3]) );
  INV_X1 U663 ( .A(n113), .ZN(n135) );
  XNOR2_X1 U664 ( .A(n540), .B(n51), .ZN(product[10]) );
  INV_X1 U665 ( .A(n540), .ZN(n87) );
  XNOR2_X1 U666 ( .A(n517), .B(n424), .ZN(n375) );
  XNOR2_X1 U667 ( .A(n564), .B(n419), .ZN(n370) );
  XNOR2_X1 U668 ( .A(n564), .B(n420), .ZN(n371) );
  XNOR2_X1 U669 ( .A(n517), .B(n423), .ZN(n374) );
  XNOR2_X1 U670 ( .A(n565), .B(n422), .ZN(n373) );
  XNOR2_X1 U671 ( .A(n517), .B(n421), .ZN(n372) );
  XNOR2_X1 U672 ( .A(n63), .B(n46), .ZN(product[15]) );
  INV_X1 U673 ( .A(n7), .ZN(n563) );
  XNOR2_X1 U674 ( .A(n77), .B(n48), .ZN(product[13]) );
  OR2_X1 U675 ( .A1(n555), .A2(n512), .ZN(n409) );
  INV_X1 U676 ( .A(n560), .ZN(n559) );
  OAI22_X1 U677 ( .A1(n23), .A2(n356), .B1(n355), .B2(n520), .ZN(n280) );
  OAI22_X1 U678 ( .A1(n23), .A2(n358), .B1(n357), .B2(n520), .ZN(n282) );
  OAI22_X1 U679 ( .A1(n23), .A2(n362), .B1(n361), .B2(n520), .ZN(n286) );
  OAI22_X1 U680 ( .A1(n23), .A2(n360), .B1(n359), .B2(n520), .ZN(n284) );
  OAI22_X1 U681 ( .A1(n23), .A2(n504), .B1(n364), .B2(n520), .ZN(n255) );
  OAI22_X1 U682 ( .A1(n23), .A2(n361), .B1(n360), .B2(n520), .ZN(n285) );
  OAI22_X1 U683 ( .A1(n23), .A2(n355), .B1(n354), .B2(n520), .ZN(n279) );
  OAI22_X1 U684 ( .A1(n23), .A2(n357), .B1(n356), .B2(n520), .ZN(n281) );
  OAI22_X1 U685 ( .A1(n23), .A2(n363), .B1(n362), .B2(n520), .ZN(n287) );
  OAI22_X1 U686 ( .A1(n23), .A2(n359), .B1(n358), .B2(n520), .ZN(n283) );
  XOR2_X1 U687 ( .A(n56), .B(n495), .Z(product[5]) );
  OAI21_X1 U688 ( .B1(n105), .B2(n107), .A(n106), .ZN(n104) );
  NAND2_X1 U689 ( .A1(n232), .A2(n233), .ZN(n111) );
  XNOR2_X1 U690 ( .A(n558), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U691 ( .A(n559), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U692 ( .A(n558), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U693 ( .A(n558), .B(n418), .ZN(n401) );
  XNOR2_X1 U694 ( .A(n559), .B(n419), .ZN(n402) );
  XNOR2_X1 U695 ( .A(n559), .B(n420), .ZN(n403) );
  XNOR2_X1 U696 ( .A(n558), .B(n555), .ZN(n408) );
  XNOR2_X1 U697 ( .A(n559), .B(n422), .ZN(n405) );
  XNOR2_X1 U698 ( .A(n559), .B(n421), .ZN(n404) );
  XNOR2_X1 U699 ( .A(n558), .B(n424), .ZN(n407) );
  XNOR2_X1 U700 ( .A(n558), .B(n423), .ZN(n406) );
  NAND2_X1 U701 ( .A1(n151), .A2(n139), .ZN(n62) );
  OAI22_X1 U702 ( .A1(n515), .A2(n370), .B1(n369), .B2(n16), .ZN(n293) );
  OAI22_X1 U703 ( .A1(n514), .A2(n367), .B1(n366), .B2(n16), .ZN(n290) );
  OAI22_X1 U704 ( .A1(n514), .A2(n375), .B1(n374), .B2(n16), .ZN(n298) );
  OAI22_X1 U705 ( .A1(n18), .A2(n372), .B1(n371), .B2(n16), .ZN(n295) );
  OAI22_X1 U706 ( .A1(n515), .A2(n368), .B1(n367), .B2(n16), .ZN(n291) );
  OAI22_X1 U707 ( .A1(n18), .A2(n374), .B1(n373), .B2(n16), .ZN(n297) );
  OAI22_X1 U708 ( .A1(n515), .A2(n369), .B1(n368), .B2(n16), .ZN(n292) );
  OAI22_X1 U709 ( .A1(n514), .A2(n373), .B1(n372), .B2(n16), .ZN(n296) );
  OAI22_X1 U710 ( .A1(n18), .A2(n371), .B1(n370), .B2(n16), .ZN(n294) );
  OAI22_X1 U711 ( .A1(n515), .A2(n376), .B1(n375), .B2(n16), .ZN(n299) );
  OAI22_X1 U712 ( .A1(n514), .A2(n505), .B1(n377), .B2(n16), .ZN(n256) );
  OAI22_X1 U713 ( .A1(n514), .A2(n366), .B1(n365), .B2(n16), .ZN(n289) );
  NAND2_X1 U714 ( .A1(n135), .A2(n114), .ZN(n58) );
  OAI21_X1 U715 ( .B1(n71), .B2(n45), .A(n72), .ZN(n70) );
  OAI21_X1 U716 ( .B1(n542), .B2(n78), .A(n79), .ZN(n77) );
  XNOR2_X1 U717 ( .A(n70), .B(n47), .ZN(product[14]) );
  OAI21_X1 U718 ( .B1(n64), .B2(n510), .A(n65), .ZN(n63) );
  XNOR2_X1 U719 ( .A(n533), .B(n53), .ZN(product[8]) );
  OAI22_X1 U720 ( .A1(n6), .A2(n395), .B1(n394), .B2(n530), .ZN(n316) );
  OAI22_X1 U721 ( .A1(n541), .A2(n394), .B1(n393), .B2(n530), .ZN(n315) );
  OAI22_X1 U722 ( .A1(n541), .A2(n396), .B1(n395), .B2(n530), .ZN(n317) );
  OAI22_X1 U723 ( .A1(n541), .A2(n397), .B1(n396), .B2(n530), .ZN(n318) );
  OAI22_X1 U724 ( .A1(n398), .A2(n6), .B1(n397), .B2(n530), .ZN(n319) );
  OAI22_X1 U725 ( .A1(n541), .A2(n400), .B1(n399), .B2(n530), .ZN(n321) );
  OAI22_X1 U726 ( .A1(n401), .A2(n6), .B1(n400), .B2(n530), .ZN(n322) );
  OAI22_X1 U727 ( .A1(n541), .A2(n399), .B1(n398), .B2(n530), .ZN(n320) );
  OAI22_X1 U728 ( .A1(n402), .A2(n6), .B1(n401), .B2(n530), .ZN(n323) );
  OAI22_X1 U729 ( .A1(n541), .A2(n404), .B1(n403), .B2(n530), .ZN(n325) );
  OAI22_X1 U730 ( .A1(n6), .A2(n403), .B1(n402), .B2(n530), .ZN(n324) );
  OAI22_X1 U731 ( .A1(n541), .A2(n406), .B1(n405), .B2(n530), .ZN(n327) );
  OAI22_X1 U732 ( .A1(n541), .A2(n405), .B1(n404), .B2(n530), .ZN(n326) );
  OAI22_X1 U733 ( .A1(n541), .A2(n407), .B1(n406), .B2(n530), .ZN(n328) );
  OAI22_X1 U734 ( .A1(n541), .A2(n408), .B1(n407), .B2(n530), .ZN(n329) );
  INV_X1 U735 ( .A(n122), .ZN(n120) );
  NAND2_X1 U736 ( .A1(n329), .A2(n258), .ZN(n122) );
  OAI21_X1 U737 ( .B1(n99), .B2(n97), .A(n98), .ZN(n96) );
  OAI22_X1 U738 ( .A1(n6), .A2(n512), .B1(n409), .B2(n530), .ZN(n258) );
  XOR2_X1 U739 ( .A(n527), .B(n54), .Z(product[7]) );
  OAI22_X1 U740 ( .A1(n537), .A2(n379), .B1(n378), .B2(n500), .ZN(n301) );
  OAI22_X1 U741 ( .A1(n536), .A2(n380), .B1(n379), .B2(n500), .ZN(n302) );
  OAI22_X1 U742 ( .A1(n536), .A2(n385), .B1(n384), .B2(n500), .ZN(n307) );
  OAI22_X1 U743 ( .A1(n537), .A2(n382), .B1(n381), .B2(n500), .ZN(n304) );
  OAI22_X1 U744 ( .A1(n536), .A2(n381), .B1(n380), .B2(n500), .ZN(n303) );
  NAND2_X1 U745 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U746 ( .A1(n537), .A2(n383), .B1(n382), .B2(n500), .ZN(n305) );
  OAI22_X1 U747 ( .A1(n536), .A2(n384), .B1(n383), .B2(n500), .ZN(n306) );
  OAI22_X1 U748 ( .A1(n536), .A2(n386), .B1(n385), .B2(n500), .ZN(n308) );
  OAI22_X1 U749 ( .A1(n537), .A2(n387), .B1(n386), .B2(n500), .ZN(n309) );
  OAI22_X1 U750 ( .A1(n537), .A2(n502), .B1(n392), .B2(n500), .ZN(n257) );
  OAI22_X1 U751 ( .A1(n12), .A2(n389), .B1(n388), .B2(n9), .ZN(n311) );
  OAI22_X1 U752 ( .A1(n12), .A2(n388), .B1(n387), .B2(n9), .ZN(n310) );
  OAI22_X1 U753 ( .A1(n12), .A2(n390), .B1(n389), .B2(n9), .ZN(n312) );
  OAI22_X1 U754 ( .A1(n536), .A2(n391), .B1(n390), .B2(n9), .ZN(n313) );
  INV_X1 U755 ( .A(n566), .ZN(n564) );
  INV_X1 U756 ( .A(n566), .ZN(n565) );
  INV_X1 U757 ( .A(n571), .ZN(n570) );
  INV_X1 U758 ( .A(n31), .ZN(n571) );
  INV_X1 U759 ( .A(n573), .ZN(n572) );
  INV_X1 U760 ( .A(n36), .ZN(n573) );
  INV_X1 U761 ( .A(n575), .ZN(n574) );
  INV_X1 U762 ( .A(n40), .ZN(n575) );
  XOR2_X1 U763 ( .A(n259), .B(n251), .Z(n148) );
  XOR2_X1 U764 ( .A(n289), .B(n279), .Z(n146) );
  XOR2_X1 U765 ( .A(n159), .B(n150), .Z(n142) );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_6_DW01_add_2 ( A, B, CI, 
        SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n5, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n19,
         n20, n22, n24, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n44, n45, n47, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n65, n67, n68, n69, n70, n71,
         n73, n75, n76, n77, n78, n79, n81, n83, n84, n86, n90, n94, n95, n96,
         n98, n100, n157, n158, n159, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177;

  XNOR2_X1 U122 ( .A(n164), .B(n157), .ZN(SUM[13]) );
  AND2_X1 U123 ( .A1(n174), .A2(n29), .ZN(n157) );
  OR2_X1 U124 ( .A1(A[11]), .A2(B[11]), .ZN(n158) );
  XNOR2_X1 U125 ( .A(n37), .B(n159), .ZN(SUM[11]) );
  AND2_X1 U126 ( .A1(n158), .A2(n36), .ZN(n159) );
  AND2_X1 U127 ( .A1(n165), .A2(n86), .ZN(SUM[0]) );
  OR2_X1 U128 ( .A1(A[15]), .A2(B[15]), .ZN(n161) );
  INV_X1 U129 ( .A(n158), .ZN(n162) );
  NOR2_X1 U130 ( .A1(A[11]), .A2(B[11]), .ZN(n35) );
  NOR2_X1 U131 ( .A1(A[8]), .A2(B[8]), .ZN(n163) );
  OR2_X2 U132 ( .A1(A[10]), .A2(B[10]), .ZN(n171) );
  AOI21_X1 U133 ( .B1(n38), .B2(n30), .A(n31), .ZN(n164) );
  OR2_X1 U134 ( .A1(A[0]), .A2(B[0]), .ZN(n165) );
  INV_X1 U135 ( .A(n51), .ZN(n50) );
  AOI21_X1 U136 ( .B1(n168), .B2(n76), .A(n73), .ZN(n71) );
  INV_X1 U137 ( .A(n75), .ZN(n73) );
  AOI21_X1 U138 ( .B1(n167), .B2(n84), .A(n81), .ZN(n79) );
  INV_X1 U139 ( .A(n83), .ZN(n81) );
  OAI21_X1 U140 ( .B1(n79), .B2(n77), .A(n78), .ZN(n76) );
  AOI21_X1 U141 ( .B1(n170), .B2(n68), .A(n65), .ZN(n63) );
  INV_X1 U142 ( .A(n67), .ZN(n65) );
  OAI21_X1 U143 ( .B1(n71), .B2(n69), .A(n70), .ZN(n68) );
  AOI21_X1 U144 ( .B1(n50), .B2(n166), .A(n47), .ZN(n45) );
  NAND2_X1 U145 ( .A1(n94), .A2(n55), .ZN(n9) );
  INV_X1 U146 ( .A(n86), .ZN(n84) );
  INV_X1 U147 ( .A(n173), .ZN(n44) );
  OAI21_X1 U148 ( .B1(n59), .B2(n57), .A(n58), .ZN(n56) );
  INV_X1 U149 ( .A(n49), .ZN(n47) );
  NAND2_X1 U150 ( .A1(n98), .A2(n70), .ZN(n13) );
  INV_X1 U151 ( .A(n69), .ZN(n98) );
  NAND2_X1 U152 ( .A1(n100), .A2(n78), .ZN(n15) );
  INV_X1 U153 ( .A(n77), .ZN(n100) );
  NAND2_X1 U154 ( .A1(n166), .A2(n49), .ZN(n8) );
  NAND2_X1 U155 ( .A1(n168), .A2(n75), .ZN(n14) );
  NAND2_X1 U156 ( .A1(n95), .A2(n58), .ZN(n10) );
  INV_X1 U157 ( .A(n57), .ZN(n95) );
  NAND2_X1 U158 ( .A1(n170), .A2(n67), .ZN(n12) );
  NAND2_X1 U159 ( .A1(n167), .A2(n83), .ZN(n16) );
  NAND2_X1 U160 ( .A1(n96), .A2(n62), .ZN(n11) );
  INV_X1 U161 ( .A(n61), .ZN(n96) );
  XNOR2_X1 U162 ( .A(n12), .B(n68), .ZN(SUM[5]) );
  XOR2_X1 U163 ( .A(n13), .B(n71), .Z(SUM[4]) );
  XOR2_X1 U164 ( .A(n15), .B(n79), .Z(SUM[2]) );
  AOI21_X1 U165 ( .B1(n38), .B2(n30), .A(n31), .ZN(n1) );
  NOR2_X1 U166 ( .A1(A[7]), .A2(B[7]), .ZN(n57) );
  NOR2_X1 U167 ( .A1(A[8]), .A2(B[8]), .ZN(n54) );
  OR2_X1 U168 ( .A1(A[9]), .A2(B[9]), .ZN(n166) );
  NOR2_X1 U169 ( .A1(A[2]), .A2(B[2]), .ZN(n77) );
  NOR2_X1 U170 ( .A1(A[4]), .A2(B[4]), .ZN(n69) );
  NAND2_X1 U171 ( .A1(n169), .A2(n26), .ZN(n3) );
  XOR2_X1 U172 ( .A(n45), .B(n7), .Z(SUM[10]) );
  XOR2_X1 U173 ( .A(n59), .B(n10), .Z(SUM[7]) );
  OR2_X1 U174 ( .A1(A[1]), .A2(B[1]), .ZN(n167) );
  OR2_X1 U175 ( .A1(A[3]), .A2(B[3]), .ZN(n168) );
  OR2_X1 U176 ( .A1(A[14]), .A2(B[14]), .ZN(n169) );
  NAND2_X1 U177 ( .A1(A[14]), .A2(B[14]), .ZN(n26) );
  XNOR2_X1 U178 ( .A(n14), .B(n76), .ZN(SUM[3]) );
  XNOR2_X1 U179 ( .A(n16), .B(n84), .ZN(SUM[1]) );
  NOR2_X1 U180 ( .A1(A[6]), .A2(B[6]), .ZN(n61) );
  NAND2_X1 U181 ( .A1(A[7]), .A2(B[7]), .ZN(n58) );
  OR2_X1 U182 ( .A1(A[5]), .A2(B[5]), .ZN(n170) );
  NAND2_X1 U183 ( .A1(A[2]), .A2(B[2]), .ZN(n78) );
  NAND2_X1 U184 ( .A1(A[4]), .A2(B[4]), .ZN(n70) );
  NAND2_X1 U185 ( .A1(A[5]), .A2(B[5]), .ZN(n67) );
  NAND2_X1 U186 ( .A1(A[1]), .A2(B[1]), .ZN(n83) );
  NAND2_X1 U187 ( .A1(A[0]), .A2(B[0]), .ZN(n86) );
  NAND2_X1 U188 ( .A1(A[13]), .A2(B[13]), .ZN(n29) );
  NAND2_X1 U189 ( .A1(A[6]), .A2(B[6]), .ZN(n62) );
  XNOR2_X1 U190 ( .A(n56), .B(n9), .ZN(SUM[8]) );
  XNOR2_X1 U191 ( .A(n50), .B(n8), .ZN(SUM[9]) );
  NAND2_X1 U192 ( .A1(n161), .A2(n19), .ZN(n2) );
  NAND2_X1 U193 ( .A1(A[15]), .A2(B[15]), .ZN(n19) );
  OR2_X1 U194 ( .A1(A[13]), .A2(B[13]), .ZN(n174) );
  NOR2_X1 U195 ( .A1(A[14]), .A2(B[14]), .ZN(n172) );
  AND2_X1 U196 ( .A1(A[10]), .A2(B[10]), .ZN(n173) );
  INV_X1 U197 ( .A(n24), .ZN(n22) );
  NOR2_X1 U198 ( .A1(A[12]), .A2(B[12]), .ZN(n175) );
  NOR2_X1 U199 ( .A1(A[12]), .A2(B[12]), .ZN(n32) );
  NAND2_X1 U200 ( .A1(n90), .A2(n33), .ZN(n5) );
  INV_X1 U201 ( .A(n175), .ZN(n90) );
  CLKBUF_X1 U202 ( .A(n36), .Z(n176) );
  NAND2_X1 U203 ( .A1(A[9]), .A2(B[9]), .ZN(n49) );
  NAND2_X1 U204 ( .A1(n169), .A2(n174), .ZN(n177) );
  NOR2_X1 U205 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  INV_X1 U206 ( .A(n60), .ZN(n59) );
  AOI21_X1 U207 ( .B1(n52), .B2(n60), .A(n53), .ZN(n51) );
  NAND2_X1 U208 ( .A1(A[3]), .A2(B[3]), .ZN(n75) );
  NAND2_X1 U209 ( .A1(A[12]), .A2(B[12]), .ZN(n33) );
  INV_X1 U210 ( .A(n163), .ZN(n94) );
  NOR2_X1 U211 ( .A1(n163), .A2(n57), .ZN(n52) );
  OAI21_X1 U212 ( .B1(n54), .B2(n58), .A(n55), .ZN(n53) );
  NAND2_X1 U213 ( .A1(A[8]), .A2(B[8]), .ZN(n55) );
  OAI21_X1 U214 ( .B1(n172), .B2(n29), .A(n26), .ZN(n24) );
  XOR2_X1 U215 ( .A(n11), .B(n63), .Z(SUM[6]) );
  OAI21_X1 U216 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  INV_X1 U217 ( .A(n38), .ZN(n37) );
  NAND2_X1 U218 ( .A1(A[11]), .A2(B[11]), .ZN(n36) );
  OAI21_X1 U219 ( .B1(n32), .B2(n36), .A(n33), .ZN(n31) );
  OAI21_X1 U220 ( .B1(n37), .B2(n162), .A(n176), .ZN(n34) );
  NOR2_X1 U221 ( .A1(n175), .A2(n35), .ZN(n30) );
  OAI21_X1 U222 ( .B1(n39), .B2(n51), .A(n40), .ZN(n38) );
  AOI21_X1 U223 ( .B1(n171), .B2(n47), .A(n173), .ZN(n40) );
  XNOR2_X1 U224 ( .A(n34), .B(n5), .ZN(SUM[12]) );
  XNOR2_X1 U225 ( .A(n20), .B(n2), .ZN(SUM[15]) );
  NAND2_X1 U226 ( .A1(n171), .A2(n44), .ZN(n7) );
  NAND2_X1 U227 ( .A1(n171), .A2(n166), .ZN(n39) );
  XNOR2_X1 U228 ( .A(n27), .B(n3), .ZN(SUM[14]) );
  OAI21_X1 U229 ( .B1(n1), .B2(n28), .A(n29), .ZN(n27) );
  OAI21_X1 U230 ( .B1(n1), .B2(n177), .A(n22), .ZN(n20) );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_6 ( clk, clear_acc, 
        data_out_x, data_out, data_out_w, data_out_b, wr_en_y, m_valid, 
        m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [4:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
         N39, N40, N41, N42, N43, N44, n1, n2, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n85, n102, n111, n112, n113, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n23), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n226), .CK(clk), .Q(n26) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n227), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n228), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n229), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n230), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n231), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n232), .CK(clk), .Q(n34) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n233), .CK(clk), .Q(n35) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n234), .CK(clk), .Q(n36) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n235), .CK(clk), .Q(n37) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n236), .CK(clk), .Q(n38) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n237), .CK(clk), .Q(n39) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n238), .CK(clk), .Q(n40) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n239), .CK(clk), .Q(n41) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n240), .CK(clk), .Q(n42) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n241), .CK(clk), .Q(n43) );
  DFF_X1 \f_reg[0]  ( .D(n112), .CK(clk), .Q(f[0]), .QN(n214) );
  DFF_X1 \f_reg[1]  ( .D(n111), .CK(clk), .Q(f[1]), .QN(n215) );
  DFF_X1 \f_reg[2]  ( .D(n102), .CK(clk), .Q(f[2]), .QN(n216) );
  DFF_X1 \f_reg[3]  ( .D(n85), .CK(clk), .Q(f[3]), .QN(n217) );
  DFF_X1 \f_reg[8]  ( .D(n79), .CK(clk), .Q(f[8]), .QN(n219) );
  DFF_X1 \f_reg[9]  ( .D(n78), .CK(clk), .Q(f[9]), .QN(n220) );
  DFF_X1 \f_reg[10]  ( .D(n77), .CK(clk), .Q(n52), .QN(n221) );
  DFF_X1 \f_reg[11]  ( .D(n76), .CK(clk), .Q(n50), .QN(n222) );
  DFF_X1 \f_reg[12]  ( .D(n4), .CK(clk), .Q(n49), .QN(n223) );
  DFF_X1 \f_reg[13]  ( .D(n18), .CK(clk), .Q(n48), .QN(n224) );
  DFF_X1 \f_reg[14]  ( .D(n9), .CK(clk), .Q(n47), .QN(n225) );
  DFF_X1 \f_reg[15]  ( .D(n75), .CK(clk), .Q(f[15]), .QN(n72) );
  DFF_X1 \data_out_reg[15]  ( .D(n166), .CK(clk), .Q(data_out[15]), .QN(n197)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n167), .CK(clk), .Q(data_out[14]), .QN(n196)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n168), .CK(clk), .Q(data_out[13]), .QN(n195)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n169), .CK(clk), .Q(data_out[12]), .QN(n194)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n170), .CK(clk), .Q(data_out[11]), .QN(n193)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n171), .CK(clk), .Q(data_out[10]), .QN(n192)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n172), .CK(clk), .Q(data_out[9]), .QN(n191) );
  DFF_X1 \data_out_reg[8]  ( .D(n173), .CK(clk), .Q(data_out[8]), .QN(n190) );
  DFF_X1 \data_out_reg[7]  ( .D(n174), .CK(clk), .Q(data_out[7]), .QN(n189) );
  DFF_X1 \data_out_reg[6]  ( .D(n175), .CK(clk), .Q(data_out[6]), .QN(n188) );
  DFF_X1 \data_out_reg[5]  ( .D(n176), .CK(clk), .Q(data_out[5]), .QN(n187) );
  DFF_X1 \data_out_reg[4]  ( .D(n177), .CK(clk), .Q(data_out[4]), .QN(n186) );
  DFF_X1 \data_out_reg[3]  ( .D(n178), .CK(clk), .Q(data_out[3]), .QN(n185) );
  DFF_X1 \data_out_reg[2]  ( .D(n179), .CK(clk), .Q(data_out[2]), .QN(n184) );
  DFF_X1 \data_out_reg[1]  ( .D(n180), .CK(clk), .Q(data_out[1]), .QN(n183) );
  DFF_X1 \data_out_reg[0]  ( .D(n181), .CK(clk), .Q(data_out[0]), .QN(n182) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_6_DW_mult_tc_1 mult_2021 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_6_DW01_add_2 add_2022 ( .A({n204, 
        n203, n202, n201, n200, n199, n213, n212, n211, n210, n209, n208, n207, 
        n206, n205, n198}), .B({f[15], n47, n48, n49, n50, n52, f[9:0]}), .CI(
        1'b0), .SUM(adder) );
  DFF_X1 delay_reg ( .D(n113), .CK(clk), .Q(n5), .QN(n242) );
  DFF_X1 \f_reg[4]  ( .D(n83), .CK(clk), .Q(f[4]), .QN(n65) );
  DFF_X1 \f_reg[5]  ( .D(n82), .CK(clk), .Q(f[5]), .QN(n66) );
  DFF_X1 \f_reg[6]  ( .D(n81), .CK(clk), .Q(f[6]), .QN(n67) );
  DFF_X1 \f_reg[7]  ( .D(n80), .CK(clk), .Q(f[7]), .QN(n218) );
  MUX2_X2 U3 ( .A(n28), .B(N42), .S(n242), .Z(n202) );
  AND2_X1 U4 ( .A1(clear_acc_delay), .A2(n242), .ZN(n1) );
  AND2_X1 U5 ( .A1(n46), .A2(n24), .ZN(n17) );
  AND2_X1 U6 ( .A1(n13), .A2(n11), .ZN(n2) );
  MUX2_X1 U8 ( .A(N39), .B(n33), .S(n5), .Z(n199) );
  MUX2_X2 U9 ( .A(n32), .B(N40), .S(n242), .Z(n200) );
  NAND3_X1 U10 ( .A1(n7), .A2(n6), .A3(n8), .ZN(n4) );
  NAND2_X1 U11 ( .A1(n12), .A2(n2), .ZN(n9) );
  MUX2_X2 U12 ( .A(n27), .B(N43), .S(n242), .Z(n203) );
  MUX2_X2 U13 ( .A(n35), .B(N37), .S(n242), .Z(n212) );
  NAND2_X1 U14 ( .A1(data_out_b[12]), .A2(n23), .ZN(n6) );
  NAND2_X1 U15 ( .A1(adder[12]), .A2(n17), .ZN(n7) );
  NAND2_X1 U16 ( .A1(n63), .A2(n49), .ZN(n8) );
  AND2_X1 U17 ( .A1(n16), .A2(n14), .ZN(n10) );
  NAND2_X1 U18 ( .A1(n15), .A2(n10), .ZN(n75) );
  MUX2_X2 U19 ( .A(n29), .B(N41), .S(n242), .Z(n201) );
  NAND2_X1 U20 ( .A1(data_out_b[14]), .A2(n23), .ZN(n11) );
  NAND2_X1 U21 ( .A1(adder[14]), .A2(n17), .ZN(n12) );
  NAND2_X1 U22 ( .A1(n63), .A2(n47), .ZN(n13) );
  NAND2_X1 U23 ( .A1(data_out_b[15]), .A2(n23), .ZN(n14) );
  NAND2_X1 U24 ( .A1(adder[15]), .A2(n17), .ZN(n15) );
  NAND2_X1 U25 ( .A1(n63), .A2(f[15]), .ZN(n16) );
  NAND2_X1 U26 ( .A1(n113), .A2(n22), .ZN(n244) );
  INV_X1 U27 ( .A(clear_acc), .ZN(n24) );
  OAI22_X1 U28 ( .A1(n185), .A2(n244), .B1(n217), .B2(n243), .ZN(n178) );
  OAI22_X1 U29 ( .A1(n186), .A2(n244), .B1(n65), .B2(n243), .ZN(n177) );
  OAI22_X1 U30 ( .A1(n187), .A2(n244), .B1(n66), .B2(n243), .ZN(n176) );
  OAI22_X1 U31 ( .A1(n188), .A2(n244), .B1(n67), .B2(n243), .ZN(n175) );
  OAI22_X1 U32 ( .A1(n189), .A2(n244), .B1(n218), .B2(n243), .ZN(n174) );
  OAI22_X1 U33 ( .A1(n190), .A2(n244), .B1(n219), .B2(n243), .ZN(n173) );
  OAI22_X1 U34 ( .A1(n191), .A2(n244), .B1(n220), .B2(n243), .ZN(n172) );
  NAND3_X1 U35 ( .A1(n20), .A2(n19), .A3(n21), .ZN(n18) );
  NAND2_X1 U36 ( .A1(data_out_b[13]), .A2(n23), .ZN(n19) );
  NAND2_X1 U37 ( .A1(adder[13]), .A2(n17), .ZN(n20) );
  NAND2_X1 U38 ( .A1(n63), .A2(n48), .ZN(n21) );
  INV_X1 U39 ( .A(n24), .ZN(n23) );
  INV_X1 U40 ( .A(n46), .ZN(n63) );
  INV_X1 U41 ( .A(wr_en_y), .ZN(n22) );
  INV_X1 U42 ( .A(m_ready), .ZN(n25) );
  NAND2_X1 U43 ( .A1(m_valid), .A2(n25), .ZN(n44) );
  OAI21_X1 U44 ( .B1(sel[4]), .B2(n74), .A(n44), .ZN(n113) );
  MUX2_X1 U45 ( .A(n26), .B(N44), .S(n1), .Z(n226) );
  MUX2_X1 U46 ( .A(n26), .B(N44), .S(n242), .Z(n204) );
  MUX2_X1 U47 ( .A(n27), .B(N43), .S(n1), .Z(n227) );
  MUX2_X1 U48 ( .A(n28), .B(N42), .S(n1), .Z(n228) );
  MUX2_X1 U49 ( .A(n29), .B(N41), .S(n1), .Z(n229) );
  MUX2_X1 U50 ( .A(n32), .B(N40), .S(n1), .Z(n230) );
  MUX2_X1 U51 ( .A(n33), .B(N39), .S(n1), .Z(n231) );
  MUX2_X1 U52 ( .A(n34), .B(N38), .S(n1), .Z(n232) );
  MUX2_X1 U53 ( .A(n34), .B(N38), .S(n242), .Z(n213) );
  MUX2_X1 U54 ( .A(n35), .B(N37), .S(n1), .Z(n233) );
  MUX2_X1 U55 ( .A(n36), .B(N36), .S(n1), .Z(n234) );
  MUX2_X1 U56 ( .A(n36), .B(N36), .S(n242), .Z(n211) );
  MUX2_X1 U57 ( .A(n37), .B(N35), .S(n1), .Z(n235) );
  MUX2_X1 U58 ( .A(n37), .B(N35), .S(n242), .Z(n210) );
  MUX2_X1 U59 ( .A(n38), .B(N34), .S(n1), .Z(n236) );
  MUX2_X1 U60 ( .A(n38), .B(N34), .S(n242), .Z(n209) );
  MUX2_X1 U61 ( .A(n39), .B(N33), .S(n1), .Z(n237) );
  MUX2_X1 U62 ( .A(n39), .B(N33), .S(n242), .Z(n208) );
  MUX2_X1 U63 ( .A(n40), .B(N32), .S(n1), .Z(n238) );
  MUX2_X1 U64 ( .A(n40), .B(N32), .S(n242), .Z(n207) );
  MUX2_X1 U65 ( .A(n41), .B(N31), .S(n1), .Z(n239) );
  MUX2_X1 U66 ( .A(n41), .B(N31), .S(n242), .Z(n206) );
  MUX2_X1 U67 ( .A(n42), .B(N30), .S(n1), .Z(n240) );
  MUX2_X1 U68 ( .A(n42), .B(N30), .S(n242), .Z(n205) );
  MUX2_X1 U69 ( .A(n43), .B(N29), .S(n1), .Z(n241) );
  MUX2_X1 U70 ( .A(n43), .B(N29), .S(n242), .Z(n198) );
  INV_X1 U71 ( .A(n44), .ZN(n45) );
  OAI21_X1 U72 ( .B1(n45), .B2(n5), .A(n24), .ZN(n46) );
  AOI222_X1 U73 ( .A1(data_out_b[11]), .A2(n23), .B1(adder[11]), .B2(n17), 
        .C1(n63), .C2(n50), .ZN(n51) );
  INV_X1 U74 ( .A(n51), .ZN(n76) );
  AOI222_X1 U75 ( .A1(data_out_b[10]), .A2(n23), .B1(adder[10]), .B2(n17), 
        .C1(n63), .C2(n52), .ZN(n53) );
  INV_X1 U76 ( .A(n53), .ZN(n77) );
  AOI222_X1 U77 ( .A1(data_out_b[8]), .A2(n23), .B1(adder[8]), .B2(n17), .C1(
        n63), .C2(f[8]), .ZN(n54) );
  INV_X1 U78 ( .A(n54), .ZN(n79) );
  AOI222_X1 U79 ( .A1(data_out_b[7]), .A2(n23), .B1(adder[7]), .B2(n17), .C1(
        n63), .C2(f[7]), .ZN(n55) );
  INV_X1 U80 ( .A(n55), .ZN(n80) );
  AOI222_X1 U81 ( .A1(data_out_b[6]), .A2(n23), .B1(adder[6]), .B2(n17), .C1(
        n63), .C2(f[6]), .ZN(n56) );
  INV_X1 U82 ( .A(n56), .ZN(n81) );
  AOI222_X1 U83 ( .A1(data_out_b[5]), .A2(n23), .B1(adder[5]), .B2(n17), .C1(
        n63), .C2(f[5]), .ZN(n57) );
  INV_X1 U84 ( .A(n57), .ZN(n82) );
  AOI222_X1 U85 ( .A1(data_out_b[4]), .A2(n23), .B1(adder[4]), .B2(n17), .C1(
        n63), .C2(f[4]), .ZN(n58) );
  INV_X1 U86 ( .A(n58), .ZN(n83) );
  AOI222_X1 U87 ( .A1(data_out_b[3]), .A2(n23), .B1(adder[3]), .B2(n17), .C1(
        n63), .C2(f[3]), .ZN(n59) );
  INV_X1 U88 ( .A(n59), .ZN(n85) );
  AOI222_X1 U89 ( .A1(data_out_b[2]), .A2(n23), .B1(adder[2]), .B2(n17), .C1(
        n63), .C2(f[2]), .ZN(n60) );
  INV_X1 U90 ( .A(n60), .ZN(n102) );
  AOI222_X1 U91 ( .A1(data_out_b[1]), .A2(n23), .B1(adder[1]), .B2(n17), .C1(
        n63), .C2(f[1]), .ZN(n61) );
  INV_X1 U92 ( .A(n61), .ZN(n111) );
  AOI222_X1 U93 ( .A1(data_out_b[0]), .A2(n23), .B1(adder[0]), .B2(n17), .C1(
        n63), .C2(f[0]), .ZN(n62) );
  INV_X1 U94 ( .A(n62), .ZN(n112) );
  AOI222_X1 U95 ( .A1(data_out_b[9]), .A2(n23), .B1(adder[9]), .B2(n17), .C1(
        n63), .C2(f[9]), .ZN(n64) );
  INV_X1 U96 ( .A(n64), .ZN(n78) );
  NOR4_X1 U97 ( .A1(n50), .A2(n49), .A3(n48), .A4(n47), .ZN(n71) );
  NOR4_X1 U98 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n52), .ZN(n70) );
  NAND4_X1 U99 ( .A1(n67), .A2(n66), .A3(n65), .A4(n217), .ZN(n68) );
  NOR4_X1 U100 ( .A1(n68), .A2(f[0]), .A3(f[1]), .A4(f[2]), .ZN(n69) );
  NAND3_X1 U101 ( .A1(n71), .A2(n70), .A3(n69), .ZN(n73) );
  NAND3_X1 U102 ( .A1(wr_en_y), .A2(n73), .A3(n72), .ZN(n243) );
  OAI22_X1 U103 ( .A1(n182), .A2(n244), .B1(n214), .B2(n243), .ZN(n181) );
  OAI22_X1 U104 ( .A1(n183), .A2(n244), .B1(n215), .B2(n243), .ZN(n180) );
  OAI22_X1 U105 ( .A1(n184), .A2(n244), .B1(n216), .B2(n243), .ZN(n179) );
  OAI22_X1 U106 ( .A1(n192), .A2(n244), .B1(n221), .B2(n243), .ZN(n171) );
  OAI22_X1 U107 ( .A1(n193), .A2(n244), .B1(n222), .B2(n243), .ZN(n170) );
  OAI22_X1 U108 ( .A1(n194), .A2(n244), .B1(n223), .B2(n243), .ZN(n169) );
  OAI22_X1 U109 ( .A1(n195), .A2(n244), .B1(n224), .B2(n243), .ZN(n168) );
  OAI22_X1 U110 ( .A1(n196), .A2(n244), .B1(n225), .B2(n243), .ZN(n167) );
  OAI22_X1 U111 ( .A1(n197), .A2(n244), .B1(n72), .B2(n243), .ZN(n166) );
  AND4_X1 U112 ( .A1(sel[3]), .A2(sel[2]), .A3(sel[1]), .A4(sel[0]), .ZN(n74)
         );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_5_DW_mult_tc_1 ( a, b, 
        product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n9, n12, n13, n16, n18, n19, n21, n23, n25, n27, n29, n31,
         n32, n34, n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n50,
         n53, n54, n55, n56, n58, n59, n62, n63, n64, n65, n67, n69, n70, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n93, n95, n96, n97, n98, n99, n103, n104,
         n105, n106, n107, n111, n112, n113, n114, n115, n117, n119, n120,
         n122, n125, n127, n135, n139, n141, n142, n143, n144, n145, n146,
         n148, n149, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n241,
         n245, n247, n249, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n418, n419, n420,
         n421, n422, n423, n424, n426, n427, n429, n431, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U148 ( .A(n265), .B(n144), .Z(n145) );
  XOR2_X1 U152 ( .A(n301), .B(n148), .Z(n149) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U162 ( .A(n170), .B(n172), .CI(n179), .CO(n165), .S(n166) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n263), .CI(n291), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n317), .B(n252), .CO(n173), .S(n174) );
  FA_X1 U167 ( .A(n180), .B(n187), .CI(n178), .CO(n175), .S(n176) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U169 ( .A(n193), .B(n282), .CI(n191), .CO(n179), .S(n180) );
  FA_X1 U170 ( .A(n268), .B(n292), .CI(n274), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U174 ( .A(n275), .B(n293), .CI(n194), .CO(n189), .S(n190) );
  FA_X1 U175 ( .A(n305), .B(n283), .CI(n253), .CO(n191), .S(n192) );
  HA_X1 U176 ( .A(n269), .B(n319), .CO(n193), .S(n194) );
  FA_X1 U177 ( .A(n205), .B(n200), .CI(n198), .CO(n195), .S(n196) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U179 ( .A(n276), .B(n294), .CI(n284), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n320), .B(n270), .CI(n306), .CO(n201), .S(n202) );
  FA_X1 U181 ( .A(n208), .B(n213), .CI(n206), .CO(n203), .S(n204) );
  FA_X1 U182 ( .A(n215), .B(n307), .CI(n210), .CO(n205), .S(n206) );
  FA_X1 U183 ( .A(n285), .B(n295), .CI(n254), .CO(n207), .S(n208) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U185 ( .A(n216), .B(n219), .CI(n214), .CO(n211), .S(n212) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n322), .B(n278), .CI(n308), .CO(n215), .S(n216) );
  FA_X1 U188 ( .A(n225), .B(n222), .CI(n220), .CO(n217), .S(n218) );
  FA_X1 U189 ( .A(n309), .B(n255), .CI(n297), .CO(n219), .S(n220) );
  HA_X1 U190 ( .A(n287), .B(n323), .CO(n221), .S(n222) );
  FA_X1 U192 ( .A(n324), .B(n288), .CI(n310), .CO(n225), .S(n226) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  HA_X1 U194 ( .A(n311), .B(n325), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n326), .B(n300), .CI(n312), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  NAND2_X1 U414 ( .A1(n431), .A2(n572), .ZN(n516) );
  BUF_X1 U415 ( .A(n573), .Z(n490) );
  BUF_X1 U416 ( .A(n16), .Z(n572) );
  BUF_X1 U417 ( .A(n12), .Z(n513) );
  BUF_X1 U418 ( .A(n12), .Z(n523) );
  BUF_X1 U419 ( .A(n12), .Z(n522) );
  OR2_X2 U420 ( .A1(n491), .A2(n541), .ZN(n34) );
  XNOR2_X1 U421 ( .A(n31), .B(a[10]), .ZN(n491) );
  BUF_X2 U422 ( .A(n582), .Z(n526) );
  BUF_X1 U423 ( .A(n582), .Z(n525) );
  BUF_X1 U424 ( .A(n574), .Z(n555) );
  BUF_X2 U425 ( .A(n574), .Z(n557) );
  BUF_X2 U426 ( .A(n574), .Z(n556) );
  INV_X2 U427 ( .A(n241), .ZN(n528) );
  NOR2_X1 U428 ( .A1(n186), .A2(n195), .ZN(n82) );
  OR2_X1 U429 ( .A1(n328), .A2(n314), .ZN(n492) );
  OR2_X1 U430 ( .A1(n329), .A2(n258), .ZN(n493) );
  OR2_X1 U431 ( .A1(n218), .A2(n223), .ZN(n494) );
  OR2_X1 U432 ( .A1(n75), .A2(n78), .ZN(n495) );
  AOI21_X1 U433 ( .B1(n104), .B2(n575), .A(n512), .ZN(n496) );
  CLKBUF_X1 U434 ( .A(n86), .Z(n497) );
  INV_X1 U435 ( .A(n527), .ZN(n37) );
  BUF_X2 U436 ( .A(n587), .Z(n498) );
  BUF_X2 U437 ( .A(n587), .Z(n499) );
  OAI21_X1 U438 ( .B1(n99), .B2(n97), .A(n98), .ZN(n500) );
  OAI21_X1 U439 ( .B1(n496), .B2(n97), .A(n98), .ZN(n96) );
  INV_X1 U440 ( .A(n559), .ZN(n501) );
  XNOR2_X1 U441 ( .A(n149), .B(n502), .ZN(n144) );
  XNOR2_X1 U442 ( .A(n271), .B(n146), .ZN(n502) );
  NAND2_X1 U443 ( .A1(n429), .A2(n27), .ZN(n29) );
  NAND2_X1 U444 ( .A1(n431), .A2(n572), .ZN(n18) );
  XOR2_X1 U445 ( .A(n588), .B(a[6]), .Z(n542) );
  CLKBUF_X1 U446 ( .A(n104), .Z(n503) );
  CLKBUF_X1 U447 ( .A(n32), .Z(n504) );
  AOI21_X1 U448 ( .B1(n500), .B2(n565), .A(n93), .ZN(n505) );
  NOR2_X1 U449 ( .A1(n196), .A2(n203), .ZN(n85) );
  OR2_X1 U450 ( .A1(n542), .A2(n559), .ZN(n537) );
  OR2_X1 U451 ( .A1(n228), .A2(n231), .ZN(n506) );
  XOR2_X1 U452 ( .A(n229), .B(n298), .Z(n507) );
  XOR2_X1 U453 ( .A(n226), .B(n507), .Z(n224) );
  NAND2_X1 U454 ( .A1(n226), .A2(n229), .ZN(n508) );
  NAND2_X1 U455 ( .A1(n226), .A2(n298), .ZN(n509) );
  NAND2_X1 U456 ( .A1(n229), .A2(n298), .ZN(n510) );
  NAND3_X1 U457 ( .A1(n508), .A2(n509), .A3(n510), .ZN(n223) );
  OR2_X2 U458 ( .A1(n543), .A2(n249), .ZN(n511) );
  OR2_X1 U459 ( .A1(n543), .A2(n249), .ZN(n6) );
  INV_X1 U460 ( .A(n588), .ZN(n587) );
  INV_X1 U461 ( .A(n512), .ZN(n103) );
  AND2_X1 U462 ( .A1(n224), .A2(n227), .ZN(n512) );
  CLKBUF_X1 U463 ( .A(n45), .Z(n514) );
  OR2_X1 U464 ( .A1(n196), .A2(n203), .ZN(n515) );
  INV_X1 U465 ( .A(n590), .ZN(n517) );
  INV_X1 U466 ( .A(n590), .ZN(n589) );
  INV_X1 U467 ( .A(n591), .ZN(n518) );
  INV_X1 U468 ( .A(n591), .ZN(n519) );
  XNOR2_X1 U469 ( .A(n166), .B(n520), .ZN(n164) );
  XNOR2_X1 U470 ( .A(n177), .B(n168), .ZN(n520) );
  OR2_X1 U471 ( .A1(n204), .A2(n211), .ZN(n521) );
  NAND2_X1 U472 ( .A1(n562), .A2(n9), .ZN(n12) );
  BUF_X2 U473 ( .A(n582), .Z(n524) );
  INV_X1 U474 ( .A(n583), .ZN(n582) );
  XNOR2_X1 U475 ( .A(n591), .B(a[12]), .ZN(n527) );
  XOR2_X1 U476 ( .A(n588), .B(a[8]), .Z(n27) );
  INV_X1 U477 ( .A(n541), .ZN(n32) );
  XNOR2_X1 U478 ( .A(n45), .B(n529), .ZN(product[12]) );
  AND2_X1 U479 ( .A1(n530), .A2(n79), .ZN(n529) );
  OR2_X1 U480 ( .A1(n176), .A2(n185), .ZN(n530) );
  OAI21_X1 U481 ( .B1(n505), .B2(n89), .A(n90), .ZN(n531) );
  CLKBUF_X1 U482 ( .A(n496), .Z(n532) );
  OAI21_X1 U483 ( .B1(n91), .B2(n89), .A(n90), .ZN(n88) );
  CLKBUF_X1 U484 ( .A(n500), .Z(n533) );
  INV_X1 U485 ( .A(n580), .ZN(n579) );
  INV_X2 U486 ( .A(n580), .ZN(n547) );
  NAND2_X1 U487 ( .A1(n166), .A2(n177), .ZN(n534) );
  NAND2_X1 U488 ( .A1(n166), .A2(n168), .ZN(n535) );
  NAND2_X1 U489 ( .A1(n177), .A2(n168), .ZN(n536) );
  NAND3_X1 U490 ( .A1(n534), .A2(n535), .A3(n536), .ZN(n163) );
  OR2_X1 U491 ( .A1(n542), .A2(n559), .ZN(n538) );
  OR2_X1 U492 ( .A1(n542), .A2(n559), .ZN(n23) );
  AND2_X1 U493 ( .A1(n232), .A2(n233), .ZN(n539) );
  OAI21_X1 U494 ( .B1(n107), .B2(n105), .A(n106), .ZN(n104) );
  CLKBUF_X1 U495 ( .A(n112), .Z(n540) );
  XNOR2_X1 U496 ( .A(n586), .B(a[4]), .ZN(n431) );
  XNOR2_X1 U497 ( .A(n590), .B(a[10]), .ZN(n541) );
  INV_X1 U498 ( .A(n559), .ZN(n21) );
  XOR2_X1 U499 ( .A(n580), .B(n249), .Z(n543) );
  INV_X1 U500 ( .A(n249), .ZN(n578) );
  NOR2_X1 U501 ( .A1(n164), .A2(n175), .ZN(n544) );
  NOR2_X1 U502 ( .A1(n164), .A2(n175), .ZN(n75) );
  OR2_X1 U503 ( .A1(n224), .A2(n227), .ZN(n575) );
  XNOR2_X1 U504 ( .A(n545), .B(n192), .ZN(n188) );
  XNOR2_X1 U505 ( .A(n199), .B(n201), .ZN(n545) );
  XNOR2_X1 U506 ( .A(n546), .B(n188), .ZN(n186) );
  XNOR2_X1 U507 ( .A(n197), .B(n190), .ZN(n546) );
  NAND2_X1 U508 ( .A1(n199), .A2(n201), .ZN(n548) );
  NAND2_X1 U509 ( .A1(n199), .A2(n192), .ZN(n549) );
  NAND2_X1 U510 ( .A1(n201), .A2(n192), .ZN(n550) );
  NAND3_X1 U511 ( .A1(n548), .A2(n549), .A3(n550), .ZN(n187) );
  NAND2_X1 U512 ( .A1(n197), .A2(n190), .ZN(n551) );
  NAND2_X1 U513 ( .A1(n197), .A2(n188), .ZN(n552) );
  NAND2_X1 U514 ( .A1(n190), .A2(n188), .ZN(n553) );
  NAND3_X1 U515 ( .A1(n551), .A2(n552), .A3(n553), .ZN(n185) );
  INV_X1 U516 ( .A(n583), .ZN(n581) );
  XOR2_X1 U517 ( .A(n580), .B(a[2]), .Z(n9) );
  CLKBUF_X1 U518 ( .A(n107), .Z(n554) );
  XNOR2_X1 U519 ( .A(n583), .B(a[2]), .ZN(n562) );
  BUF_X1 U520 ( .A(n9), .Z(n574) );
  AOI21_X1 U521 ( .B1(n531), .B2(n80), .A(n81), .ZN(n558) );
  XNOR2_X1 U522 ( .A(n586), .B(a[6]), .ZN(n559) );
  OR2_X1 U523 ( .A1(n152), .A2(n163), .ZN(n563) );
  XOR2_X1 U524 ( .A(n505), .B(n560), .Z(product[9]) );
  NAND2_X1 U525 ( .A1(n521), .A2(n90), .ZN(n560) );
  XOR2_X1 U526 ( .A(n561), .B(n540), .Z(product[4]) );
  AND2_X1 U527 ( .A1(n567), .A2(n111), .ZN(n561) );
  OR2_X1 U528 ( .A1(n212), .A2(n217), .ZN(n565) );
  AOI21_X1 U529 ( .B1(n74), .B2(n563), .A(n67), .ZN(n65) );
  INV_X1 U530 ( .A(n69), .ZN(n67) );
  NAND2_X1 U531 ( .A1(n563), .A2(n69), .ZN(n47) );
  NAND2_X1 U532 ( .A1(n73), .A2(n563), .ZN(n64) );
  INV_X1 U533 ( .A(n74), .ZN(n72) );
  AOI21_X1 U534 ( .B1(n80), .B2(n531), .A(n81), .ZN(n45) );
  NOR2_X1 U535 ( .A1(n82), .A2(n85), .ZN(n80) );
  OAI21_X1 U536 ( .B1(n86), .B2(n82), .A(n83), .ZN(n81) );
  AOI21_X1 U537 ( .B1(n96), .B2(n565), .A(n93), .ZN(n91) );
  INV_X1 U538 ( .A(n95), .ZN(n93) );
  XNOR2_X1 U539 ( .A(n87), .B(n564), .ZN(product[10]) );
  AND2_X1 U540 ( .A1(n515), .A2(n86), .ZN(n564) );
  OAI21_X1 U541 ( .B1(n544), .B2(n79), .A(n76), .ZN(n74) );
  NOR2_X1 U542 ( .A1(n75), .A2(n78), .ZN(n73) );
  XNOR2_X1 U543 ( .A(n84), .B(n50), .ZN(product[11]) );
  NAND2_X1 U544 ( .A1(n127), .A2(n83), .ZN(n50) );
  INV_X1 U545 ( .A(n82), .ZN(n127) );
  XNOR2_X1 U546 ( .A(n533), .B(n53), .ZN(product[8]) );
  NAND2_X1 U547 ( .A1(n565), .A2(n95), .ZN(n53) );
  XNOR2_X1 U548 ( .A(n77), .B(n48), .ZN(product[13]) );
  NAND2_X1 U549 ( .A1(n125), .A2(n76), .ZN(n48) );
  INV_X1 U550 ( .A(n544), .ZN(n125) );
  NAND2_X1 U551 ( .A1(n152), .A2(n163), .ZN(n69) );
  OAI21_X1 U552 ( .B1(n113), .B2(n115), .A(n114), .ZN(n112) );
  NAND2_X1 U553 ( .A1(n135), .A2(n114), .ZN(n58) );
  INV_X1 U554 ( .A(n113), .ZN(n135) );
  NAND2_X1 U555 ( .A1(n506), .A2(n106), .ZN(n56) );
  NAND2_X1 U556 ( .A1(n494), .A2(n98), .ZN(n54) );
  AOI21_X1 U557 ( .B1(n567), .B2(n112), .A(n539), .ZN(n107) );
  NOR2_X1 U558 ( .A1(n176), .A2(n185), .ZN(n78) );
  NAND2_X1 U559 ( .A1(n575), .A2(n103), .ZN(n55) );
  AOI21_X1 U560 ( .B1(n492), .B2(n120), .A(n117), .ZN(n115) );
  INV_X1 U561 ( .A(n119), .ZN(n117) );
  INV_X1 U562 ( .A(n122), .ZN(n120) );
  XNOR2_X1 U563 ( .A(n120), .B(n59), .ZN(product[2]) );
  NAND2_X1 U564 ( .A1(n492), .A2(n119), .ZN(n59) );
  NAND2_X1 U565 ( .A1(n196), .A2(n203), .ZN(n86) );
  NAND2_X1 U566 ( .A1(n176), .A2(n185), .ZN(n79) );
  NAND2_X1 U567 ( .A1(n164), .A2(n175), .ZN(n76) );
  NAND2_X1 U568 ( .A1(n186), .A2(n195), .ZN(n83) );
  NAND2_X1 U569 ( .A1(n212), .A2(n217), .ZN(n95) );
  NAND2_X1 U570 ( .A1(n204), .A2(n211), .ZN(n90) );
  NAND2_X1 U571 ( .A1(n566), .A2(n62), .ZN(n46) );
  NOR2_X1 U572 ( .A1(n218), .A2(n223), .ZN(n97) );
  OR2_X1 U573 ( .A1(n151), .A2(n139), .ZN(n566) );
  NOR2_X1 U574 ( .A1(n228), .A2(n231), .ZN(n105) );
  NAND2_X1 U575 ( .A1(n218), .A2(n223), .ZN(n98) );
  NAND2_X1 U576 ( .A1(n228), .A2(n231), .ZN(n106) );
  OR2_X1 U577 ( .A1(n232), .A2(n233), .ZN(n567) );
  INV_X1 U578 ( .A(n41), .ZN(n235) );
  AND2_X1 U579 ( .A1(n493), .A2(n122), .ZN(product[1]) );
  XNOR2_X1 U580 ( .A(n592), .B(a[14]), .ZN(n41) );
  OR2_X1 U581 ( .A1(n577), .A2(n583), .ZN(n392) );
  XNOR2_X1 U582 ( .A(n519), .B(n577), .ZN(n343) );
  AND2_X1 U583 ( .A1(n577), .A2(n541), .ZN(n270) );
  XNOR2_X1 U584 ( .A(n585), .B(n577), .ZN(n376) );
  XNOR2_X1 U585 ( .A(n517), .B(n577), .ZN(n352) );
  XNOR2_X1 U586 ( .A(n155), .B(n569), .ZN(n139) );
  XNOR2_X1 U587 ( .A(n153), .B(n141), .ZN(n569) );
  XNOR2_X1 U588 ( .A(n157), .B(n570), .ZN(n141) );
  XNOR2_X1 U589 ( .A(n145), .B(n143), .ZN(n570) );
  OAI22_X1 U590 ( .A1(n39), .A2(n593), .B1(n337), .B2(n37), .ZN(n252) );
  OR2_X1 U591 ( .A1(n577), .A2(n593), .ZN(n337) );
  OAI22_X1 U592 ( .A1(n42), .A2(n595), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U593 ( .A1(n577), .A2(n595), .ZN(n332) );
  AND2_X1 U594 ( .A1(n43), .A2(n245), .ZN(n300) );
  XOR2_X1 U595 ( .A(n589), .B(a[8]), .Z(n429) );
  XNOR2_X1 U596 ( .A(n159), .B(n571), .ZN(n142) );
  XNOR2_X1 U597 ( .A(n315), .B(n261), .ZN(n571) );
  XNOR2_X1 U598 ( .A(n592), .B(n577), .ZN(n336) );
  NAND2_X1 U599 ( .A1(n427), .A2(n37), .ZN(n39) );
  XOR2_X1 U600 ( .A(n592), .B(a[12]), .Z(n427) );
  AND2_X1 U601 ( .A1(n577), .A2(n241), .ZN(n278) );
  OAI22_X1 U602 ( .A1(n39), .A2(n336), .B1(n37), .B2(n335), .ZN(n263) );
  AND2_X1 U603 ( .A1(n43), .A2(n527), .ZN(n264) );
  AND2_X1 U604 ( .A1(n43), .A2(n559), .ZN(n288) );
  AND2_X1 U605 ( .A1(n43), .A2(n235), .ZN(n260) );
  OAI22_X1 U606 ( .A1(n39), .A2(n335), .B1(n37), .B2(n334), .ZN(n262) );
  INV_X1 U607 ( .A(n19), .ZN(n588) );
  INV_X1 U608 ( .A(n25), .ZN(n590) );
  NAND2_X1 U609 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U610 ( .A(n594), .B(a[14]), .Z(n426) );
  INV_X1 U611 ( .A(n7), .ZN(n583) );
  XNOR2_X1 U612 ( .A(n498), .B(n577), .ZN(n363) );
  AND2_X1 U613 ( .A1(n43), .A2(n247), .ZN(n314) );
  AND2_X1 U614 ( .A1(n43), .A2(n249), .ZN(product[0]) );
  OR2_X1 U615 ( .A1(n577), .A2(n586), .ZN(n377) );
  OR2_X1 U616 ( .A1(n577), .A2(n590), .ZN(n353) );
  OR2_X1 U617 ( .A1(n577), .A2(n588), .ZN(n364) );
  OR2_X1 U618 ( .A1(n577), .A2(n591), .ZN(n344) );
  XNOR2_X1 U619 ( .A(n498), .B(b[9]), .ZN(n354) );
  OAI22_X1 U620 ( .A1(n39), .A2(n334), .B1(n37), .B2(n333), .ZN(n261) );
  XNOR2_X1 U621 ( .A(n592), .B(n422), .ZN(n333) );
  XNOR2_X1 U622 ( .A(n585), .B(b[11]), .ZN(n365) );
  XNOR2_X1 U623 ( .A(n592), .B(n424), .ZN(n335) );
  XNOR2_X1 U624 ( .A(n592), .B(n423), .ZN(n334) );
  OAI22_X1 U625 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U626 ( .A(n594), .B(n424), .ZN(n330) );
  XNOR2_X1 U627 ( .A(n594), .B(n577), .ZN(n331) );
  XNOR2_X1 U628 ( .A(n517), .B(n418), .ZN(n345) );
  XNOR2_X1 U629 ( .A(n519), .B(n420), .ZN(n338) );
  XNOR2_X1 U630 ( .A(n525), .B(b[13]), .ZN(n378) );
  XNOR2_X1 U631 ( .A(n587), .B(n424), .ZN(n362) );
  XNOR2_X1 U632 ( .A(n517), .B(n424), .ZN(n351) );
  XNOR2_X1 U633 ( .A(n518), .B(n424), .ZN(n342) );
  XNOR2_X1 U634 ( .A(n519), .B(n423), .ZN(n341) );
  XNOR2_X1 U635 ( .A(n518), .B(n422), .ZN(n340) );
  XNOR2_X1 U636 ( .A(n519), .B(n421), .ZN(n339) );
  XNOR2_X1 U637 ( .A(n525), .B(n419), .ZN(n385) );
  XNOR2_X1 U638 ( .A(n526), .B(n418), .ZN(n384) );
  XNOR2_X1 U639 ( .A(n524), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U640 ( .A(n525), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U641 ( .A(n526), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U642 ( .A(n524), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U643 ( .A(n524), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U644 ( .A(n498), .B(n422), .ZN(n360) );
  XNOR2_X1 U645 ( .A(n517), .B(n422), .ZN(n349) );
  XNOR2_X1 U646 ( .A(n585), .B(n418), .ZN(n369) );
  XNOR2_X1 U647 ( .A(n585), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U648 ( .A(n585), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U649 ( .A(n585), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U650 ( .A(n499), .B(n423), .ZN(n361) );
  XNOR2_X1 U651 ( .A(n517), .B(n423), .ZN(n350) );
  XNOR2_X1 U652 ( .A(n547), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U653 ( .A(n547), .B(b[11]), .ZN(n397) );
  XNOR2_X1 U654 ( .A(n547), .B(b[13]), .ZN(n395) );
  XNOR2_X1 U655 ( .A(n547), .B(b[14]), .ZN(n394) );
  XNOR2_X1 U656 ( .A(n499), .B(n421), .ZN(n359) );
  XNOR2_X1 U657 ( .A(n517), .B(n421), .ZN(n348) );
  XNOR2_X1 U658 ( .A(n498), .B(n420), .ZN(n358) );
  XNOR2_X1 U659 ( .A(n517), .B(n420), .ZN(n347) );
  XNOR2_X1 U660 ( .A(n499), .B(n418), .ZN(n356) );
  XNOR2_X1 U661 ( .A(n498), .B(n419), .ZN(n357) );
  XNOR2_X1 U662 ( .A(n517), .B(n419), .ZN(n346) );
  XNOR2_X1 U663 ( .A(n499), .B(b[8]), .ZN(n355) );
  XNOR2_X1 U664 ( .A(n547), .B(b[15]), .ZN(n393) );
  CLKBUF_X3 U665 ( .A(n16), .Z(n573) );
  XNOR2_X1 U666 ( .A(n581), .B(a[4]), .ZN(n16) );
  NAND2_X1 U667 ( .A1(n328), .A2(n314), .ZN(n119) );
  OAI22_X1 U668 ( .A1(n34), .A2(n339), .B1(n338), .B2(n504), .ZN(n265) );
  OAI22_X1 U669 ( .A1(n34), .A2(n340), .B1(n339), .B2(n504), .ZN(n266) );
  OAI22_X1 U670 ( .A1(n34), .A2(n341), .B1(n340), .B2(n504), .ZN(n267) );
  OAI22_X1 U671 ( .A1(n34), .A2(n342), .B1(n341), .B2(n32), .ZN(n268) );
  OAI22_X1 U672 ( .A1(n34), .A2(n343), .B1(n342), .B2(n32), .ZN(n269) );
  OAI22_X1 U673 ( .A1(n34), .A2(n591), .B1(n344), .B2(n504), .ZN(n253) );
  INV_X1 U674 ( .A(n13), .ZN(n586) );
  XNOR2_X1 U675 ( .A(n503), .B(n55), .ZN(product[6]) );
  NOR2_X1 U676 ( .A1(n204), .A2(n211), .ZN(n89) );
  OAI22_X1 U677 ( .A1(n29), .A2(n346), .B1(n345), .B2(n528), .ZN(n271) );
  OAI22_X1 U678 ( .A1(n29), .A2(n350), .B1(n349), .B2(n528), .ZN(n275) );
  OAI22_X1 U679 ( .A1(n29), .A2(n347), .B1(n346), .B2(n528), .ZN(n272) );
  OAI22_X1 U680 ( .A1(n29), .A2(n348), .B1(n347), .B2(n528), .ZN(n273) );
  OAI22_X1 U681 ( .A1(n29), .A2(n349), .B1(n348), .B2(n528), .ZN(n274) );
  OAI22_X1 U682 ( .A1(n29), .A2(n351), .B1(n350), .B2(n528), .ZN(n276) );
  OAI22_X1 U683 ( .A1(n29), .A2(n590), .B1(n353), .B2(n528), .ZN(n254) );
  INV_X1 U684 ( .A(n27), .ZN(n241) );
  OAI22_X1 U685 ( .A1(n29), .A2(n352), .B1(n351), .B2(n528), .ZN(n277) );
  XNOR2_X1 U686 ( .A(n63), .B(n46), .ZN(product[15]) );
  INV_X1 U687 ( .A(n579), .ZN(n576) );
  INV_X1 U688 ( .A(n1), .ZN(n580) );
  XNOR2_X1 U689 ( .A(n584), .B(n424), .ZN(n375) );
  XNOR2_X1 U690 ( .A(n584), .B(n419), .ZN(n370) );
  XNOR2_X1 U691 ( .A(n584), .B(n420), .ZN(n371) );
  XNOR2_X1 U692 ( .A(n584), .B(n423), .ZN(n374) );
  XNOR2_X1 U693 ( .A(n584), .B(n422), .ZN(n373) );
  XNOR2_X1 U694 ( .A(n584), .B(n421), .ZN(n372) );
  OAI21_X1 U695 ( .B1(n87), .B2(n85), .A(n497), .ZN(n84) );
  OR2_X1 U696 ( .A1(n577), .A2(n576), .ZN(n409) );
  XNOR2_X1 U697 ( .A(n70), .B(n47), .ZN(product[14]) );
  INV_X1 U698 ( .A(n88), .ZN(n87) );
  NAND2_X1 U699 ( .A1(n151), .A2(n139), .ZN(n62) );
  OAI22_X1 U700 ( .A1(n537), .A2(n358), .B1(n357), .B2(n501), .ZN(n282) );
  OAI22_X1 U701 ( .A1(n538), .A2(n356), .B1(n355), .B2(n501), .ZN(n280) );
  OAI22_X1 U702 ( .A1(n538), .A2(n362), .B1(n361), .B2(n501), .ZN(n286) );
  OAI22_X1 U703 ( .A1(n538), .A2(n357), .B1(n356), .B2(n501), .ZN(n281) );
  OAI22_X1 U704 ( .A1(n538), .A2(n588), .B1(n364), .B2(n21), .ZN(n255) );
  OAI22_X1 U705 ( .A1(n537), .A2(n360), .B1(n359), .B2(n501), .ZN(n284) );
  OAI22_X1 U706 ( .A1(n537), .A2(n361), .B1(n360), .B2(n21), .ZN(n285) );
  OAI22_X1 U707 ( .A1(n23), .A2(n363), .B1(n362), .B2(n21), .ZN(n287) );
  OAI22_X1 U708 ( .A1(n23), .A2(n359), .B1(n358), .B2(n21), .ZN(n283) );
  OAI22_X1 U709 ( .A1(n537), .A2(n355), .B1(n354), .B2(n21), .ZN(n279) );
  AOI21_X1 U710 ( .B1(n104), .B2(n575), .A(n512), .ZN(n99) );
  XOR2_X1 U711 ( .A(n532), .B(n54), .Z(product[7]) );
  OAI22_X1 U712 ( .A1(n516), .A2(n370), .B1(n369), .B2(n490), .ZN(n293) );
  OAI22_X1 U713 ( .A1(n516), .A2(n367), .B1(n366), .B2(n573), .ZN(n290) );
  OAI22_X1 U714 ( .A1(n18), .A2(n372), .B1(n371), .B2(n573), .ZN(n295) );
  OAI22_X1 U715 ( .A1(n516), .A2(n368), .B1(n367), .B2(n490), .ZN(n291) );
  OAI22_X1 U716 ( .A1(n516), .A2(n371), .B1(n370), .B2(n573), .ZN(n294) );
  OAI22_X1 U717 ( .A1(n18), .A2(n369), .B1(n368), .B2(n573), .ZN(n292) );
  OAI22_X1 U718 ( .A1(n516), .A2(n373), .B1(n372), .B2(n573), .ZN(n296) );
  OAI22_X1 U719 ( .A1(n516), .A2(n375), .B1(n374), .B2(n573), .ZN(n298) );
  OAI22_X1 U720 ( .A1(n18), .A2(n374), .B1(n373), .B2(n573), .ZN(n297) );
  OAI22_X1 U721 ( .A1(n18), .A2(n366), .B1(n365), .B2(n573), .ZN(n289) );
  OAI22_X1 U722 ( .A1(n516), .A2(n586), .B1(n377), .B2(n490), .ZN(n256) );
  OAI22_X1 U723 ( .A1(n516), .A2(n376), .B1(n375), .B2(n573), .ZN(n299) );
  XNOR2_X1 U724 ( .A(n525), .B(n420), .ZN(n386) );
  XNOR2_X1 U725 ( .A(n524), .B(n577), .ZN(n391) );
  INV_X1 U726 ( .A(n573), .ZN(n245) );
  XNOR2_X1 U727 ( .A(n524), .B(n424), .ZN(n390) );
  XNOR2_X1 U728 ( .A(n526), .B(n422), .ZN(n388) );
  XNOR2_X1 U729 ( .A(n526), .B(n423), .ZN(n389) );
  XNOR2_X1 U730 ( .A(n524), .B(n421), .ZN(n387) );
  NAND2_X1 U731 ( .A1(n232), .A2(n233), .ZN(n111) );
  XNOR2_X1 U732 ( .A(n579), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U733 ( .A(n547), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U734 ( .A(n547), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U735 ( .A(n547), .B(n418), .ZN(n401) );
  XNOR2_X1 U736 ( .A(n547), .B(n577), .ZN(n408) );
  XNOR2_X1 U737 ( .A(n579), .B(n421), .ZN(n404) );
  XNOR2_X1 U738 ( .A(n547), .B(n422), .ZN(n405) );
  XNOR2_X1 U739 ( .A(n579), .B(n420), .ZN(n403) );
  XNOR2_X1 U740 ( .A(n579), .B(n419), .ZN(n402) );
  XNOR2_X1 U741 ( .A(n547), .B(n424), .ZN(n407) );
  XNOR2_X1 U742 ( .A(n547), .B(n423), .ZN(n406) );
  OAI21_X1 U743 ( .B1(n558), .B2(n495), .A(n72), .ZN(n70) );
  OAI21_X1 U744 ( .B1(n558), .B2(n78), .A(n79), .ZN(n77) );
  OAI21_X1 U745 ( .B1(n64), .B2(n514), .A(n65), .ZN(n63) );
  NOR2_X1 U746 ( .A1(n234), .A2(n257), .ZN(n113) );
  XOR2_X1 U747 ( .A(n56), .B(n554), .Z(product[5]) );
  XOR2_X1 U748 ( .A(n58), .B(n115), .Z(product[3]) );
  OAI22_X1 U749 ( .A1(n511), .A2(n395), .B1(n394), .B2(n578), .ZN(n316) );
  OAI22_X1 U750 ( .A1(n511), .A2(n394), .B1(n393), .B2(n578), .ZN(n315) );
  OAI22_X1 U751 ( .A1(n511), .A2(n396), .B1(n395), .B2(n578), .ZN(n317) );
  OAI22_X1 U752 ( .A1(n511), .A2(n397), .B1(n396), .B2(n578), .ZN(n318) );
  OAI22_X1 U753 ( .A1(n6), .A2(n398), .B1(n397), .B2(n578), .ZN(n319) );
  OAI22_X1 U754 ( .A1(n511), .A2(n400), .B1(n399), .B2(n578), .ZN(n321) );
  OAI22_X1 U755 ( .A1(n511), .A2(n399), .B1(n398), .B2(n578), .ZN(n320) );
  OAI22_X1 U756 ( .A1(n6), .A2(n401), .B1(n400), .B2(n578), .ZN(n322) );
  OAI22_X1 U757 ( .A1(n6), .A2(n402), .B1(n401), .B2(n578), .ZN(n323) );
  NAND2_X1 U758 ( .A1(n329), .A2(n258), .ZN(n122) );
  OAI22_X1 U759 ( .A1(n6), .A2(n404), .B1(n403), .B2(n578), .ZN(n325) );
  OAI22_X1 U760 ( .A1(n6), .A2(n403), .B1(n402), .B2(n578), .ZN(n324) );
  OAI22_X1 U761 ( .A1(n511), .A2(n406), .B1(n405), .B2(n578), .ZN(n327) );
  OAI22_X1 U762 ( .A1(n511), .A2(n405), .B1(n404), .B2(n578), .ZN(n326) );
  OAI22_X1 U763 ( .A1(n511), .A2(n407), .B1(n406), .B2(n578), .ZN(n328) );
  OAI22_X1 U764 ( .A1(n511), .A2(n408), .B1(n407), .B2(n578), .ZN(n329) );
  OAI22_X1 U765 ( .A1(n6), .A2(n576), .B1(n409), .B2(n578), .ZN(n258) );
  OAI22_X1 U766 ( .A1(n522), .A2(n379), .B1(n378), .B2(n557), .ZN(n301) );
  OAI22_X1 U767 ( .A1(n523), .A2(n380), .B1(n379), .B2(n556), .ZN(n302) );
  OAI22_X1 U768 ( .A1(n523), .A2(n385), .B1(n384), .B2(n556), .ZN(n307) );
  OAI22_X1 U769 ( .A1(n523), .A2(n382), .B1(n381), .B2(n556), .ZN(n304) );
  OAI22_X1 U770 ( .A1(n522), .A2(n381), .B1(n380), .B2(n557), .ZN(n303) );
  NAND2_X1 U771 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U772 ( .A1(n522), .A2(n383), .B1(n382), .B2(n556), .ZN(n305) );
  OAI22_X1 U773 ( .A1(n513), .A2(n384), .B1(n555), .B2(n383), .ZN(n306) );
  OAI22_X1 U774 ( .A1(n513), .A2(n386), .B1(n385), .B2(n557), .ZN(n308) );
  OAI22_X1 U775 ( .A1(n522), .A2(n387), .B1(n386), .B2(n556), .ZN(n309) );
  OAI22_X1 U776 ( .A1(n523), .A2(n583), .B1(n392), .B2(n556), .ZN(n257) );
  OAI22_X1 U777 ( .A1(n389), .A2(n513), .B1(n388), .B2(n555), .ZN(n311) );
  OAI22_X1 U778 ( .A1(n522), .A2(n388), .B1(n387), .B2(n557), .ZN(n310) );
  OAI22_X1 U779 ( .A1(n513), .A2(n390), .B1(n389), .B2(n557), .ZN(n312) );
  INV_X1 U780 ( .A(n557), .ZN(n247) );
  OAI22_X1 U781 ( .A1(n523), .A2(n391), .B1(n390), .B2(n556), .ZN(n313) );
  BUF_X4 U782 ( .A(n43), .Z(n577) );
  INV_X1 U783 ( .A(n586), .ZN(n584) );
  INV_X1 U784 ( .A(n586), .ZN(n585) );
  INV_X1 U785 ( .A(n31), .ZN(n591) );
  INV_X1 U786 ( .A(n593), .ZN(n592) );
  INV_X1 U787 ( .A(n36), .ZN(n593) );
  INV_X1 U788 ( .A(n595), .ZN(n594) );
  INV_X1 U789 ( .A(n40), .ZN(n595) );
  XOR2_X1 U790 ( .A(n259), .B(n251), .Z(n148) );
  XOR2_X1 U791 ( .A(n289), .B(n279), .Z(n146) );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_5_DW01_add_2 ( A, B, CI, 
        SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n5, n8, n9, n10, n11, n12, n13, n14, n15, n16, n19, n20,
         n22, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34, n35, n36, n37,
         n38, n39, n40, n44, n45, n47, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n65, n67, n68, n69, n70, n71, n73,
         n75, n76, n77, n78, n79, n81, n83, n84, n86, n90, n91, n94, n95, n96,
         n98, n100, n157, n158, n159, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181;

  AOI21_X1 U122 ( .B1(n52), .B2(n60), .A(n53), .ZN(n157) );
  OR2_X1 U123 ( .A1(A[13]), .A2(B[13]), .ZN(n158) );
  BUF_X1 U124 ( .A(n171), .Z(n167) );
  NOR2_X1 U125 ( .A1(A[12]), .A2(B[12]), .ZN(n159) );
  NOR2_X1 U126 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  NOR2_X1 U127 ( .A1(A[11]), .A2(B[11]), .ZN(n35) );
  AND2_X1 U128 ( .A1(n175), .A2(n86), .ZN(SUM[0]) );
  XNOR2_X1 U129 ( .A(n45), .B(n161), .ZN(SUM[10]) );
  AND2_X1 U130 ( .A1(n44), .A2(n168), .ZN(n161) );
  XNOR2_X1 U131 ( .A(n37), .B(n162), .ZN(SUM[11]) );
  AND2_X1 U132 ( .A1(n91), .A2(n36), .ZN(n162) );
  XNOR2_X1 U133 ( .A(n1), .B(n163), .ZN(SUM[13]) );
  AND2_X1 U134 ( .A1(n158), .A2(n29), .ZN(n163) );
  NOR2_X1 U135 ( .A1(A[8]), .A2(B[8]), .ZN(n164) );
  NOR2_X1 U136 ( .A1(A[14]), .A2(B[14]), .ZN(n165) );
  NOR2_X1 U137 ( .A1(B[12]), .A2(A[12]), .ZN(n166) );
  NOR2_X1 U138 ( .A1(A[14]), .A2(B[14]), .ZN(n25) );
  OR2_X1 U139 ( .A1(A[10]), .A2(B[10]), .ZN(n168) );
  OR2_X1 U140 ( .A1(A[10]), .A2(B[10]), .ZN(n179) );
  OR2_X1 U141 ( .A1(A[14]), .A2(B[14]), .ZN(n169) );
  INV_X1 U142 ( .A(n167), .ZN(n44) );
  OAI21_X1 U143 ( .B1(n159), .B2(n36), .A(n33), .ZN(n170) );
  AND2_X1 U144 ( .A1(A[10]), .A2(B[10]), .ZN(n171) );
  AOI21_X1 U145 ( .B1(n38), .B2(n30), .A(n170), .ZN(n172) );
  AOI21_X1 U146 ( .B1(n38), .B2(n30), .A(n31), .ZN(n173) );
  INV_X1 U147 ( .A(n24), .ZN(n22) );
  NOR2_X1 U148 ( .A1(A[7]), .A2(B[7]), .ZN(n57) );
  OR2_X1 U149 ( .A1(A[15]), .A2(B[15]), .ZN(n174) );
  OR2_X1 U150 ( .A1(A[9]), .A2(B[9]), .ZN(n180) );
  OR2_X1 U151 ( .A1(A[0]), .A2(B[0]), .ZN(n175) );
  INV_X1 U152 ( .A(n60), .ZN(n59) );
  INV_X1 U153 ( .A(n157), .ZN(n50) );
  INV_X1 U154 ( .A(n67), .ZN(n65) );
  AOI21_X1 U155 ( .B1(n38), .B2(n30), .A(n170), .ZN(n1) );
  AOI21_X1 U156 ( .B1(n177), .B2(n76), .A(n73), .ZN(n71) );
  INV_X1 U157 ( .A(n75), .ZN(n73) );
  OAI21_X1 U158 ( .B1(n79), .B2(n77), .A(n78), .ZN(n76) );
  OR2_X1 U159 ( .A1(n25), .A2(n28), .ZN(n176) );
  AOI21_X1 U160 ( .B1(n52), .B2(n60), .A(n53), .ZN(n51) );
  OAI21_X1 U161 ( .B1(n71), .B2(n69), .A(n70), .ZN(n68) );
  NAND2_X1 U162 ( .A1(n94), .A2(n55), .ZN(n9) );
  INV_X1 U163 ( .A(n86), .ZN(n84) );
  OAI21_X1 U164 ( .B1(n59), .B2(n57), .A(n58), .ZN(n56) );
  AOI21_X1 U165 ( .B1(n178), .B2(n84), .A(n81), .ZN(n79) );
  INV_X1 U166 ( .A(n83), .ZN(n81) );
  NAND2_X1 U167 ( .A1(n98), .A2(n70), .ZN(n13) );
  INV_X1 U168 ( .A(n69), .ZN(n98) );
  INV_X1 U169 ( .A(n166), .ZN(n90) );
  NAND2_X1 U170 ( .A1(n95), .A2(n58), .ZN(n10) );
  INV_X1 U171 ( .A(n57), .ZN(n95) );
  NAND2_X1 U172 ( .A1(n180), .A2(n49), .ZN(n8) );
  NAND2_X1 U173 ( .A1(n100), .A2(n78), .ZN(n15) );
  INV_X1 U174 ( .A(n77), .ZN(n100) );
  NAND2_X1 U175 ( .A1(n181), .A2(n67), .ZN(n12) );
  NAND2_X1 U176 ( .A1(n177), .A2(n75), .ZN(n14) );
  NAND2_X1 U177 ( .A1(n178), .A2(n83), .ZN(n16) );
  NAND2_X1 U178 ( .A1(n96), .A2(n62), .ZN(n11) );
  INV_X1 U179 ( .A(n61), .ZN(n96) );
  XNOR2_X1 U180 ( .A(n12), .B(n68), .ZN(SUM[5]) );
  XOR2_X1 U181 ( .A(n13), .B(n71), .Z(SUM[4]) );
  XOR2_X1 U182 ( .A(n15), .B(n79), .Z(SUM[2]) );
  NAND2_X1 U183 ( .A1(n90), .A2(n33), .ZN(n5) );
  NAND2_X1 U184 ( .A1(n169), .A2(n26), .ZN(n3) );
  NOR2_X1 U185 ( .A1(A[8]), .A2(B[8]), .ZN(n54) );
  NOR2_X1 U186 ( .A1(A[4]), .A2(B[4]), .ZN(n69) );
  NOR2_X1 U187 ( .A1(A[2]), .A2(B[2]), .ZN(n77) );
  NAND2_X1 U188 ( .A1(A[13]), .A2(B[13]), .ZN(n29) );
  NAND2_X1 U189 ( .A1(A[11]), .A2(B[11]), .ZN(n36) );
  OR2_X1 U190 ( .A1(A[3]), .A2(B[3]), .ZN(n177) );
  OR2_X1 U191 ( .A1(A[1]), .A2(B[1]), .ZN(n178) );
  XNOR2_X1 U192 ( .A(n56), .B(n9), .ZN(SUM[8]) );
  XNOR2_X1 U193 ( .A(n14), .B(n76), .ZN(SUM[3]) );
  NOR2_X1 U194 ( .A1(A[6]), .A2(B[6]), .ZN(n61) );
  NAND2_X1 U195 ( .A1(A[7]), .A2(B[7]), .ZN(n58) );
  NAND2_X1 U196 ( .A1(A[4]), .A2(B[4]), .ZN(n70) );
  NAND2_X1 U197 ( .A1(A[2]), .A2(B[2]), .ZN(n78) );
  NAND2_X1 U198 ( .A1(A[15]), .A2(B[15]), .ZN(n19) );
  NAND2_X1 U199 ( .A1(A[5]), .A2(B[5]), .ZN(n67) );
  NAND2_X1 U200 ( .A1(A[3]), .A2(B[3]), .ZN(n75) );
  NAND2_X1 U201 ( .A1(A[1]), .A2(B[1]), .ZN(n83) );
  NAND2_X1 U202 ( .A1(A[0]), .A2(B[0]), .ZN(n86) );
  OR2_X1 U203 ( .A1(A[5]), .A2(B[5]), .ZN(n181) );
  NAND2_X1 U204 ( .A1(A[9]), .A2(B[9]), .ZN(n49) );
  NAND2_X1 U205 ( .A1(A[6]), .A2(B[6]), .ZN(n62) );
  NAND2_X1 U206 ( .A1(A[12]), .A2(B[12]), .ZN(n33) );
  NAND2_X1 U207 ( .A1(A[14]), .A2(B[14]), .ZN(n26) );
  XNOR2_X1 U208 ( .A(n50), .B(n8), .ZN(SUM[9]) );
  XOR2_X1 U209 ( .A(n59), .B(n10), .Z(SUM[7]) );
  XNOR2_X1 U210 ( .A(n16), .B(n84), .ZN(SUM[1]) );
  XOR2_X1 U211 ( .A(n11), .B(n63), .Z(SUM[6]) );
  OAI21_X1 U212 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  AOI21_X1 U213 ( .B1(n181), .B2(n68), .A(n65), .ZN(n63) );
  AOI21_X1 U214 ( .B1(n50), .B2(n180), .A(n47), .ZN(n45) );
  NAND2_X1 U215 ( .A1(n174), .A2(n19), .ZN(n2) );
  XNOR2_X1 U216 ( .A(n20), .B(n2), .ZN(SUM[15]) );
  INV_X1 U217 ( .A(n49), .ZN(n47) );
  INV_X1 U218 ( .A(n164), .ZN(n94) );
  NOR2_X1 U219 ( .A1(n164), .A2(n57), .ZN(n52) );
  OAI21_X1 U220 ( .B1(n54), .B2(n58), .A(n55), .ZN(n53) );
  NAND2_X1 U221 ( .A1(A[8]), .A2(B[8]), .ZN(n55) );
  OAI21_X1 U222 ( .B1(n166), .B2(n36), .A(n33), .ZN(n31) );
  OAI21_X1 U223 ( .B1(n165), .B2(n29), .A(n26), .ZN(n24) );
  OAI21_X1 U224 ( .B1(n37), .B2(n35), .A(n36), .ZN(n34) );
  INV_X1 U225 ( .A(n35), .ZN(n91) );
  NOR2_X1 U226 ( .A1(n159), .A2(n35), .ZN(n30) );
  INV_X1 U227 ( .A(n38), .ZN(n37) );
  NAND2_X1 U228 ( .A1(n168), .A2(n180), .ZN(n39) );
  AOI21_X1 U229 ( .B1(n179), .B2(n47), .A(n171), .ZN(n40) );
  OAI21_X1 U230 ( .B1(n39), .B2(n51), .A(n40), .ZN(n38) );
  XNOR2_X1 U231 ( .A(n34), .B(n5), .ZN(SUM[12]) );
  XNOR2_X1 U232 ( .A(n27), .B(n3), .ZN(SUM[14]) );
  OAI21_X1 U233 ( .B1(n173), .B2(n176), .A(n22), .ZN(n20) );
  OAI21_X1 U234 ( .B1(n172), .B2(n28), .A(n29), .ZN(n27) );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_5 ( clk, clear_acc, 
        data_out_x, data_out, data_out_w, data_out_b, wr_en_y, m_valid, 
        m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [4:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
         N39, N40, N41, N42, N43, N44, n1, n2, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n85, n102, n111, n112, n113, n114, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n22), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n225), .CK(clk), .Q(n26) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n226), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n227), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n228), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n229), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n230), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n231), .CK(clk), .Q(n34) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n232), .CK(clk), .Q(n35) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n233), .CK(clk), .Q(n36) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n234), .CK(clk), .Q(n37) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n235), .CK(clk), .Q(n38) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n236), .CK(clk), .Q(n39) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n237), .CK(clk), .Q(n40) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n238), .CK(clk), .Q(n41) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n239), .CK(clk), .Q(n42) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n240), .CK(clk), .Q(n44) );
  DFF_X1 \f_reg[0]  ( .D(n113), .CK(clk), .Q(f[0]), .QN(n214) );
  DFF_X1 \f_reg[1]  ( .D(n112), .CK(clk), .Q(f[1]), .QN(n215) );
  DFF_X1 \f_reg[2]  ( .D(n111), .CK(clk), .Q(f[2]), .QN(n216) );
  DFF_X1 \f_reg[7]  ( .D(n81), .CK(clk), .Q(f[7]), .QN(n217) );
  DFF_X1 \f_reg[8]  ( .D(n80), .CK(clk), .Q(f[8]), .QN(n218) );
  DFF_X1 \f_reg[9]  ( .D(n79), .CK(clk), .Q(f[9]), .QN(n219) );
  DFF_X1 \f_reg[10]  ( .D(n78), .CK(clk), .Q(n53), .QN(n220) );
  DFF_X1 \f_reg[11]  ( .D(n77), .CK(clk), .Q(n51), .QN(n221) );
  DFF_X1 \f_reg[12]  ( .D(n1), .CK(clk), .Q(n50), .QN(n222) );
  DFF_X1 \f_reg[14]  ( .D(n4), .CK(clk), .Q(n48), .QN(n224) );
  DFF_X1 \f_reg[15]  ( .D(n2), .CK(clk), .Q(f[15]), .QN(n74) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_5_DW_mult_tc_1 mult_2021 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_5_DW01_add_2 add_2022 ( .A({n204, 
        n203, n202, n201, n200, n199, n213, n212, n211, n210, n209, n208, n207, 
        n206, n205, n198}), .B({f[15], n48, n49, n50, n51, n53, f[9:0]}), .CI(
        1'b0), .SUM(adder) );
  DFF_X1 delay_reg ( .D(n114), .CK(clk), .Q(n11), .QN(n241) );
  DFF_X1 \data_out_reg[15]  ( .D(n166), .CK(clk), .Q(data_out[15]), .QN(n197)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n167), .CK(clk), .Q(data_out[14]), .QN(n196)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n168), .CK(clk), .Q(data_out[13]), .QN(n195)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n169), .CK(clk), .Q(data_out[12]), .QN(n194)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n170), .CK(clk), .Q(data_out[11]), .QN(n193)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n171), .CK(clk), .Q(data_out[10]), .QN(n192)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n172), .CK(clk), .Q(data_out[9]), .QN(n191) );
  DFF_X1 \data_out_reg[8]  ( .D(n173), .CK(clk), .Q(data_out[8]), .QN(n190) );
  DFF_X1 \data_out_reg[7]  ( .D(n174), .CK(clk), .Q(data_out[7]), .QN(n189) );
  DFF_X1 \data_out_reg[6]  ( .D(n175), .CK(clk), .Q(data_out[6]), .QN(n188) );
  DFF_X1 \data_out_reg[5]  ( .D(n176), .CK(clk), .Q(data_out[5]), .QN(n187) );
  DFF_X1 \data_out_reg[4]  ( .D(n177), .CK(clk), .Q(data_out[4]), .QN(n186) );
  DFF_X1 \data_out_reg[3]  ( .D(n178), .CK(clk), .Q(data_out[3]), .QN(n185) );
  DFF_X1 \data_out_reg[2]  ( .D(n179), .CK(clk), .Q(data_out[2]), .QN(n184) );
  DFF_X1 \data_out_reg[1]  ( .D(n180), .CK(clk), .Q(data_out[1]), .QN(n183) );
  DFF_X1 \data_out_reg[0]  ( .D(n181), .CK(clk), .Q(data_out[0]), .QN(n182) );
  DFF_X1 \f_reg[3]  ( .D(n102), .CK(clk), .Q(f[3]), .QN(n66) );
  DFF_X1 \f_reg[4]  ( .D(n85), .CK(clk), .Q(f[4]), .QN(n67) );
  DFF_X1 \f_reg[5]  ( .D(n83), .CK(clk), .Q(f[5]), .QN(n68) );
  DFF_X1 \f_reg[6]  ( .D(n82), .CK(clk), .Q(f[6]), .QN(n69) );
  DFF_X2 \f_reg[13]  ( .D(n12), .CK(clk), .Q(n49), .QN(n223) );
  MUX2_X1 U3 ( .A(N39), .B(n33), .S(n11), .Z(n199) );
  AND2_X1 U4 ( .A1(n47), .A2(n23), .ZN(n19) );
  NAND3_X1 U5 ( .A1(n6), .A2(n5), .A3(n7), .ZN(n1) );
  NAND3_X1 U6 ( .A1(n9), .A2(n8), .A3(n10), .ZN(n2) );
  NAND3_X1 U8 ( .A1(n17), .A2(n16), .A3(n18), .ZN(n4) );
  MUX2_X2 U9 ( .A(n35), .B(N37), .S(n241), .Z(n212) );
  MUX2_X2 U10 ( .A(n27), .B(N43), .S(n241), .Z(n203) );
  MUX2_X2 U11 ( .A(n28), .B(N42), .S(n241), .Z(n202) );
  NAND2_X1 U12 ( .A1(data_out_b[12]), .A2(n22), .ZN(n5) );
  NAND2_X1 U13 ( .A1(adder[12]), .A2(n19), .ZN(n6) );
  NAND2_X1 U14 ( .A1(n64), .A2(n50), .ZN(n7) );
  NAND2_X1 U15 ( .A1(data_out_b[15]), .A2(n22), .ZN(n8) );
  NAND2_X1 U16 ( .A1(adder[15]), .A2(n19), .ZN(n9) );
  NAND2_X1 U17 ( .A1(n64), .A2(f[15]), .ZN(n10) );
  INV_X1 U18 ( .A(n47), .ZN(n64) );
  MUX2_X2 U19 ( .A(n29), .B(N41), .S(n241), .Z(n201) );
  MUX2_X2 U20 ( .A(n32), .B(N40), .S(n241), .Z(n200) );
  NAND3_X1 U21 ( .A1(n14), .A2(n13), .A3(n15), .ZN(n12) );
  NAND2_X1 U22 ( .A1(data_out_b[13]), .A2(n22), .ZN(n13) );
  NAND2_X1 U23 ( .A1(adder[13]), .A2(n19), .ZN(n14) );
  NAND2_X1 U24 ( .A1(n64), .A2(n49), .ZN(n15) );
  NAND2_X1 U25 ( .A1(data_out_b[14]), .A2(n22), .ZN(n16) );
  NAND2_X1 U26 ( .A1(adder[14]), .A2(n19), .ZN(n17) );
  NAND2_X1 U27 ( .A1(n64), .A2(n48), .ZN(n18) );
  INV_X1 U28 ( .A(n23), .ZN(n22) );
  NAND2_X1 U29 ( .A1(n114), .A2(n21), .ZN(n243) );
  INV_X1 U30 ( .A(clear_acc), .ZN(n23) );
  INV_X1 U31 ( .A(n25), .ZN(n43) );
  OAI22_X1 U32 ( .A1(n185), .A2(n243), .B1(n66), .B2(n242), .ZN(n178) );
  OAI22_X1 U33 ( .A1(n186), .A2(n243), .B1(n67), .B2(n242), .ZN(n177) );
  OAI22_X1 U34 ( .A1(n187), .A2(n243), .B1(n68), .B2(n242), .ZN(n176) );
  OAI22_X1 U35 ( .A1(n188), .A2(n243), .B1(n69), .B2(n242), .ZN(n175) );
  OAI22_X1 U36 ( .A1(n189), .A2(n243), .B1(n217), .B2(n242), .ZN(n174) );
  OAI22_X1 U37 ( .A1(n190), .A2(n243), .B1(n218), .B2(n242), .ZN(n173) );
  OAI22_X1 U38 ( .A1(n191), .A2(n243), .B1(n219), .B2(n242), .ZN(n172) );
  CLKBUF_X1 U39 ( .A(N39), .Z(n20) );
  INV_X1 U40 ( .A(wr_en_y), .ZN(n21) );
  INV_X1 U41 ( .A(m_ready), .ZN(n24) );
  NAND2_X1 U42 ( .A1(m_valid), .A2(n24), .ZN(n45) );
  OAI21_X1 U43 ( .B1(sel[4]), .B2(n76), .A(n45), .ZN(n114) );
  NAND2_X1 U44 ( .A1(clear_acc_delay), .A2(n241), .ZN(n25) );
  MUX2_X1 U45 ( .A(n26), .B(N44), .S(n43), .Z(n225) );
  MUX2_X1 U46 ( .A(n26), .B(N44), .S(n241), .Z(n204) );
  MUX2_X1 U47 ( .A(n27), .B(N43), .S(n43), .Z(n226) );
  MUX2_X1 U48 ( .A(n28), .B(N42), .S(n43), .Z(n227) );
  MUX2_X1 U49 ( .A(n29), .B(N41), .S(n43), .Z(n228) );
  MUX2_X1 U50 ( .A(n32), .B(N40), .S(n43), .Z(n229) );
  MUX2_X1 U51 ( .A(n33), .B(n20), .S(n43), .Z(n230) );
  MUX2_X1 U52 ( .A(n34), .B(N38), .S(n43), .Z(n231) );
  MUX2_X1 U53 ( .A(n34), .B(N38), .S(n241), .Z(n213) );
  MUX2_X1 U54 ( .A(n35), .B(N37), .S(n43), .Z(n232) );
  MUX2_X1 U55 ( .A(n36), .B(N36), .S(n43), .Z(n233) );
  MUX2_X1 U56 ( .A(n36), .B(N36), .S(n241), .Z(n211) );
  MUX2_X1 U57 ( .A(n37), .B(N35), .S(n43), .Z(n234) );
  MUX2_X1 U58 ( .A(n37), .B(N35), .S(n241), .Z(n210) );
  MUX2_X1 U59 ( .A(n38), .B(N34), .S(n43), .Z(n235) );
  MUX2_X1 U60 ( .A(n38), .B(N34), .S(n241), .Z(n209) );
  MUX2_X1 U61 ( .A(n39), .B(N33), .S(n43), .Z(n236) );
  MUX2_X1 U62 ( .A(n39), .B(N33), .S(n241), .Z(n208) );
  MUX2_X1 U63 ( .A(n40), .B(N32), .S(n43), .Z(n237) );
  MUX2_X1 U64 ( .A(n40), .B(N32), .S(n241), .Z(n207) );
  MUX2_X1 U65 ( .A(n41), .B(N31), .S(n43), .Z(n238) );
  MUX2_X1 U66 ( .A(n41), .B(N31), .S(n241), .Z(n206) );
  MUX2_X1 U67 ( .A(n42), .B(N30), .S(n43), .Z(n239) );
  MUX2_X1 U68 ( .A(n42), .B(N30), .S(n241), .Z(n205) );
  MUX2_X1 U69 ( .A(n44), .B(N29), .S(n43), .Z(n240) );
  MUX2_X1 U70 ( .A(n44), .B(N29), .S(n241), .Z(n198) );
  INV_X1 U71 ( .A(n45), .ZN(n46) );
  OAI21_X1 U72 ( .B1(n46), .B2(n11), .A(n23), .ZN(n47) );
  AOI222_X1 U73 ( .A1(data_out_b[11]), .A2(n22), .B1(adder[11]), .B2(n19), 
        .C1(n64), .C2(n51), .ZN(n52) );
  INV_X1 U74 ( .A(n52), .ZN(n77) );
  AOI222_X1 U75 ( .A1(data_out_b[10]), .A2(n22), .B1(adder[10]), .B2(n19), 
        .C1(n64), .C2(n53), .ZN(n54) );
  INV_X1 U76 ( .A(n54), .ZN(n78) );
  AOI222_X1 U77 ( .A1(data_out_b[8]), .A2(n22), .B1(adder[8]), .B2(n19), .C1(
        n64), .C2(f[8]), .ZN(n55) );
  INV_X1 U78 ( .A(n55), .ZN(n80) );
  AOI222_X1 U79 ( .A1(data_out_b[7]), .A2(n22), .B1(adder[7]), .B2(n19), .C1(
        n64), .C2(f[7]), .ZN(n56) );
  INV_X1 U80 ( .A(n56), .ZN(n81) );
  AOI222_X1 U81 ( .A1(data_out_b[6]), .A2(n22), .B1(adder[6]), .B2(n19), .C1(
        n64), .C2(f[6]), .ZN(n57) );
  INV_X1 U82 ( .A(n57), .ZN(n82) );
  AOI222_X1 U83 ( .A1(data_out_b[5]), .A2(n22), .B1(adder[5]), .B2(n19), .C1(
        n64), .C2(f[5]), .ZN(n58) );
  INV_X1 U84 ( .A(n58), .ZN(n83) );
  AOI222_X1 U85 ( .A1(data_out_b[4]), .A2(n22), .B1(adder[4]), .B2(n19), .C1(
        n64), .C2(f[4]), .ZN(n59) );
  INV_X1 U86 ( .A(n59), .ZN(n85) );
  AOI222_X1 U87 ( .A1(data_out_b[3]), .A2(n22), .B1(adder[3]), .B2(n19), .C1(
        n64), .C2(f[3]), .ZN(n60) );
  INV_X1 U88 ( .A(n60), .ZN(n102) );
  AOI222_X1 U89 ( .A1(data_out_b[2]), .A2(n22), .B1(adder[2]), .B2(n19), .C1(
        n64), .C2(f[2]), .ZN(n61) );
  INV_X1 U90 ( .A(n61), .ZN(n111) );
  AOI222_X1 U91 ( .A1(data_out_b[1]), .A2(n22), .B1(adder[1]), .B2(n19), .C1(
        n64), .C2(f[1]), .ZN(n62) );
  INV_X1 U92 ( .A(n62), .ZN(n112) );
  AOI222_X1 U93 ( .A1(data_out_b[0]), .A2(n22), .B1(adder[0]), .B2(n19), .C1(
        n64), .C2(f[0]), .ZN(n63) );
  INV_X1 U94 ( .A(n63), .ZN(n113) );
  AOI222_X1 U95 ( .A1(data_out_b[9]), .A2(n22), .B1(adder[9]), .B2(n19), .C1(
        n64), .C2(f[9]), .ZN(n65) );
  INV_X1 U96 ( .A(n65), .ZN(n79) );
  NOR4_X1 U97 ( .A1(n51), .A2(n50), .A3(n49), .A4(n48), .ZN(n73) );
  NOR4_X1 U98 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n53), .ZN(n72) );
  NAND4_X1 U99 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(n70) );
  NOR4_X1 U100 ( .A1(n70), .A2(f[0]), .A3(f[1]), .A4(f[2]), .ZN(n71) );
  NAND3_X1 U101 ( .A1(n73), .A2(n72), .A3(n71), .ZN(n75) );
  NAND3_X1 U102 ( .A1(wr_en_y), .A2(n75), .A3(n74), .ZN(n242) );
  OAI22_X1 U103 ( .A1(n182), .A2(n243), .B1(n214), .B2(n242), .ZN(n181) );
  OAI22_X1 U104 ( .A1(n183), .A2(n243), .B1(n215), .B2(n242), .ZN(n180) );
  OAI22_X1 U105 ( .A1(n184), .A2(n243), .B1(n216), .B2(n242), .ZN(n179) );
  OAI22_X1 U106 ( .A1(n192), .A2(n243), .B1(n220), .B2(n242), .ZN(n171) );
  OAI22_X1 U107 ( .A1(n193), .A2(n243), .B1(n221), .B2(n242), .ZN(n170) );
  OAI22_X1 U108 ( .A1(n194), .A2(n243), .B1(n222), .B2(n242), .ZN(n169) );
  OAI22_X1 U109 ( .A1(n195), .A2(n243), .B1(n223), .B2(n242), .ZN(n168) );
  OAI22_X1 U110 ( .A1(n196), .A2(n243), .B1(n224), .B2(n242), .ZN(n167) );
  OAI22_X1 U111 ( .A1(n197), .A2(n243), .B1(n74), .B2(n242), .ZN(n166) );
  AND4_X1 U112 ( .A1(sel[3]), .A2(sel[2]), .A3(sel[1]), .A4(sel[0]), .ZN(n76)
         );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_4_DW_mult_tc_1 ( a, b, 
        product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n9, n12, n13, n16, n18, n19, n21, n25, n27, n29, n31, n32,
         n34, n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n50, n52,
         n53, n54, n55, n56, n57, n58, n59, n62, n63, n64, n65, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n93, n95, n96, n97, n98, n99, n101,
         n103, n104, n105, n106, n107, n111, n112, n113, n114, n115, n117,
         n119, n120, n122, n125, n126, n127, n131, n135, n139, n141, n142,
         n144, n146, n149, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n237, n239, n245, n247, n249, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n418,
         n419, n420, n421, n422, n423, n424, n426, n427, n428, n433, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n263), .CI(n291), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n317), .B(n252), .CO(n173), .S(n174) );
  FA_X1 U169 ( .A(n193), .B(n282), .CI(n191), .CO(n179), .S(n180) );
  FA_X1 U170 ( .A(n268), .B(n292), .CI(n274), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U174 ( .A(n275), .B(n293), .CI(n194), .CO(n189), .S(n190) );
  FA_X1 U175 ( .A(n305), .B(n253), .CI(n283), .CO(n191), .S(n192) );
  HA_X1 U176 ( .A(n269), .B(n319), .CO(n193), .S(n194) );
  FA_X1 U177 ( .A(n205), .B(n200), .CI(n198), .CO(n195), .S(n196) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U179 ( .A(n284), .B(n294), .CI(n276), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n306), .B(n270), .CI(n320), .CO(n201), .S(n202) );
  FA_X1 U181 ( .A(n208), .B(n213), .CI(n206), .CO(n203), .S(n204) );
  FA_X1 U182 ( .A(n215), .B(n307), .CI(n210), .CO(n205), .S(n206) );
  FA_X1 U183 ( .A(n254), .B(n295), .CI(n285), .CO(n207), .S(n208) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U185 ( .A(n216), .B(n219), .CI(n214), .CO(n211), .S(n212) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n308), .B(n278), .CI(n322), .CO(n215), .S(n216) );
  FA_X1 U188 ( .A(n225), .B(n222), .CI(n220), .CO(n217), .S(n218) );
  FA_X1 U189 ( .A(n255), .B(n309), .CI(n297), .CO(n219), .S(n220) );
  HA_X1 U190 ( .A(n323), .B(n287), .CO(n221), .S(n222) );
  FA_X1 U192 ( .A(n310), .B(n288), .CI(n324), .CO(n225), .S(n226) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  HA_X1 U194 ( .A(n325), .B(n311), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n312), .B(n300), .CI(n326), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  BUF_X1 U414 ( .A(n85), .Z(n490) );
  INV_X1 U415 ( .A(n594), .ZN(n491) );
  BUF_X1 U416 ( .A(n497), .Z(n492) );
  BUF_X2 U417 ( .A(n1), .Z(n493) );
  BUF_X1 U418 ( .A(n1), .Z(n497) );
  OR2_X1 U419 ( .A1(n329), .A2(n258), .ZN(n494) );
  CLKBUF_X1 U420 ( .A(n12), .Z(n495) );
  FA_X1 U421 ( .A(n205), .B(n200), .CI(n198), .S(n496) );
  INV_X1 U422 ( .A(n601), .ZN(n498) );
  XNOR2_X1 U423 ( .A(n301), .B(n499), .ZN(n149) );
  XNOR2_X1 U424 ( .A(n259), .B(n251), .ZN(n499) );
  XNOR2_X1 U425 ( .A(n500), .B(n501), .ZN(n585) );
  XNOR2_X1 U426 ( .A(n265), .B(n144), .ZN(n500) );
  XNOR2_X1 U427 ( .A(n161), .B(n142), .ZN(n501) );
  XNOR2_X1 U428 ( .A(n502), .B(n188), .ZN(n186) );
  XNOR2_X1 U429 ( .A(n197), .B(n190), .ZN(n502) );
  XOR2_X1 U430 ( .A(n596), .B(a[4]), .Z(n16) );
  XNOR2_X1 U431 ( .A(n503), .B(n166), .ZN(n164) );
  XNOR2_X1 U432 ( .A(n177), .B(n168), .ZN(n503) );
  INV_X1 U433 ( .A(n509), .ZN(n504) );
  NAND2_X1 U434 ( .A1(n196), .A2(n203), .ZN(n505) );
  BUF_X2 U435 ( .A(n9), .Z(n506) );
  CLKBUF_X1 U436 ( .A(n9), .Z(n588) );
  OAI21_X1 U437 ( .B1(n82), .B2(n505), .A(n83), .ZN(n507) );
  AOI21_X1 U438 ( .B1(n582), .B2(n104), .A(n101), .ZN(n508) );
  CLKBUF_X1 U439 ( .A(n602), .Z(n509) );
  INV_X1 U440 ( .A(n515), .ZN(n510) );
  XNOR2_X1 U441 ( .A(n149), .B(n511), .ZN(n144) );
  XNOR2_X1 U442 ( .A(n146), .B(n271), .ZN(n511) );
  INV_X1 U443 ( .A(n603), .ZN(n512) );
  INV_X1 U444 ( .A(n603), .ZN(n602) );
  BUF_X1 U445 ( .A(n37), .Z(n513) );
  OR2_X1 U446 ( .A1(n496), .A2(n203), .ZN(n514) );
  INV_X1 U447 ( .A(n595), .ZN(n515) );
  XNOR2_X1 U448 ( .A(n516), .B(n179), .ZN(n166) );
  XNOR2_X1 U449 ( .A(n170), .B(n172), .ZN(n516) );
  INV_X1 U450 ( .A(n541), .ZN(n517) );
  XNOR2_X1 U451 ( .A(n518), .B(n189), .ZN(n178) );
  XNOR2_X1 U452 ( .A(n182), .B(n184), .ZN(n518) );
  NOR2_X1 U453 ( .A1(n186), .A2(n195), .ZN(n519) );
  NOR2_X1 U454 ( .A1(n186), .A2(n195), .ZN(n82) );
  INV_X1 U455 ( .A(n549), .ZN(n520) );
  BUF_X2 U456 ( .A(n600), .Z(n549) );
  XNOR2_X1 U457 ( .A(n596), .B(a[2]), .ZN(n575) );
  XOR2_X1 U458 ( .A(n199), .B(n201), .Z(n521) );
  XOR2_X1 U459 ( .A(n521), .B(n192), .Z(n188) );
  NAND2_X1 U460 ( .A1(n199), .A2(n201), .ZN(n522) );
  NAND2_X1 U461 ( .A1(n199), .A2(n192), .ZN(n523) );
  NAND2_X1 U462 ( .A1(n201), .A2(n192), .ZN(n524) );
  NAND3_X1 U463 ( .A1(n522), .A2(n523), .A3(n524), .ZN(n187) );
  NAND2_X1 U464 ( .A1(n197), .A2(n190), .ZN(n525) );
  NAND2_X1 U465 ( .A1(n197), .A2(n188), .ZN(n526) );
  NAND2_X1 U466 ( .A1(n190), .A2(n188), .ZN(n527) );
  NAND3_X1 U467 ( .A1(n525), .A2(n526), .A3(n527), .ZN(n185) );
  INV_X1 U468 ( .A(n239), .ZN(n545) );
  XNOR2_X1 U469 ( .A(n45), .B(n528), .ZN(product[12]) );
  AND2_X1 U470 ( .A1(n126), .A2(n79), .ZN(n528) );
  OR2_X2 U471 ( .A1(n542), .A2(n574), .ZN(n538) );
  OR2_X2 U472 ( .A1(n529), .A2(n563), .ZN(n29) );
  XNOR2_X1 U473 ( .A(n602), .B(a[8]), .ZN(n529) );
  NAND2_X1 U474 ( .A1(n170), .A2(n172), .ZN(n530) );
  NAND2_X1 U475 ( .A1(n170), .A2(n179), .ZN(n531) );
  NAND2_X1 U476 ( .A1(n172), .A2(n179), .ZN(n532) );
  NAND3_X1 U477 ( .A1(n530), .A2(n531), .A3(n532), .ZN(n165) );
  NAND2_X1 U478 ( .A1(n177), .A2(n168), .ZN(n533) );
  NAND2_X1 U479 ( .A1(n177), .A2(n166), .ZN(n534) );
  NAND2_X1 U480 ( .A1(n168), .A2(n166), .ZN(n535) );
  NAND3_X1 U481 ( .A1(n533), .A2(n534), .A3(n535), .ZN(n163) );
  INV_X1 U482 ( .A(n574), .ZN(n21) );
  BUF_X1 U483 ( .A(n16), .Z(n536) );
  INV_X1 U484 ( .A(n594), .ZN(n537) );
  INV_X1 U485 ( .A(n594), .ZN(n593) );
  OR2_X1 U486 ( .A1(n204), .A2(n211), .ZN(n539) );
  NOR2_X1 U487 ( .A1(n164), .A2(n175), .ZN(n540) );
  NOR2_X1 U488 ( .A1(n164), .A2(n175), .ZN(n75) );
  INV_X1 U489 ( .A(n599), .ZN(n541) );
  XNOR2_X1 U490 ( .A(n498), .B(a[6]), .ZN(n542) );
  CLKBUF_X1 U491 ( .A(n573), .Z(n543) );
  AOI21_X1 U492 ( .B1(n96), .B2(n578), .A(n93), .ZN(n544) );
  XOR2_X1 U493 ( .A(n603), .B(a[10]), .Z(n32) );
  INV_X1 U494 ( .A(n605), .ZN(n546) );
  INV_X1 U495 ( .A(n605), .ZN(n547) );
  INV_X2 U496 ( .A(n563), .ZN(n27) );
  OAI21_X1 U497 ( .B1(n91), .B2(n89), .A(n90), .ZN(n548) );
  OAI21_X1 U498 ( .B1(n544), .B2(n89), .A(n90), .ZN(n88) );
  BUF_X2 U499 ( .A(n600), .Z(n550) );
  INV_X1 U500 ( .A(n601), .ZN(n600) );
  NAND2_X1 U501 ( .A1(n576), .A2(n536), .ZN(n551) );
  INV_X2 U502 ( .A(n596), .ZN(n595) );
  XOR2_X1 U503 ( .A(n180), .B(n187), .Z(n552) );
  XOR2_X1 U504 ( .A(n552), .B(n178), .Z(n176) );
  NAND2_X1 U505 ( .A1(n182), .A2(n184), .ZN(n553) );
  NAND2_X1 U506 ( .A1(n182), .A2(n189), .ZN(n554) );
  NAND2_X1 U507 ( .A1(n184), .A2(n189), .ZN(n555) );
  NAND3_X1 U508 ( .A1(n553), .A2(n554), .A3(n555), .ZN(n177) );
  NAND2_X1 U509 ( .A1(n180), .A2(n187), .ZN(n556) );
  NAND2_X1 U510 ( .A1(n180), .A2(n178), .ZN(n557) );
  NAND2_X1 U511 ( .A1(n187), .A2(n178), .ZN(n558) );
  NAND3_X1 U512 ( .A1(n556), .A2(n557), .A3(n558), .ZN(n175) );
  CLKBUF_X1 U513 ( .A(n104), .Z(n559) );
  CLKBUF_X1 U514 ( .A(n562), .Z(n560) );
  INV_X2 U515 ( .A(n249), .ZN(n592) );
  XNOR2_X1 U516 ( .A(n88), .B(n561), .ZN(product[10]) );
  NAND2_X1 U517 ( .A1(n514), .A2(n86), .ZN(n561) );
  NAND2_X1 U518 ( .A1(n575), .A2(n9), .ZN(n562) );
  NAND2_X1 U519 ( .A1(n9), .A2(n575), .ZN(n12) );
  XNOR2_X1 U520 ( .A(n601), .B(a[8]), .ZN(n563) );
  NAND2_X1 U521 ( .A1(n433), .A2(n592), .ZN(n564) );
  NAND2_X1 U522 ( .A1(n433), .A2(n592), .ZN(n565) );
  NAND2_X1 U523 ( .A1(n433), .A2(n592), .ZN(n6) );
  AND2_X1 U524 ( .A1(n232), .A2(n233), .ZN(n566) );
  OR2_X1 U525 ( .A1(n228), .A2(n231), .ZN(n567) );
  XOR2_X1 U526 ( .A(n229), .B(n298), .Z(n568) );
  XOR2_X1 U527 ( .A(n226), .B(n568), .Z(n224) );
  NAND2_X1 U528 ( .A1(n226), .A2(n229), .ZN(n569) );
  NAND2_X1 U529 ( .A1(n226), .A2(n298), .ZN(n570) );
  NAND2_X1 U530 ( .A1(n229), .A2(n298), .ZN(n571) );
  NAND3_X1 U531 ( .A1(n569), .A2(n570), .A3(n571), .ZN(n223) );
  CLKBUF_X3 U532 ( .A(n16), .Z(n587) );
  CLKBUF_X1 U533 ( .A(n107), .Z(n572) );
  AOI21_X1 U534 ( .B1(n548), .B2(n80), .A(n507), .ZN(n573) );
  XNOR2_X1 U535 ( .A(n599), .B(a[6]), .ZN(n574) );
  NAND2_X1 U536 ( .A1(n576), .A2(n536), .ZN(n18) );
  XOR2_X1 U537 ( .A(n597), .B(a[4]), .Z(n576) );
  BUF_X1 U538 ( .A(n43), .Z(n590) );
  INV_X1 U539 ( .A(n69), .ZN(n67) );
  NAND2_X1 U540 ( .A1(n577), .A2(n69), .ZN(n47) );
  INV_X1 U541 ( .A(n73), .ZN(n71) );
  NAND2_X1 U542 ( .A1(n577), .A2(n73), .ZN(n64) );
  INV_X1 U543 ( .A(n74), .ZN(n72) );
  AOI21_X1 U544 ( .B1(n80), .B2(n88), .A(n81), .ZN(n45) );
  NAND2_X1 U545 ( .A1(n90), .A2(n539), .ZN(n52) );
  INV_X1 U546 ( .A(n78), .ZN(n126) );
  OR2_X1 U547 ( .A1(n152), .A2(n163), .ZN(n577) );
  OAI21_X1 U548 ( .B1(n540), .B2(n79), .A(n76), .ZN(n74) );
  NAND2_X1 U549 ( .A1(n125), .A2(n76), .ZN(n48) );
  INV_X1 U550 ( .A(n75), .ZN(n125) );
  NOR2_X1 U551 ( .A1(n75), .A2(n78), .ZN(n73) );
  XNOR2_X1 U552 ( .A(n84), .B(n50), .ZN(product[11]) );
  NAND2_X1 U553 ( .A1(n127), .A2(n83), .ZN(n50) );
  NAND2_X1 U554 ( .A1(n152), .A2(n163), .ZN(n69) );
  INV_X1 U555 ( .A(n95), .ZN(n93) );
  AOI21_X1 U556 ( .B1(n582), .B2(n104), .A(n101), .ZN(n99) );
  OAI21_X1 U557 ( .B1(n113), .B2(n115), .A(n114), .ZN(n112) );
  NOR2_X1 U558 ( .A1(n176), .A2(n185), .ZN(n78) );
  NAND2_X1 U559 ( .A1(n578), .A2(n95), .ZN(n53) );
  AOI21_X1 U560 ( .B1(n579), .B2(n120), .A(n117), .ZN(n115) );
  INV_X1 U561 ( .A(n119), .ZN(n117) );
  INV_X1 U562 ( .A(n122), .ZN(n120) );
  NOR2_X1 U563 ( .A1(n196), .A2(n203), .ZN(n85) );
  XNOR2_X1 U564 ( .A(n63), .B(n46), .ZN(product[15]) );
  NAND2_X1 U565 ( .A1(n581), .A2(n62), .ZN(n46) );
  AOI21_X1 U566 ( .B1(n74), .B2(n577), .A(n67), .ZN(n65) );
  XNOR2_X1 U567 ( .A(n57), .B(n112), .ZN(product[4]) );
  NAND2_X1 U568 ( .A1(n580), .A2(n111), .ZN(n57) );
  XNOR2_X1 U569 ( .A(n59), .B(n120), .ZN(product[2]) );
  NAND2_X1 U570 ( .A1(n579), .A2(n119), .ZN(n59) );
  NAND2_X1 U571 ( .A1(n176), .A2(n185), .ZN(n79) );
  NAND2_X1 U572 ( .A1(n164), .A2(n175), .ZN(n76) );
  NAND2_X1 U573 ( .A1(n212), .A2(n217), .ZN(n95) );
  OR2_X1 U574 ( .A1(n212), .A2(n217), .ZN(n578) );
  NAND2_X1 U575 ( .A1(n204), .A2(n211), .ZN(n90) );
  NAND2_X1 U576 ( .A1(n496), .A2(n203), .ZN(n86) );
  NAND2_X1 U577 ( .A1(n135), .A2(n114), .ZN(n58) );
  NAND2_X1 U578 ( .A1(n131), .A2(n98), .ZN(n54) );
  INV_X1 U579 ( .A(n97), .ZN(n131) );
  NAND2_X1 U580 ( .A1(n567), .A2(n106), .ZN(n56) );
  NOR2_X1 U581 ( .A1(n218), .A2(n223), .ZN(n97) );
  OR2_X1 U582 ( .A1(n328), .A2(n314), .ZN(n579) );
  NOR2_X1 U583 ( .A1(n228), .A2(n231), .ZN(n105) );
  NAND2_X1 U584 ( .A1(n218), .A2(n223), .ZN(n98) );
  NAND2_X1 U585 ( .A1(n228), .A2(n231), .ZN(n106) );
  INV_X1 U586 ( .A(n37), .ZN(n237) );
  OR2_X1 U587 ( .A1(n232), .A2(n233), .ZN(n580) );
  INV_X1 U588 ( .A(n41), .ZN(n235) );
  OR2_X1 U589 ( .A1(n139), .A2(n151), .ZN(n581) );
  OR2_X1 U590 ( .A1(n224), .A2(n227), .ZN(n582) );
  AND2_X1 U591 ( .A1(n494), .A2(n122), .ZN(product[1]) );
  XNOR2_X1 U592 ( .A(n604), .B(a[12]), .ZN(n37) );
  XNOR2_X1 U593 ( .A(n606), .B(a[14]), .ZN(n41) );
  OR2_X1 U594 ( .A1(n590), .A2(n515), .ZN(n392) );
  OR2_X1 U595 ( .A1(n590), .A2(n517), .ZN(n377) );
  XOR2_X1 U596 ( .A(n604), .B(a[10]), .Z(n428) );
  XNOR2_X1 U597 ( .A(n512), .B(n590), .ZN(n352) );
  OAI22_X1 U598 ( .A1(n39), .A2(n336), .B1(n513), .B2(n335), .ZN(n263) );
  OAI22_X1 U599 ( .A1(n42), .A2(n609), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U600 ( .A1(n590), .A2(n609), .ZN(n332) );
  XNOR2_X1 U601 ( .A(n546), .B(n590), .ZN(n343) );
  AND2_X1 U602 ( .A1(n591), .A2(n245), .ZN(n300) );
  XNOR2_X1 U603 ( .A(n155), .B(n584), .ZN(n139) );
  XNOR2_X1 U604 ( .A(n153), .B(n141), .ZN(n584) );
  XNOR2_X1 U605 ( .A(n157), .B(n585), .ZN(n141) );
  XNOR2_X1 U606 ( .A(n159), .B(n586), .ZN(n142) );
  XNOR2_X1 U607 ( .A(n315), .B(n261), .ZN(n586) );
  XNOR2_X1 U608 ( .A(n606), .B(n590), .ZN(n336) );
  NAND2_X1 U609 ( .A1(n427), .A2(n37), .ZN(n39) );
  XOR2_X1 U610 ( .A(n606), .B(a[12]), .Z(n427) );
  XNOR2_X1 U611 ( .A(n598), .B(n590), .ZN(n376) );
  AND2_X1 U612 ( .A1(n591), .A2(n237), .ZN(n264) );
  AND2_X1 U613 ( .A1(n591), .A2(n235), .ZN(n260) );
  OAI22_X1 U614 ( .A1(n39), .A2(n335), .B1(n513), .B2(n334), .ZN(n262) );
  AND2_X1 U615 ( .A1(n591), .A2(n574), .ZN(n288) );
  AND2_X1 U616 ( .A1(n591), .A2(n239), .ZN(n270) );
  INV_X1 U617 ( .A(n19), .ZN(n601) );
  INV_X1 U618 ( .A(n25), .ZN(n603) );
  AND2_X1 U619 ( .A1(n591), .A2(n563), .ZN(n278) );
  INV_X1 U620 ( .A(n1), .ZN(n594) );
  NAND2_X1 U621 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U622 ( .A(n608), .B(a[14]), .Z(n426) );
  INV_X1 U623 ( .A(n7), .ZN(n596) );
  XNOR2_X1 U624 ( .A(n549), .B(n590), .ZN(n363) );
  OAI22_X1 U625 ( .A1(n39), .A2(n607), .B1(n337), .B2(n513), .ZN(n252) );
  OR2_X1 U626 ( .A1(n590), .A2(n607), .ZN(n337) );
  AND2_X1 U627 ( .A1(n591), .A2(n247), .ZN(n314) );
  AND2_X1 U628 ( .A1(n591), .A2(n249), .ZN(product[0]) );
  OR2_X1 U629 ( .A1(n590), .A2(n605), .ZN(n344) );
  OR2_X1 U630 ( .A1(n590), .A2(n520), .ZN(n364) );
  OR2_X1 U631 ( .A1(n590), .A2(n504), .ZN(n353) );
  XNOR2_X1 U632 ( .A(n549), .B(b[9]), .ZN(n354) );
  OAI22_X1 U633 ( .A1(n39), .A2(n334), .B1(n513), .B2(n333), .ZN(n261) );
  XNOR2_X1 U634 ( .A(n606), .B(n422), .ZN(n333) );
  XNOR2_X1 U635 ( .A(n598), .B(b[11]), .ZN(n365) );
  XNOR2_X1 U636 ( .A(n606), .B(n424), .ZN(n335) );
  XNOR2_X1 U637 ( .A(n606), .B(n423), .ZN(n334) );
  OAI22_X1 U638 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U639 ( .A(n608), .B(n424), .ZN(n330) );
  XNOR2_X1 U640 ( .A(n608), .B(n590), .ZN(n331) );
  XNOR2_X1 U641 ( .A(n512), .B(n418), .ZN(n345) );
  XNOR2_X1 U642 ( .A(n546), .B(n420), .ZN(n338) );
  XNOR2_X1 U643 ( .A(n510), .B(b[13]), .ZN(n378) );
  XNOR2_X1 U644 ( .A(n547), .B(n424), .ZN(n342) );
  XNOR2_X1 U645 ( .A(n550), .B(n424), .ZN(n362) );
  XNOR2_X1 U646 ( .A(n602), .B(n424), .ZN(n351) );
  XNOR2_X1 U647 ( .A(n546), .B(n423), .ZN(n341) );
  XNOR2_X1 U648 ( .A(n547), .B(n422), .ZN(n340) );
  XNOR2_X1 U649 ( .A(n547), .B(n421), .ZN(n339) );
  XNOR2_X1 U650 ( .A(n595), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U651 ( .A(n595), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U652 ( .A(n595), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U653 ( .A(n595), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U654 ( .A(n510), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U655 ( .A(n595), .B(n418), .ZN(n384) );
  XNOR2_X1 U656 ( .A(n595), .B(n419), .ZN(n385) );
  XNOR2_X1 U657 ( .A(n550), .B(n423), .ZN(n361) );
  XNOR2_X1 U658 ( .A(n512), .B(n423), .ZN(n350) );
  XNOR2_X1 U659 ( .A(n598), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U660 ( .A(n598), .B(n418), .ZN(n369) );
  XNOR2_X1 U661 ( .A(n598), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U662 ( .A(n598), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U663 ( .A(n602), .B(n422), .ZN(n349) );
  XNOR2_X1 U664 ( .A(n549), .B(n422), .ZN(n360) );
  XNOR2_X1 U665 ( .A(n550), .B(n421), .ZN(n359) );
  XNOR2_X1 U666 ( .A(n509), .B(n421), .ZN(n348) );
  XNOR2_X1 U667 ( .A(n593), .B(b[11]), .ZN(n397) );
  XNOR2_X1 U668 ( .A(n491), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U669 ( .A(n497), .B(b[13]), .ZN(n395) );
  XNOR2_X1 U670 ( .A(n491), .B(b[14]), .ZN(n394) );
  XNOR2_X1 U671 ( .A(n549), .B(n420), .ZN(n358) );
  XNOR2_X1 U672 ( .A(n512), .B(n420), .ZN(n347) );
  XNOR2_X1 U673 ( .A(n550), .B(n418), .ZN(n356) );
  XNOR2_X1 U674 ( .A(n549), .B(n419), .ZN(n357) );
  XNOR2_X1 U675 ( .A(n512), .B(n419), .ZN(n346) );
  XNOR2_X1 U676 ( .A(n550), .B(b[8]), .ZN(n355) );
  BUF_X1 U677 ( .A(n43), .Z(n591) );
  XNOR2_X1 U678 ( .A(n593), .B(b[15]), .ZN(n393) );
  OAI22_X1 U679 ( .A1(n34), .A2(n339), .B1(n338), .B2(n545), .ZN(n265) );
  OAI22_X1 U680 ( .A1(n34), .A2(n340), .B1(n339), .B2(n545), .ZN(n266) );
  OAI22_X1 U681 ( .A1(n34), .A2(n341), .B1(n340), .B2(n545), .ZN(n267) );
  OAI22_X1 U682 ( .A1(n34), .A2(n342), .B1(n341), .B2(n545), .ZN(n268) );
  INV_X1 U683 ( .A(n32), .ZN(n239) );
  OAI22_X1 U684 ( .A1(n34), .A2(n343), .B1(n342), .B2(n545), .ZN(n269) );
  OAI22_X1 U685 ( .A1(n34), .A2(n605), .B1(n344), .B2(n545), .ZN(n253) );
  NAND2_X1 U686 ( .A1(n428), .A2(n32), .ZN(n34) );
  XNOR2_X1 U687 ( .A(n1), .B(a[2]), .ZN(n9) );
  INV_X1 U688 ( .A(n13), .ZN(n599) );
  NAND2_X1 U689 ( .A1(n582), .A2(n103), .ZN(n55) );
  INV_X1 U690 ( .A(n103), .ZN(n101) );
  NAND2_X1 U691 ( .A1(n224), .A2(n227), .ZN(n103) );
  AOI21_X1 U692 ( .B1(n580), .B2(n112), .A(n566), .ZN(n107) );
  INV_X1 U693 ( .A(n519), .ZN(n127) );
  NOR2_X1 U694 ( .A1(n519), .A2(n85), .ZN(n80) );
  OAI21_X1 U695 ( .B1(n82), .B2(n86), .A(n83), .ZN(n81) );
  NAND2_X1 U696 ( .A1(n186), .A2(n195), .ZN(n83) );
  OAI21_X1 U697 ( .B1(n99), .B2(n97), .A(n98), .ZN(n589) );
  OAI21_X1 U698 ( .B1(n508), .B2(n97), .A(n98), .ZN(n96) );
  NOR2_X1 U699 ( .A1(n204), .A2(n211), .ZN(n89) );
  OAI22_X1 U700 ( .A1(n29), .A2(n346), .B1(n345), .B2(n27), .ZN(n271) );
  OAI22_X1 U701 ( .A1(n29), .A2(n350), .B1(n349), .B2(n27), .ZN(n275) );
  OAI22_X1 U702 ( .A1(n29), .A2(n347), .B1(n346), .B2(n27), .ZN(n272) );
  OAI22_X1 U703 ( .A1(n29), .A2(n348), .B1(n347), .B2(n27), .ZN(n273) );
  OAI22_X1 U704 ( .A1(n29), .A2(n349), .B1(n348), .B2(n27), .ZN(n274) );
  OAI22_X1 U705 ( .A1(n29), .A2(n504), .B1(n353), .B2(n27), .ZN(n254) );
  OAI22_X1 U706 ( .A1(n29), .A2(n351), .B1(n350), .B2(n27), .ZN(n276) );
  OAI22_X1 U707 ( .A1(n29), .A2(n352), .B1(n351), .B2(n27), .ZN(n277) );
  INV_X1 U708 ( .A(n113), .ZN(n135) );
  AOI21_X1 U709 ( .B1(n96), .B2(n578), .A(n93), .ZN(n91) );
  OR2_X1 U710 ( .A1(n590), .A2(n594), .ZN(n409) );
  XNOR2_X1 U711 ( .A(n77), .B(n48), .ZN(product[13]) );
  XNOR2_X1 U712 ( .A(n55), .B(n559), .ZN(product[6]) );
  XOR2_X1 U713 ( .A(n56), .B(n572), .Z(product[5]) );
  OAI21_X1 U714 ( .B1(n105), .B2(n107), .A(n106), .ZN(n104) );
  XNOR2_X1 U715 ( .A(n70), .B(n47), .ZN(product[14]) );
  OAI21_X1 U716 ( .B1(n87), .B2(n490), .A(n505), .ZN(n84) );
  NAND2_X1 U717 ( .A1(n151), .A2(n139), .ZN(n62) );
  OAI22_X1 U718 ( .A1(n538), .A2(n358), .B1(n357), .B2(n21), .ZN(n282) );
  OAI22_X1 U719 ( .A1(n538), .A2(n362), .B1(n361), .B2(n21), .ZN(n286) );
  OAI22_X1 U720 ( .A1(n538), .A2(n356), .B1(n355), .B2(n21), .ZN(n280) );
  OAI22_X1 U721 ( .A1(n538), .A2(n520), .B1(n364), .B2(n21), .ZN(n255) );
  OAI22_X1 U722 ( .A1(n538), .A2(n360), .B1(n359), .B2(n21), .ZN(n284) );
  OAI22_X1 U723 ( .A1(n538), .A2(n361), .B1(n360), .B2(n21), .ZN(n285) );
  OAI22_X1 U724 ( .A1(n538), .A2(n357), .B1(n356), .B2(n21), .ZN(n281) );
  OAI22_X1 U725 ( .A1(n538), .A2(n363), .B1(n362), .B2(n21), .ZN(n287) );
  XNOR2_X1 U726 ( .A(n541), .B(n423), .ZN(n374) );
  XNOR2_X1 U727 ( .A(n597), .B(n422), .ZN(n373) );
  XNOR2_X1 U728 ( .A(n541), .B(n421), .ZN(n372) );
  OAI22_X1 U729 ( .A1(n538), .A2(n359), .B1(n358), .B2(n21), .ZN(n283) );
  XNOR2_X1 U730 ( .A(n541), .B(n424), .ZN(n375) );
  XNOR2_X1 U731 ( .A(n597), .B(n419), .ZN(n370) );
  OAI22_X1 U732 ( .A1(n538), .A2(n355), .B1(n354), .B2(n21), .ZN(n279) );
  XNOR2_X1 U733 ( .A(n597), .B(n420), .ZN(n371) );
  INV_X1 U734 ( .A(n548), .ZN(n87) );
  NAND2_X1 U735 ( .A1(n232), .A2(n233), .ZN(n111) );
  OAI22_X1 U736 ( .A1(n18), .A2(n370), .B1(n369), .B2(n587), .ZN(n293) );
  OAI22_X1 U737 ( .A1(n18), .A2(n367), .B1(n366), .B2(n587), .ZN(n290) );
  OAI22_X1 U738 ( .A1(n18), .A2(n368), .B1(n367), .B2(n587), .ZN(n291) );
  OAI22_X1 U739 ( .A1(n369), .A2(n551), .B1(n368), .B2(n587), .ZN(n292) );
  OAI22_X1 U740 ( .A1(n551), .A2(n372), .B1(n371), .B2(n587), .ZN(n295) );
  OAI22_X1 U741 ( .A1(n551), .A2(n371), .B1(n370), .B2(n587), .ZN(n294) );
  OAI22_X1 U742 ( .A1(n18), .A2(n375), .B1(n374), .B2(n587), .ZN(n298) );
  OAI22_X1 U743 ( .A1(n18), .A2(n373), .B1(n372), .B2(n587), .ZN(n296) );
  OAI22_X1 U744 ( .A1(n551), .A2(n374), .B1(n373), .B2(n587), .ZN(n297) );
  OAI22_X1 U745 ( .A1(n18), .A2(n517), .B1(n377), .B2(n587), .ZN(n256) );
  OAI22_X1 U746 ( .A1(n18), .A2(n376), .B1(n375), .B2(n587), .ZN(n299) );
  OAI22_X1 U747 ( .A1(n551), .A2(n366), .B1(n365), .B2(n587), .ZN(n289) );
  XNOR2_X1 U748 ( .A(n595), .B(n420), .ZN(n386) );
  XNOR2_X1 U749 ( .A(n595), .B(n590), .ZN(n391) );
  INV_X1 U750 ( .A(n16), .ZN(n245) );
  XNOR2_X1 U751 ( .A(n595), .B(n422), .ZN(n388) );
  XNOR2_X1 U752 ( .A(n595), .B(n421), .ZN(n387) );
  XNOR2_X1 U753 ( .A(n595), .B(n423), .ZN(n389) );
  XNOR2_X1 U754 ( .A(n595), .B(n424), .ZN(n390) );
  NAND2_X1 U755 ( .A1(n328), .A2(n314), .ZN(n119) );
  XNOR2_X1 U756 ( .A(n493), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U757 ( .A(n537), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U758 ( .A(n492), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U759 ( .A(n493), .B(n418), .ZN(n401) );
  XNOR2_X1 U760 ( .A(n537), .B(n420), .ZN(n403) );
  XNOR2_X1 U761 ( .A(n493), .B(n419), .ZN(n402) );
  XNOR2_X1 U762 ( .A(n492), .B(n421), .ZN(n404) );
  XNOR2_X1 U763 ( .A(n491), .B(n422), .ZN(n405) );
  XNOR2_X1 U764 ( .A(n593), .B(n590), .ZN(n408) );
  XNOR2_X1 U765 ( .A(n493), .B(n424), .ZN(n407) );
  XNOR2_X1 U766 ( .A(n493), .B(n423), .ZN(n406) );
  XOR2_X1 U767 ( .A(n1), .B(n249), .Z(n433) );
  NOR2_X1 U768 ( .A1(n234), .A2(n257), .ZN(n113) );
  OAI21_X1 U769 ( .B1(n64), .B2(n543), .A(n65), .ZN(n63) );
  OAI21_X1 U770 ( .B1(n573), .B2(n71), .A(n72), .ZN(n70) );
  OAI21_X1 U771 ( .B1(n45), .B2(n78), .A(n79), .ZN(n77) );
  XOR2_X1 U772 ( .A(n91), .B(n52), .Z(product[9]) );
  XNOR2_X1 U773 ( .A(n53), .B(n589), .ZN(product[8]) );
  XOR2_X1 U774 ( .A(n58), .B(n115), .Z(product[3]) );
  OAI22_X1 U775 ( .A1(n565), .A2(n395), .B1(n394), .B2(n592), .ZN(n316) );
  OAI22_X1 U776 ( .A1(n564), .A2(n394), .B1(n393), .B2(n592), .ZN(n315) );
  OAI22_X1 U777 ( .A1(n564), .A2(n396), .B1(n395), .B2(n592), .ZN(n317) );
  OAI22_X1 U778 ( .A1(n565), .A2(n397), .B1(n396), .B2(n592), .ZN(n318) );
  OAI22_X1 U779 ( .A1(n565), .A2(n398), .B1(n397), .B2(n592), .ZN(n319) );
  OAI22_X1 U780 ( .A1(n565), .A2(n400), .B1(n399), .B2(n592), .ZN(n321) );
  OAI22_X1 U781 ( .A1(n6), .A2(n399), .B1(n398), .B2(n592), .ZN(n320) );
  OAI22_X1 U782 ( .A1(n564), .A2(n401), .B1(n400), .B2(n592), .ZN(n322) );
  OAI22_X1 U783 ( .A1(n564), .A2(n402), .B1(n401), .B2(n592), .ZN(n323) );
  NAND2_X1 U784 ( .A1(n329), .A2(n258), .ZN(n122) );
  OAI22_X1 U785 ( .A1(n6), .A2(n404), .B1(n403), .B2(n592), .ZN(n325) );
  OAI22_X1 U786 ( .A1(n564), .A2(n403), .B1(n402), .B2(n592), .ZN(n324) );
  OAI22_X1 U787 ( .A1(n6), .A2(n406), .B1(n405), .B2(n592), .ZN(n327) );
  OAI22_X1 U788 ( .A1(n565), .A2(n405), .B1(n404), .B2(n592), .ZN(n326) );
  OAI22_X1 U789 ( .A1(n564), .A2(n407), .B1(n406), .B2(n592), .ZN(n328) );
  OAI22_X1 U790 ( .A1(n6), .A2(n408), .B1(n407), .B2(n592), .ZN(n329) );
  OAI22_X1 U791 ( .A1(n6), .A2(n594), .B1(n409), .B2(n592), .ZN(n258) );
  XOR2_X1 U792 ( .A(n99), .B(n54), .Z(product[7]) );
  OAI22_X1 U793 ( .A1(n560), .A2(n379), .B1(n378), .B2(n506), .ZN(n301) );
  OAI22_X1 U794 ( .A1(n495), .A2(n380), .B1(n379), .B2(n506), .ZN(n302) );
  OAI22_X1 U795 ( .A1(n560), .A2(n385), .B1(n384), .B2(n506), .ZN(n307) );
  OAI22_X1 U796 ( .A1(n12), .A2(n382), .B1(n381), .B2(n506), .ZN(n304) );
  OAI22_X1 U797 ( .A1(n562), .A2(n381), .B1(n380), .B2(n506), .ZN(n303) );
  NAND2_X1 U798 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U799 ( .A1(n12), .A2(n383), .B1(n382), .B2(n506), .ZN(n305) );
  OAI22_X1 U800 ( .A1(n12), .A2(n384), .B1(n383), .B2(n588), .ZN(n306) );
  OAI22_X1 U801 ( .A1(n12), .A2(n386), .B1(n385), .B2(n588), .ZN(n308) );
  OAI22_X1 U802 ( .A1(n562), .A2(n387), .B1(n386), .B2(n506), .ZN(n309) );
  OAI22_X1 U803 ( .A1(n562), .A2(n515), .B1(n392), .B2(n506), .ZN(n257) );
  OAI22_X1 U804 ( .A1(n12), .A2(n389), .B1(n388), .B2(n588), .ZN(n311) );
  OAI22_X1 U805 ( .A1(n562), .A2(n388), .B1(n387), .B2(n506), .ZN(n310) );
  OAI22_X1 U806 ( .A1(n562), .A2(n390), .B1(n389), .B2(n506), .ZN(n312) );
  INV_X1 U807 ( .A(n506), .ZN(n247) );
  OAI22_X1 U808 ( .A1(n562), .A2(n391), .B1(n390), .B2(n506), .ZN(n313) );
  INV_X1 U809 ( .A(n599), .ZN(n597) );
  INV_X1 U810 ( .A(n599), .ZN(n598) );
  INV_X1 U811 ( .A(n605), .ZN(n604) );
  INV_X1 U812 ( .A(n31), .ZN(n605) );
  INV_X1 U813 ( .A(n607), .ZN(n606) );
  INV_X1 U814 ( .A(n36), .ZN(n607) );
  INV_X1 U815 ( .A(n609), .ZN(n608) );
  INV_X1 U816 ( .A(n40), .ZN(n609) );
  XOR2_X1 U817 ( .A(n289), .B(n279), .Z(n146) );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_4_DW01_add_2 ( A, B, CI, 
        SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n19, n20, n22, n24, n25, n26, n27, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n44, n45, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n65, n67, n68, n69, n70, n71,
         n73, n75, n76, n77, n78, n79, n81, n83, n84, n86, n90, n94, n95, n96,
         n98, n100, n157, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185;

  CLKBUF_X1 U122 ( .A(n30), .Z(n157) );
  NOR2_X1 U123 ( .A1(A[14]), .A2(B[14]), .ZN(n25) );
  AND2_X1 U124 ( .A1(n180), .A2(n86), .ZN(SUM[0]) );
  OR2_X1 U125 ( .A1(n25), .A2(n167), .ZN(n159) );
  OR2_X1 U126 ( .A1(A[15]), .A2(B[15]), .ZN(n160) );
  NOR2_X1 U127 ( .A1(A[8]), .A2(B[8]), .ZN(n161) );
  NOR2_X1 U128 ( .A1(A[8]), .A2(B[8]), .ZN(n54) );
  OR2_X1 U129 ( .A1(A[13]), .A2(B[13]), .ZN(n162) );
  XNOR2_X1 U130 ( .A(n172), .B(n6), .ZN(SUM[11]) );
  XNOR2_X1 U131 ( .A(n1), .B(n163), .ZN(SUM[13]) );
  AND2_X1 U132 ( .A1(n162), .A2(n29), .ZN(n163) );
  AOI21_X1 U133 ( .B1(n52), .B2(n60), .A(n53), .ZN(n164) );
  AOI21_X1 U134 ( .B1(n52), .B2(n60), .A(n53), .ZN(n165) );
  OR2_X1 U135 ( .A1(A[11]), .A2(B[11]), .ZN(n166) );
  NOR2_X1 U136 ( .A1(A[13]), .A2(B[13]), .ZN(n167) );
  NOR2_X1 U137 ( .A1(n35), .A2(n170), .ZN(n30) );
  AOI21_X1 U138 ( .B1(n184), .B2(n47), .A(n177), .ZN(n168) );
  NOR2_X1 U139 ( .A1(A[12]), .A2(B[12]), .ZN(n169) );
  NOR2_X1 U140 ( .A1(A[12]), .A2(B[12]), .ZN(n170) );
  NOR2_X1 U141 ( .A1(A[12]), .A2(B[12]), .ZN(n32) );
  OR2_X1 U142 ( .A1(A[14]), .A2(B[14]), .ZN(n171) );
  OAI21_X1 U143 ( .B1(n39), .B2(n164), .A(n40), .ZN(n172) );
  NAND2_X1 U144 ( .A1(A[11]), .A2(B[11]), .ZN(n173) );
  NAND2_X1 U145 ( .A1(A[11]), .A2(B[11]), .ZN(n36) );
  OR2_X1 U146 ( .A1(A[10]), .A2(B[10]), .ZN(n174) );
  OR2_X1 U147 ( .A1(A[10]), .A2(B[10]), .ZN(n184) );
  OAI21_X1 U148 ( .B1(n32), .B2(n36), .A(n33), .ZN(n175) );
  INV_X1 U149 ( .A(n177), .ZN(n44) );
  INV_X1 U150 ( .A(n166), .ZN(n176) );
  AND2_X1 U151 ( .A1(A[10]), .A2(B[10]), .ZN(n177) );
  AOI21_X1 U152 ( .B1(n30), .B2(n38), .A(n175), .ZN(n178) );
  AOI21_X1 U153 ( .B1(n30), .B2(n38), .A(n31), .ZN(n179) );
  OR2_X1 U154 ( .A1(A[0]), .A2(B[0]), .ZN(n180) );
  OAI21_X1 U155 ( .B1(n71), .B2(n69), .A(n70), .ZN(n68) );
  AOI21_X1 U156 ( .B1(n38), .B2(n157), .A(n175), .ZN(n1) );
  AOI21_X1 U157 ( .B1(n182), .B2(n84), .A(n81), .ZN(n79) );
  INV_X1 U158 ( .A(n83), .ZN(n81) );
  OAI21_X1 U159 ( .B1(n79), .B2(n77), .A(n78), .ZN(n76) );
  AOI21_X1 U160 ( .B1(n185), .B2(n68), .A(n65), .ZN(n63) );
  INV_X1 U161 ( .A(n67), .ZN(n65) );
  INV_X1 U162 ( .A(n24), .ZN(n22) );
  AOI21_X1 U163 ( .B1(n183), .B2(n76), .A(n73), .ZN(n71) );
  INV_X1 U164 ( .A(n75), .ZN(n73) );
  AOI21_X1 U165 ( .B1(n50), .B2(n181), .A(n47), .ZN(n45) );
  NAND2_X1 U166 ( .A1(n94), .A2(n55), .ZN(n9) );
  INV_X1 U167 ( .A(n86), .ZN(n84) );
  OAI21_X1 U168 ( .B1(n59), .B2(n57), .A(n58), .ZN(n56) );
  INV_X1 U169 ( .A(n49), .ZN(n47) );
  INV_X1 U170 ( .A(n170), .ZN(n90) );
  NAND2_X1 U171 ( .A1(n183), .A2(n75), .ZN(n14) );
  NAND2_X1 U172 ( .A1(n95), .A2(n58), .ZN(n10) );
  INV_X1 U173 ( .A(n57), .ZN(n95) );
  NAND2_X1 U174 ( .A1(n181), .A2(n49), .ZN(n8) );
  NAND2_X1 U175 ( .A1(n100), .A2(n78), .ZN(n15) );
  INV_X1 U176 ( .A(n77), .ZN(n100) );
  NAND2_X1 U177 ( .A1(n185), .A2(n67), .ZN(n12) );
  NAND2_X1 U178 ( .A1(n182), .A2(n83), .ZN(n16) );
  NAND2_X1 U179 ( .A1(n98), .A2(n70), .ZN(n13) );
  INV_X1 U180 ( .A(n69), .ZN(n98) );
  NAND2_X1 U181 ( .A1(n96), .A2(n62), .ZN(n11) );
  INV_X1 U182 ( .A(n61), .ZN(n96) );
  XNOR2_X1 U183 ( .A(n12), .B(n68), .ZN(SUM[5]) );
  NAND2_X1 U184 ( .A1(n171), .A2(n26), .ZN(n3) );
  NAND2_X1 U185 ( .A1(n90), .A2(n33), .ZN(n5) );
  NOR2_X1 U186 ( .A1(A[7]), .A2(B[7]), .ZN(n57) );
  NOR2_X1 U187 ( .A1(A[11]), .A2(B[11]), .ZN(n35) );
  OR2_X1 U188 ( .A1(A[9]), .A2(B[9]), .ZN(n181) );
  NOR2_X1 U189 ( .A1(A[2]), .A2(B[2]), .ZN(n77) );
  XOR2_X1 U190 ( .A(n59), .B(n10), .Z(SUM[7]) );
  NAND2_X1 U191 ( .A1(A[13]), .A2(B[13]), .ZN(n29) );
  OR2_X1 U192 ( .A1(A[1]), .A2(B[1]), .ZN(n182) );
  OR2_X1 U193 ( .A1(A[3]), .A2(B[3]), .ZN(n183) );
  NOR2_X1 U194 ( .A1(A[4]), .A2(B[4]), .ZN(n69) );
  XNOR2_X1 U195 ( .A(n56), .B(n9), .ZN(SUM[8]) );
  XNOR2_X1 U196 ( .A(n14), .B(n76), .ZN(SUM[3]) );
  XNOR2_X1 U197 ( .A(n16), .B(n84), .ZN(SUM[1]) );
  NOR2_X1 U198 ( .A1(A[6]), .A2(B[6]), .ZN(n61) );
  NAND2_X1 U199 ( .A1(A[7]), .A2(B[7]), .ZN(n58) );
  OR2_X1 U200 ( .A1(A[5]), .A2(B[5]), .ZN(n185) );
  NAND2_X1 U201 ( .A1(A[2]), .A2(B[2]), .ZN(n78) );
  NAND2_X1 U202 ( .A1(A[9]), .A2(B[9]), .ZN(n49) );
  NAND2_X1 U203 ( .A1(A[5]), .A2(B[5]), .ZN(n67) );
  NAND2_X1 U204 ( .A1(A[1]), .A2(B[1]), .ZN(n83) );
  NAND2_X1 U205 ( .A1(A[0]), .A2(B[0]), .ZN(n86) );
  NAND2_X1 U206 ( .A1(A[4]), .A2(B[4]), .ZN(n70) );
  NAND2_X1 U207 ( .A1(A[6]), .A2(B[6]), .ZN(n62) );
  NAND2_X1 U208 ( .A1(A[14]), .A2(B[14]), .ZN(n26) );
  XOR2_X1 U209 ( .A(n45), .B(n7), .Z(SUM[10]) );
  XNOR2_X1 U210 ( .A(n50), .B(n8), .ZN(SUM[9]) );
  XOR2_X1 U211 ( .A(n15), .B(n79), .Z(SUM[2]) );
  NAND2_X1 U212 ( .A1(n160), .A2(n19), .ZN(n2) );
  INV_X1 U213 ( .A(n165), .ZN(n50) );
  INV_X1 U214 ( .A(n60), .ZN(n59) );
  OAI21_X1 U215 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  INV_X1 U216 ( .A(n161), .ZN(n94) );
  NOR2_X1 U217 ( .A1(n161), .A2(n57), .ZN(n52) );
  OAI21_X1 U218 ( .B1(n54), .B2(n58), .A(n55), .ZN(n53) );
  NAND2_X1 U219 ( .A1(A[8]), .A2(B[8]), .ZN(n55) );
  XOR2_X1 U220 ( .A(n11), .B(n63), .Z(SUM[6]) );
  NAND2_X1 U221 ( .A1(A[12]), .A2(B[12]), .ZN(n33) );
  XOR2_X1 U222 ( .A(n13), .B(n71), .Z(SUM[4]) );
  NAND2_X1 U223 ( .A1(A[3]), .A2(B[3]), .ZN(n75) );
  INV_X1 U224 ( .A(n172), .ZN(n37) );
  OAI21_X1 U225 ( .B1(n25), .B2(n29), .A(n26), .ZN(n24) );
  OAI21_X1 U226 ( .B1(n169), .B2(n173), .A(n33), .ZN(n31) );
  NAND2_X1 U227 ( .A1(n166), .A2(n173), .ZN(n6) );
  NAND2_X1 U228 ( .A1(A[15]), .A2(B[15]), .ZN(n19) );
  OAI21_X1 U229 ( .B1(n37), .B2(n176), .A(n173), .ZN(n34) );
  OAI21_X1 U230 ( .B1(n39), .B2(n164), .A(n168), .ZN(n38) );
  NAND2_X1 U231 ( .A1(n174), .A2(n181), .ZN(n39) );
  AOI21_X1 U232 ( .B1(n184), .B2(n47), .A(n177), .ZN(n40) );
  NAND2_X1 U233 ( .A1(n174), .A2(n44), .ZN(n7) );
  XNOR2_X1 U234 ( .A(n34), .B(n5), .ZN(SUM[12]) );
  XNOR2_X1 U235 ( .A(n20), .B(n2), .ZN(SUM[15]) );
  XNOR2_X1 U236 ( .A(n27), .B(n3), .ZN(SUM[14]) );
  OAI21_X1 U237 ( .B1(n179), .B2(n167), .A(n29), .ZN(n27) );
  OAI21_X1 U238 ( .B1(n178), .B2(n159), .A(n22), .ZN(n20) );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_4 ( clk, clear_acc, 
        data_out_x, data_out, data_out_w, data_out_b, wr_en_y, m_valid, 
        m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [4:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
         N39, N40, N41, N42, N43, N44, n1, n2, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n85, n102, n111, n112, n113, n114, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n22), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n221), .CK(clk), .Q(n25) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n222), .CK(clk), .Q(n26) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n223), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n224), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n225), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n226), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n227), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n228), .CK(clk), .Q(n34) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n229), .CK(clk), .Q(n35) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n230), .CK(clk), .Q(n36) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n231), .CK(clk), .Q(n37) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n232), .CK(clk), .Q(n38) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n233), .CK(clk), .Q(n39) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n234), .CK(clk), .Q(n40) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n235), .CK(clk), .Q(n41) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n236), .CK(clk), .Q(n42) );
  DFF_X1 \f_reg[0]  ( .D(n111), .CK(clk), .Q(f[0]), .QN(n210) );
  DFF_X1 \f_reg[1]  ( .D(n102), .CK(clk), .Q(f[1]), .QN(n211) );
  DFF_X1 \f_reg[2]  ( .D(n85), .CK(clk), .Q(f[2]), .QN(n212) );
  DFF_X1 \f_reg[7]  ( .D(n79), .CK(clk), .Q(f[7]), .QN(n213) );
  DFF_X1 \f_reg[8]  ( .D(n78), .CK(clk), .Q(f[8]), .QN(n214) );
  DFF_X1 \f_reg[9]  ( .D(n77), .CK(clk), .Q(f[9]), .QN(n215) );
  DFF_X1 \f_reg[10]  ( .D(n76), .CK(clk), .Q(n51), .QN(n216) );
  DFF_X1 \f_reg[11]  ( .D(n75), .CK(clk), .Q(n49), .QN(n217) );
  DFF_X1 \f_reg[12]  ( .D(n2), .CK(clk), .Q(n48), .QN(n218) );
  DFF_X1 \f_reg[13]  ( .D(n4), .CK(clk), .Q(n47), .QN(n219) );
  DFF_X1 \f_reg[14]  ( .D(n8), .CK(clk), .Q(n46), .QN(n220) );
  DFF_X1 \f_reg[15]  ( .D(n9), .CK(clk), .Q(f[15]), .QN(n72) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_4_DW_mult_tc_1 mult_2021 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_4_DW01_add_2 add_2022 ( .A({n200, 
        n199, n198, n197, n196, n195, n209, n208, n207, n206, n205, n204, n203, 
        n202, n201, n194}), .B({f[15], n46, n47, n48, n49, n51, f[9:0]}), .CI(
        1'b0), .SUM(adder) );
  DFF_X1 delay_reg ( .D(n112), .CK(clk), .Q(n19), .QN(n237) );
  DFF_X1 \data_out_reg[15]  ( .D(n113), .CK(clk), .Q(data_out[15]), .QN(n193)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n114), .CK(clk), .Q(data_out[14]), .QN(n192)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n164), .CK(clk), .Q(data_out[13]), .QN(n191)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n165), .CK(clk), .Q(data_out[12]), .QN(n190)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n166), .CK(clk), .Q(data_out[11]), .QN(n189)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n167), .CK(clk), .Q(data_out[10]), .QN(n188)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n168), .CK(clk), .Q(data_out[9]), .QN(n187) );
  DFF_X1 \data_out_reg[8]  ( .D(n169), .CK(clk), .Q(data_out[8]), .QN(n186) );
  DFF_X1 \data_out_reg[7]  ( .D(n170), .CK(clk), .Q(data_out[7]), .QN(n185) );
  DFF_X1 \data_out_reg[6]  ( .D(n171), .CK(clk), .Q(data_out[6]), .QN(n184) );
  DFF_X1 \data_out_reg[5]  ( .D(n172), .CK(clk), .Q(data_out[5]), .QN(n183) );
  DFF_X1 \data_out_reg[4]  ( .D(n173), .CK(clk), .Q(data_out[4]), .QN(n182) );
  DFF_X1 \data_out_reg[3]  ( .D(n174), .CK(clk), .Q(data_out[3]), .QN(n181) );
  DFF_X1 \data_out_reg[2]  ( .D(n175), .CK(clk), .Q(data_out[2]), .QN(n180) );
  DFF_X1 \data_out_reg[1]  ( .D(n176), .CK(clk), .Q(data_out[1]), .QN(n179) );
  DFF_X1 \data_out_reg[0]  ( .D(n177), .CK(clk), .Q(data_out[0]), .QN(n178) );
  DFF_X1 \f_reg[3]  ( .D(n83), .CK(clk), .Q(f[3]), .QN(n64) );
  DFF_X1 \f_reg[4]  ( .D(n82), .CK(clk), .Q(f[4]), .QN(n65) );
  DFF_X1 \f_reg[5]  ( .D(n81), .CK(clk), .Q(f[5]), .QN(n66) );
  DFF_X1 \f_reg[6]  ( .D(n80), .CK(clk), .Q(f[6]), .QN(n67) );
  AND2_X1 U3 ( .A1(clear_acc_delay), .A2(n237), .ZN(n1) );
  INV_X1 U4 ( .A(n45), .ZN(n62) );
  AND2_X1 U5 ( .A1(n45), .A2(n23), .ZN(n20) );
  NAND3_X1 U6 ( .A1(n11), .A2(n10), .A3(n12), .ZN(n2) );
  NAND3_X1 U8 ( .A1(n6), .A2(n5), .A3(n7), .ZN(n4) );
  NAND2_X1 U9 ( .A1(data_out_b[13]), .A2(n22), .ZN(n5) );
  NAND2_X1 U10 ( .A1(adder[13]), .A2(n20), .ZN(n6) );
  NAND2_X1 U11 ( .A1(n62), .A2(n47), .ZN(n7) );
  MUX2_X2 U12 ( .A(n34), .B(N37), .S(n237), .Z(n208) );
  NAND3_X1 U13 ( .A1(n17), .A2(n16), .A3(n18), .ZN(n8) );
  NAND3_X1 U14 ( .A1(n14), .A2(n13), .A3(n15), .ZN(n9) );
  MUX2_X2 U15 ( .A(n28), .B(N41), .S(n237), .Z(n197) );
  NAND2_X1 U16 ( .A1(data_out_b[12]), .A2(n22), .ZN(n10) );
  NAND2_X1 U17 ( .A1(adder[12]), .A2(n20), .ZN(n11) );
  NAND2_X1 U18 ( .A1(n62), .A2(n48), .ZN(n12) );
  NAND2_X1 U19 ( .A1(data_out_b[15]), .A2(n22), .ZN(n13) );
  NAND2_X1 U20 ( .A1(adder[15]), .A2(n20), .ZN(n14) );
  NAND2_X1 U21 ( .A1(n62), .A2(f[15]), .ZN(n15) );
  NAND2_X1 U22 ( .A1(data_out_b[14]), .A2(n22), .ZN(n16) );
  NAND2_X1 U23 ( .A1(adder[14]), .A2(n20), .ZN(n17) );
  NAND2_X1 U24 ( .A1(n62), .A2(n46), .ZN(n18) );
  MUX2_X2 U25 ( .A(n26), .B(N43), .S(n237), .Z(n199) );
  MUX2_X2 U26 ( .A(n27), .B(N42), .S(n237), .Z(n198) );
  MUX2_X2 U27 ( .A(n29), .B(N40), .S(n237), .Z(n196) );
  MUX2_X2 U28 ( .A(N39), .B(n32), .S(n19), .Z(n195) );
  INV_X1 U29 ( .A(n23), .ZN(n22) );
  NAND2_X1 U30 ( .A1(n112), .A2(n21), .ZN(n239) );
  INV_X1 U31 ( .A(clear_acc), .ZN(n23) );
  OAI22_X1 U32 ( .A1(n181), .A2(n239), .B1(n64), .B2(n238), .ZN(n174) );
  OAI22_X1 U33 ( .A1(n182), .A2(n239), .B1(n65), .B2(n238), .ZN(n173) );
  OAI22_X1 U34 ( .A1(n183), .A2(n239), .B1(n66), .B2(n238), .ZN(n172) );
  OAI22_X1 U35 ( .A1(n184), .A2(n239), .B1(n67), .B2(n238), .ZN(n171) );
  OAI22_X1 U36 ( .A1(n185), .A2(n239), .B1(n213), .B2(n238), .ZN(n170) );
  OAI22_X1 U37 ( .A1(n186), .A2(n239), .B1(n214), .B2(n238), .ZN(n169) );
  OAI22_X1 U38 ( .A1(n187), .A2(n239), .B1(n215), .B2(n238), .ZN(n168) );
  INV_X1 U39 ( .A(wr_en_y), .ZN(n21) );
  INV_X1 U40 ( .A(m_ready), .ZN(n24) );
  NAND2_X1 U41 ( .A1(m_valid), .A2(n24), .ZN(n43) );
  OAI21_X1 U42 ( .B1(sel[4]), .B2(n74), .A(n43), .ZN(n112) );
  MUX2_X1 U43 ( .A(n25), .B(N44), .S(n1), .Z(n221) );
  MUX2_X1 U44 ( .A(n25), .B(N44), .S(n237), .Z(n200) );
  MUX2_X1 U45 ( .A(n26), .B(N43), .S(n1), .Z(n222) );
  MUX2_X1 U46 ( .A(n27), .B(N42), .S(n1), .Z(n223) );
  MUX2_X1 U47 ( .A(n28), .B(N41), .S(n1), .Z(n224) );
  MUX2_X1 U48 ( .A(n29), .B(N40), .S(n1), .Z(n225) );
  MUX2_X1 U49 ( .A(n32), .B(N39), .S(n1), .Z(n226) );
  MUX2_X1 U50 ( .A(n33), .B(N38), .S(n1), .Z(n227) );
  MUX2_X1 U51 ( .A(n33), .B(N38), .S(n237), .Z(n209) );
  MUX2_X1 U52 ( .A(n34), .B(N37), .S(n1), .Z(n228) );
  MUX2_X1 U53 ( .A(n35), .B(N36), .S(n1), .Z(n229) );
  MUX2_X1 U54 ( .A(n35), .B(N36), .S(n237), .Z(n207) );
  MUX2_X1 U55 ( .A(n36), .B(N35), .S(n1), .Z(n230) );
  MUX2_X1 U56 ( .A(n36), .B(N35), .S(n237), .Z(n206) );
  MUX2_X1 U57 ( .A(n37), .B(N34), .S(n1), .Z(n231) );
  MUX2_X1 U58 ( .A(n37), .B(N34), .S(n237), .Z(n205) );
  MUX2_X1 U59 ( .A(n38), .B(N33), .S(n1), .Z(n232) );
  MUX2_X1 U60 ( .A(n38), .B(N33), .S(n237), .Z(n204) );
  MUX2_X1 U61 ( .A(n39), .B(N32), .S(n1), .Z(n233) );
  MUX2_X1 U62 ( .A(n39), .B(N32), .S(n237), .Z(n203) );
  MUX2_X1 U63 ( .A(n40), .B(N31), .S(n1), .Z(n234) );
  MUX2_X1 U64 ( .A(n40), .B(N31), .S(n237), .Z(n202) );
  MUX2_X1 U65 ( .A(n41), .B(N30), .S(n1), .Z(n235) );
  MUX2_X1 U66 ( .A(n41), .B(N30), .S(n237), .Z(n201) );
  MUX2_X1 U67 ( .A(n42), .B(N29), .S(n1), .Z(n236) );
  MUX2_X1 U68 ( .A(n42), .B(N29), .S(n237), .Z(n194) );
  INV_X1 U69 ( .A(n43), .ZN(n44) );
  OAI21_X1 U70 ( .B1(n44), .B2(n19), .A(n23), .ZN(n45) );
  AOI222_X1 U71 ( .A1(data_out_b[11]), .A2(n22), .B1(adder[11]), .B2(n20), 
        .C1(n62), .C2(n49), .ZN(n50) );
  INV_X1 U72 ( .A(n50), .ZN(n75) );
  AOI222_X1 U73 ( .A1(data_out_b[10]), .A2(n22), .B1(adder[10]), .B2(n20), 
        .C1(n62), .C2(n51), .ZN(n52) );
  INV_X1 U74 ( .A(n52), .ZN(n76) );
  AOI222_X1 U75 ( .A1(data_out_b[8]), .A2(n22), .B1(adder[8]), .B2(n20), .C1(
        n62), .C2(f[8]), .ZN(n53) );
  INV_X1 U76 ( .A(n53), .ZN(n78) );
  AOI222_X1 U77 ( .A1(data_out_b[7]), .A2(n22), .B1(adder[7]), .B2(n20), .C1(
        n62), .C2(f[7]), .ZN(n54) );
  INV_X1 U78 ( .A(n54), .ZN(n79) );
  AOI222_X1 U79 ( .A1(data_out_b[6]), .A2(n22), .B1(adder[6]), .B2(n20), .C1(
        n62), .C2(f[6]), .ZN(n55) );
  INV_X1 U80 ( .A(n55), .ZN(n80) );
  AOI222_X1 U81 ( .A1(data_out_b[5]), .A2(n22), .B1(adder[5]), .B2(n20), .C1(
        n62), .C2(f[5]), .ZN(n56) );
  INV_X1 U82 ( .A(n56), .ZN(n81) );
  AOI222_X1 U83 ( .A1(data_out_b[4]), .A2(n22), .B1(adder[4]), .B2(n20), .C1(
        n62), .C2(f[4]), .ZN(n57) );
  INV_X1 U84 ( .A(n57), .ZN(n82) );
  AOI222_X1 U85 ( .A1(data_out_b[3]), .A2(n22), .B1(adder[3]), .B2(n20), .C1(
        n62), .C2(f[3]), .ZN(n58) );
  INV_X1 U86 ( .A(n58), .ZN(n83) );
  AOI222_X1 U87 ( .A1(data_out_b[2]), .A2(n22), .B1(adder[2]), .B2(n20), .C1(
        n62), .C2(f[2]), .ZN(n59) );
  INV_X1 U88 ( .A(n59), .ZN(n85) );
  AOI222_X1 U89 ( .A1(data_out_b[1]), .A2(n22), .B1(adder[1]), .B2(n20), .C1(
        n62), .C2(f[1]), .ZN(n60) );
  INV_X1 U90 ( .A(n60), .ZN(n102) );
  AOI222_X1 U91 ( .A1(data_out_b[0]), .A2(n22), .B1(adder[0]), .B2(n20), .C1(
        n62), .C2(f[0]), .ZN(n61) );
  INV_X1 U92 ( .A(n61), .ZN(n111) );
  AOI222_X1 U93 ( .A1(data_out_b[9]), .A2(n22), .B1(adder[9]), .B2(n20), .C1(
        n62), .C2(f[9]), .ZN(n63) );
  INV_X1 U94 ( .A(n63), .ZN(n77) );
  NOR4_X1 U95 ( .A1(n49), .A2(n48), .A3(n47), .A4(n46), .ZN(n71) );
  NOR4_X1 U96 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n51), .ZN(n70) );
  NAND4_X1 U97 ( .A1(n67), .A2(n66), .A3(n65), .A4(n64), .ZN(n68) );
  NOR4_X1 U98 ( .A1(n68), .A2(f[0]), .A3(f[1]), .A4(f[2]), .ZN(n69) );
  NAND3_X1 U99 ( .A1(n71), .A2(n70), .A3(n69), .ZN(n73) );
  NAND3_X1 U100 ( .A1(wr_en_y), .A2(n73), .A3(n72), .ZN(n238) );
  OAI22_X1 U101 ( .A1(n178), .A2(n239), .B1(n210), .B2(n238), .ZN(n177) );
  OAI22_X1 U102 ( .A1(n179), .A2(n239), .B1(n211), .B2(n238), .ZN(n176) );
  OAI22_X1 U103 ( .A1(n180), .A2(n239), .B1(n212), .B2(n238), .ZN(n175) );
  OAI22_X1 U104 ( .A1(n188), .A2(n239), .B1(n216), .B2(n238), .ZN(n167) );
  OAI22_X1 U105 ( .A1(n189), .A2(n239), .B1(n217), .B2(n238), .ZN(n166) );
  OAI22_X1 U106 ( .A1(n190), .A2(n239), .B1(n218), .B2(n238), .ZN(n165) );
  OAI22_X1 U107 ( .A1(n191), .A2(n239), .B1(n219), .B2(n238), .ZN(n164) );
  OAI22_X1 U108 ( .A1(n192), .A2(n239), .B1(n220), .B2(n238), .ZN(n114) );
  OAI22_X1 U109 ( .A1(n193), .A2(n239), .B1(n72), .B2(n238), .ZN(n113) );
  AND4_X1 U110 ( .A1(sel[3]), .A2(sel[2]), .A3(sel[1]), .A4(sel[0]), .ZN(n74)
         );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_3_DW_mult_tc_1 ( a, b, 
        product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n9, n12, n13, n16, n18, n19, n21, n23, n25, n27, n29, n31,
         n34, n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n50,
         n53, n54, n55, n56, n57, n58, n59, n62, n63, n64, n65, n67, n69, n70,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n93, n95, n96, n97, n98, n99, n101,
         n103, n104, n105, n106, n107, n109, n111, n112, n113, n114, n115,
         n117, n119, n120, n122, n125, n127, n129, n131, n133, n135, n139,
         n141, n142, n144, n146, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n237, n241, n247, n249, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n418, n419, n420, n421, n422, n423, n424, n426, n427,
         n429, n433, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U152 ( .A(n301), .B(n148), .Z(n149) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n263), .CI(n291), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n317), .B(n252), .CO(n173), .S(n174) );
  FA_X1 U167 ( .A(n180), .B(n187), .CI(n178), .CO(n175), .S(n176) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U169 ( .A(n193), .B(n282), .CI(n191), .CO(n179), .S(n180) );
  FA_X1 U170 ( .A(n268), .B(n274), .CI(n292), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U172 ( .A(n197), .B(n190), .CI(n188), .CO(n185), .S(n186) );
  FA_X1 U173 ( .A(n199), .B(n201), .CI(n192), .CO(n187), .S(n188) );
  FA_X1 U174 ( .A(n275), .B(n293), .CI(n194), .CO(n189), .S(n190) );
  FA_X1 U175 ( .A(n283), .B(n305), .CI(n253), .CO(n191), .S(n192) );
  HA_X1 U176 ( .A(n269), .B(n319), .CO(n193), .S(n194) );
  FA_X1 U177 ( .A(n205), .B(n200), .CI(n198), .CO(n195), .S(n196) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U179 ( .A(n276), .B(n284), .CI(n294), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n306), .B(n270), .CI(n320), .CO(n201), .S(n202) );
  FA_X1 U181 ( .A(n208), .B(n213), .CI(n206), .CO(n203), .S(n204) );
  FA_X1 U182 ( .A(n210), .B(n307), .CI(n215), .CO(n205), .S(n206) );
  FA_X1 U183 ( .A(n254), .B(n285), .CI(n295), .CO(n207), .S(n208) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U185 ( .A(n216), .B(n219), .CI(n214), .CO(n211), .S(n212) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n322), .B(n278), .CI(n308), .CO(n215), .S(n216) );
  FA_X1 U188 ( .A(n225), .B(n222), .CI(n220), .CO(n217), .S(n218) );
  FA_X1 U189 ( .A(n255), .B(n309), .CI(n297), .CO(n219), .S(n220) );
  HA_X1 U190 ( .A(n287), .B(n323), .CO(n221), .S(n222) );
  FA_X1 U192 ( .A(n324), .B(n288), .CI(n310), .CO(n225), .S(n226) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  HA_X1 U194 ( .A(n311), .B(n325), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n326), .B(n300), .CI(n312), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  XNOR2_X1 U414 ( .A(n506), .B(n490), .ZN(product[9]) );
  AND2_X1 U415 ( .A1(n129), .A2(n90), .ZN(n490) );
  INV_X1 U416 ( .A(n536), .ZN(n491) );
  XOR2_X1 U417 ( .A(n590), .B(a[10]), .Z(n537) );
  OR2_X1 U418 ( .A1(n176), .A2(n185), .ZN(n492) );
  OR2_X2 U419 ( .A1(n518), .A2(n508), .ZN(n514) );
  XNOR2_X1 U420 ( .A(n493), .B(n179), .ZN(n166) );
  XNOR2_X1 U421 ( .A(n170), .B(n172), .ZN(n493) );
  BUF_X1 U422 ( .A(n9), .Z(n571) );
  XOR2_X1 U423 ( .A(n177), .B(n168), .Z(n494) );
  XOR2_X1 U424 ( .A(n166), .B(n494), .Z(n164) );
  NAND2_X1 U425 ( .A1(n170), .A2(n172), .ZN(n495) );
  NAND2_X1 U426 ( .A1(n170), .A2(n179), .ZN(n496) );
  NAND2_X1 U427 ( .A1(n172), .A2(n179), .ZN(n497) );
  NAND3_X1 U428 ( .A1(n495), .A2(n496), .A3(n497), .ZN(n165) );
  NAND2_X1 U429 ( .A1(n177), .A2(n168), .ZN(n498) );
  NAND2_X1 U430 ( .A1(n177), .A2(n166), .ZN(n499) );
  NAND2_X1 U431 ( .A1(n168), .A2(n166), .ZN(n500) );
  NAND3_X1 U432 ( .A1(n498), .A2(n499), .A3(n500), .ZN(n163) );
  OR2_X1 U433 ( .A1(n517), .A2(n78), .ZN(n501) );
  OR2_X1 U434 ( .A1(n329), .A2(n258), .ZN(n502) );
  NOR2_X1 U435 ( .A1(n228), .A2(n231), .ZN(n105) );
  OR2_X1 U436 ( .A1(n539), .A2(n561), .ZN(n524) );
  CLKBUF_X1 U437 ( .A(n45), .Z(n503) );
  XNOR2_X1 U438 ( .A(n504), .B(n505), .ZN(n570) );
  XNOR2_X1 U439 ( .A(n265), .B(n144), .ZN(n504) );
  XNOR2_X1 U440 ( .A(n161), .B(n142), .ZN(n505) );
  CLKBUF_X1 U441 ( .A(n540), .Z(n506) );
  BUF_X2 U442 ( .A(n9), .Z(n507) );
  XNOR2_X1 U443 ( .A(n581), .B(a[4]), .ZN(n508) );
  INV_X1 U444 ( .A(n589), .ZN(n509) );
  XNOR2_X1 U445 ( .A(n88), .B(n510), .ZN(product[10]) );
  NAND2_X1 U446 ( .A1(n525), .A2(n86), .ZN(n510) );
  INV_X1 U447 ( .A(n25), .ZN(n511) );
  BUF_X1 U448 ( .A(n519), .Z(n512) );
  INV_X2 U449 ( .A(n586), .ZN(n547) );
  INV_X2 U450 ( .A(n7), .ZN(n581) );
  XNOR2_X1 U451 ( .A(n149), .B(n513), .ZN(n144) );
  XNOR2_X1 U452 ( .A(n271), .B(n146), .ZN(n513) );
  OR2_X1 U453 ( .A1(n518), .A2(n552), .ZN(n18) );
  AOI21_X2 U454 ( .B1(n566), .B2(n112), .A(n109), .ZN(n107) );
  INV_X2 U455 ( .A(n592), .ZN(n591) );
  CLKBUF_X1 U456 ( .A(n548), .Z(n515) );
  INV_X1 U457 ( .A(n561), .ZN(n516) );
  INV_X1 U458 ( .A(n561), .ZN(n21) );
  OR2_X1 U459 ( .A1(n539), .A2(n561), .ZN(n23) );
  NOR2_X1 U460 ( .A1(n164), .A2(n175), .ZN(n517) );
  NOR2_X1 U461 ( .A1(n164), .A2(n175), .ZN(n75) );
  XNOR2_X1 U462 ( .A(n582), .B(a[4]), .ZN(n518) );
  NOR2_X1 U463 ( .A1(n186), .A2(n195), .ZN(n519) );
  NOR2_X1 U464 ( .A1(n186), .A2(n195), .ZN(n82) );
  INV_X1 U465 ( .A(n547), .ZN(n520) );
  XOR2_X1 U466 ( .A(n586), .B(a[8]), .Z(n27) );
  INV_X1 U467 ( .A(n590), .ZN(n521) );
  INV_X1 U468 ( .A(n581), .ZN(n522) );
  INV_X1 U469 ( .A(n1), .ZN(n523) );
  INV_X1 U470 ( .A(n1), .ZN(n578) );
  OR2_X1 U471 ( .A1(n196), .A2(n203), .ZN(n525) );
  OAI21_X1 U472 ( .B1(n105), .B2(n107), .A(n106), .ZN(n526) );
  INV_X1 U473 ( .A(n511), .ZN(n527) );
  INV_X1 U474 ( .A(n588), .ZN(n528) );
  INV_X1 U475 ( .A(n588), .ZN(n587) );
  INV_X1 U476 ( .A(n590), .ZN(n529) );
  INV_X1 U477 ( .A(n590), .ZN(n589) );
  NAND2_X1 U478 ( .A1(n562), .A2(n541), .ZN(n530) );
  NAND2_X1 U479 ( .A1(n562), .A2(n541), .ZN(n550) );
  NOR2_X1 U480 ( .A1(n204), .A2(n211), .ZN(n531) );
  CLKBUF_X1 U481 ( .A(n29), .Z(n532) );
  XNOR2_X1 U482 ( .A(n521), .B(a[12]), .ZN(n533) );
  XNOR2_X1 U483 ( .A(n521), .B(a[12]), .ZN(n534) );
  XNOR2_X1 U484 ( .A(n589), .B(a[12]), .ZN(n37) );
  BUF_X2 U485 ( .A(n545), .Z(n535) );
  INV_X1 U486 ( .A(n584), .ZN(n536) );
  OR2_X2 U487 ( .A1(n537), .A2(n538), .ZN(n34) );
  XOR2_X1 U488 ( .A(n587), .B(a[10]), .Z(n538) );
  NAND2_X1 U489 ( .A1(n429), .A2(n27), .ZN(n29) );
  NOR2_X1 U490 ( .A1(n196), .A2(n203), .ZN(n85) );
  XNOR2_X1 U491 ( .A(n585), .B(a[6]), .ZN(n539) );
  AOI21_X1 U492 ( .B1(n96), .B2(n564), .A(n93), .ZN(n540) );
  INV_X2 U493 ( .A(n552), .ZN(n16) );
  XOR2_X1 U494 ( .A(n523), .B(a[2]), .Z(n541) );
  XNOR2_X1 U495 ( .A(n581), .B(a[2]), .ZN(n562) );
  INV_X1 U496 ( .A(n581), .ZN(n579) );
  AOI21_X1 U497 ( .B1(n96), .B2(n564), .A(n93), .ZN(n91) );
  INV_X1 U498 ( .A(n575), .ZN(n542) );
  INV_X1 U499 ( .A(n542), .ZN(n543) );
  INV_X2 U500 ( .A(n542), .ZN(n544) );
  XNOR2_X1 U501 ( .A(n25), .B(a[10]), .ZN(n545) );
  OAI21_X1 U502 ( .B1(n82), .B2(n86), .A(n83), .ZN(n546) );
  BUF_X2 U503 ( .A(n27), .Z(n548) );
  INV_X1 U504 ( .A(n586), .ZN(n585) );
  OAI21_X1 U505 ( .B1(n540), .B2(n531), .A(n90), .ZN(n549) );
  AOI21_X1 U506 ( .B1(n526), .B2(n572), .A(n101), .ZN(n551) );
  NAND2_X1 U507 ( .A1(n562), .A2(n541), .ZN(n12) );
  XNOR2_X1 U508 ( .A(n581), .B(a[4]), .ZN(n552) );
  XNOR2_X1 U509 ( .A(n523), .B(n249), .ZN(n433) );
  XOR2_X1 U510 ( .A(n229), .B(n298), .Z(n553) );
  XOR2_X1 U511 ( .A(n226), .B(n553), .Z(n224) );
  NAND2_X1 U512 ( .A1(n226), .A2(n229), .ZN(n554) );
  NAND2_X1 U513 ( .A1(n226), .A2(n298), .ZN(n555) );
  NAND2_X1 U514 ( .A1(n229), .A2(n298), .ZN(n556) );
  NAND3_X1 U515 ( .A1(n554), .A2(n555), .A3(n556), .ZN(n223) );
  XOR2_X1 U516 ( .A(n578), .B(a[2]), .Z(n9) );
  OAI21_X1 U517 ( .B1(n551), .B2(n97), .A(n98), .ZN(n557) );
  NAND2_X1 U518 ( .A1(n433), .A2(n543), .ZN(n558) );
  NAND2_X1 U519 ( .A1(n433), .A2(n543), .ZN(n559) );
  AOI21_X1 U520 ( .B1(n80), .B2(n549), .A(n81), .ZN(n560) );
  XNOR2_X1 U521 ( .A(n584), .B(a[6]), .ZN(n561) );
  BUF_X1 U522 ( .A(n43), .Z(n573) );
  XNOR2_X1 U523 ( .A(n70), .B(n47), .ZN(product[14]) );
  NAND2_X1 U524 ( .A1(n563), .A2(n69), .ZN(n47) );
  INV_X1 U525 ( .A(n74), .ZN(n72) );
  AOI21_X1 U526 ( .B1(n563), .B2(n74), .A(n67), .ZN(n65) );
  INV_X1 U527 ( .A(n69), .ZN(n67) );
  NAND2_X1 U528 ( .A1(n73), .A2(n563), .ZN(n64) );
  INV_X1 U529 ( .A(n95), .ZN(n93) );
  AOI21_X1 U530 ( .B1(n80), .B2(n549), .A(n546), .ZN(n45) );
  NOR2_X1 U531 ( .A1(n82), .A2(n85), .ZN(n80) );
  OAI21_X1 U532 ( .B1(n519), .B2(n86), .A(n83), .ZN(n81) );
  NAND2_X1 U533 ( .A1(n492), .A2(n79), .ZN(n49) );
  NAND2_X1 U534 ( .A1(n125), .A2(n76), .ZN(n48) );
  INV_X1 U535 ( .A(n517), .ZN(n125) );
  INV_X1 U536 ( .A(n531), .ZN(n129) );
  OR2_X1 U537 ( .A1(n152), .A2(n163), .ZN(n563) );
  OAI21_X1 U538 ( .B1(n91), .B2(n89), .A(n90), .ZN(n88) );
  OAI21_X1 U539 ( .B1(n75), .B2(n79), .A(n76), .ZN(n74) );
  NAND2_X1 U540 ( .A1(n127), .A2(n83), .ZN(n50) );
  INV_X1 U541 ( .A(n512), .ZN(n127) );
  NOR2_X1 U542 ( .A1(n517), .A2(n78), .ZN(n73) );
  XNOR2_X1 U543 ( .A(n557), .B(n53), .ZN(product[8]) );
  NAND2_X1 U544 ( .A1(n564), .A2(n95), .ZN(n53) );
  NAND2_X1 U545 ( .A1(n152), .A2(n163), .ZN(n69) );
  AOI21_X1 U546 ( .B1(n104), .B2(n572), .A(n101), .ZN(n99) );
  OAI21_X1 U547 ( .B1(n113), .B2(n115), .A(n114), .ZN(n112) );
  NAND2_X1 U548 ( .A1(n133), .A2(n106), .ZN(n56) );
  INV_X1 U549 ( .A(n105), .ZN(n133) );
  OAI21_X1 U550 ( .B1(n99), .B2(n97), .A(n98), .ZN(n96) );
  NOR2_X1 U551 ( .A1(n176), .A2(n185), .ZN(n78) );
  AOI21_X1 U552 ( .B1(n565), .B2(n120), .A(n117), .ZN(n115) );
  INV_X1 U553 ( .A(n119), .ZN(n117) );
  XOR2_X1 U554 ( .A(n54), .B(n551), .Z(product[7]) );
  NAND2_X1 U555 ( .A1(n131), .A2(n98), .ZN(n54) );
  INV_X1 U556 ( .A(n97), .ZN(n131) );
  XNOR2_X1 U557 ( .A(n57), .B(n112), .ZN(product[4]) );
  NAND2_X1 U558 ( .A1(n566), .A2(n111), .ZN(n57) );
  XNOR2_X1 U559 ( .A(n59), .B(n120), .ZN(product[2]) );
  NAND2_X1 U560 ( .A1(n565), .A2(n119), .ZN(n59) );
  NAND2_X1 U561 ( .A1(n176), .A2(n185), .ZN(n79) );
  NAND2_X1 U562 ( .A1(n186), .A2(n195), .ZN(n83) );
  NAND2_X1 U563 ( .A1(n164), .A2(n175), .ZN(n76) );
  NAND2_X1 U564 ( .A1(n196), .A2(n203), .ZN(n86) );
  NAND2_X1 U565 ( .A1(n212), .A2(n217), .ZN(n95) );
  NAND2_X1 U566 ( .A1(n204), .A2(n211), .ZN(n90) );
  OR2_X1 U567 ( .A1(n212), .A2(n217), .ZN(n564) );
  NAND2_X1 U568 ( .A1(n135), .A2(n114), .ZN(n58) );
  INV_X1 U569 ( .A(n113), .ZN(n135) );
  NOR2_X1 U570 ( .A1(n218), .A2(n223), .ZN(n97) );
  OR2_X1 U571 ( .A1(n328), .A2(n314), .ZN(n565) );
  XNOR2_X1 U572 ( .A(n63), .B(n46), .ZN(product[15]) );
  NAND2_X1 U573 ( .A1(n567), .A2(n62), .ZN(n46) );
  NAND2_X1 U574 ( .A1(n218), .A2(n223), .ZN(n98) );
  OR2_X1 U575 ( .A1(n232), .A2(n233), .ZN(n566) );
  INV_X1 U576 ( .A(n533), .ZN(n237) );
  NAND2_X1 U577 ( .A1(n232), .A2(n233), .ZN(n111) );
  INV_X1 U578 ( .A(n41), .ZN(n235) );
  OR2_X1 U579 ( .A1(n151), .A2(n139), .ZN(n567) );
  OR2_X1 U580 ( .A1(n224), .A2(n227), .ZN(n572) );
  AND2_X1 U581 ( .A1(n502), .A2(n122), .ZN(product[1]) );
  INV_X1 U582 ( .A(n249), .ZN(n575) );
  XNOR2_X1 U583 ( .A(n591), .B(a[14]), .ZN(n41) );
  OR2_X1 U584 ( .A1(n573), .A2(n581), .ZN(n392) );
  NAND2_X1 U585 ( .A1(n433), .A2(n543), .ZN(n6) );
  AND2_X1 U586 ( .A1(n574), .A2(n508), .ZN(n300) );
  OAI22_X1 U587 ( .A1(n559), .A2(n405), .B1(n404), .B2(n544), .ZN(n326) );
  OAI22_X1 U588 ( .A1(n6), .A2(n400), .B1(n399), .B2(n544), .ZN(n321) );
  XNOR2_X1 U589 ( .A(n528), .B(n573), .ZN(n352) );
  OAI22_X1 U590 ( .A1(n559), .A2(n406), .B1(n405), .B2(n544), .ZN(n327) );
  XNOR2_X1 U591 ( .A(n155), .B(n569), .ZN(n139) );
  XNOR2_X1 U592 ( .A(n153), .B(n141), .ZN(n569) );
  XNOR2_X1 U593 ( .A(n157), .B(n570), .ZN(n141) );
  OAI22_X1 U594 ( .A1(n6), .A2(n408), .B1(n407), .B2(n544), .ZN(n329) );
  OAI22_X1 U595 ( .A1(n558), .A2(n398), .B1(n397), .B2(n544), .ZN(n319) );
  OAI22_X1 U596 ( .A1(n34), .A2(n343), .B1(n342), .B2(n535), .ZN(n269) );
  XNOR2_X1 U597 ( .A(n529), .B(n573), .ZN(n343) );
  OAI22_X1 U598 ( .A1(n42), .A2(n594), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U599 ( .A1(n573), .A2(n594), .ZN(n332) );
  OAI22_X1 U600 ( .A1(n558), .A2(n404), .B1(n403), .B2(n544), .ZN(n325) );
  XOR2_X1 U601 ( .A(n587), .B(a[8]), .Z(n429) );
  XOR2_X1 U602 ( .A(n315), .B(n261), .Z(n150) );
  OAI22_X1 U603 ( .A1(n6), .A2(n394), .B1(n393), .B2(n544), .ZN(n315) );
  XNOR2_X1 U604 ( .A(n591), .B(n573), .ZN(n336) );
  NAND2_X1 U605 ( .A1(n427), .A2(n37), .ZN(n39) );
  XOR2_X1 U606 ( .A(n591), .B(a[12]), .Z(n427) );
  AND2_X1 U607 ( .A1(n574), .A2(n241), .ZN(n278) );
  OAI22_X1 U608 ( .A1(n559), .A2(n401), .B1(n400), .B2(n544), .ZN(n322) );
  OAI22_X1 U609 ( .A1(n34), .A2(n342), .B1(n341), .B2(n535), .ZN(n268) );
  OAI22_X1 U610 ( .A1(n34), .A2(n341), .B1(n340), .B2(n535), .ZN(n267) );
  OAI22_X1 U611 ( .A1(n6), .A2(n397), .B1(n396), .B2(n544), .ZN(n318) );
  AND2_X1 U612 ( .A1(n574), .A2(n237), .ZN(n264) );
  OAI22_X1 U613 ( .A1(n39), .A2(n336), .B1(n534), .B2(n335), .ZN(n263) );
  XNOR2_X1 U614 ( .A(n583), .B(n573), .ZN(n376) );
  AND2_X1 U615 ( .A1(n574), .A2(n561), .ZN(n288) );
  OAI22_X1 U616 ( .A1(n6), .A2(n403), .B1(n402), .B2(n544), .ZN(n324) );
  AND2_X1 U617 ( .A1(n574), .A2(n538), .ZN(n270) );
  OAI22_X1 U618 ( .A1(n559), .A2(n399), .B1(n398), .B2(n544), .ZN(n320) );
  OAI22_X1 U619 ( .A1(n34), .A2(n509), .B1(n344), .B2(n535), .ZN(n253) );
  AND2_X1 U620 ( .A1(n574), .A2(n235), .ZN(n260) );
  OAI22_X1 U621 ( .A1(n559), .A2(n395), .B1(n394), .B2(n544), .ZN(n316) );
  OAI22_X1 U622 ( .A1(n39), .A2(n335), .B1(n533), .B2(n334), .ZN(n262) );
  INV_X1 U623 ( .A(n19), .ZN(n586) );
  INV_X1 U624 ( .A(n25), .ZN(n588) );
  OAI22_X1 U625 ( .A1(n34), .A2(n340), .B1(n339), .B2(n535), .ZN(n266) );
  NAND2_X1 U626 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U627 ( .A(n593), .B(a[14]), .Z(n426) );
  INV_X1 U628 ( .A(n13), .ZN(n584) );
  OAI22_X1 U629 ( .A1(n6), .A2(n402), .B1(n401), .B2(n544), .ZN(n323) );
  XNOR2_X1 U630 ( .A(n547), .B(n573), .ZN(n363) );
  OAI22_X1 U631 ( .A1(n558), .A2(n396), .B1(n395), .B2(n544), .ZN(n317) );
  OAI22_X1 U632 ( .A1(n39), .A2(n592), .B1(n337), .B2(n533), .ZN(n252) );
  OR2_X1 U633 ( .A1(n573), .A2(n592), .ZN(n337) );
  AND2_X1 U634 ( .A1(n574), .A2(n247), .ZN(n314) );
  OR2_X1 U635 ( .A1(n573), .A2(n509), .ZN(n344) );
  AND2_X1 U636 ( .A1(n574), .A2(n249), .ZN(product[0]) );
  OR2_X1 U637 ( .A1(n573), .A2(n520), .ZN(n364) );
  OR2_X1 U638 ( .A1(n573), .A2(n511), .ZN(n353) );
  OR2_X1 U639 ( .A1(n573), .A2(n491), .ZN(n377) );
  XNOR2_X1 U640 ( .A(n547), .B(b[9]), .ZN(n354) );
  OAI22_X1 U641 ( .A1(n39), .A2(n334), .B1(n534), .B2(n333), .ZN(n261) );
  XNOR2_X1 U642 ( .A(n591), .B(n422), .ZN(n333) );
  XNOR2_X1 U643 ( .A(n583), .B(b[11]), .ZN(n365) );
  XNOR2_X1 U644 ( .A(n521), .B(n424), .ZN(n342) );
  XNOR2_X1 U645 ( .A(n529), .B(n423), .ZN(n341) );
  XNOR2_X1 U646 ( .A(n529), .B(n422), .ZN(n340) );
  XNOR2_X1 U647 ( .A(n529), .B(n421), .ZN(n339) );
  XNOR2_X1 U648 ( .A(n591), .B(n424), .ZN(n335) );
  XNOR2_X1 U649 ( .A(n591), .B(n423), .ZN(n334) );
  OAI22_X1 U650 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U651 ( .A(n593), .B(n424), .ZN(n330) );
  XNOR2_X1 U652 ( .A(n593), .B(n573), .ZN(n331) );
  XNOR2_X1 U653 ( .A(n577), .B(b[11]), .ZN(n397) );
  XNOR2_X1 U654 ( .A(n577), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U655 ( .A(n577), .B(b[13]), .ZN(n395) );
  XNOR2_X1 U656 ( .A(n577), .B(b[14]), .ZN(n394) );
  XNOR2_X1 U657 ( .A(n527), .B(n418), .ZN(n345) );
  OAI22_X1 U658 ( .A1(n34), .A2(n339), .B1(n338), .B2(n535), .ZN(n265) );
  XNOR2_X1 U659 ( .A(n529), .B(n420), .ZN(n338) );
  XNOR2_X1 U660 ( .A(n522), .B(b[13]), .ZN(n378) );
  XNOR2_X1 U661 ( .A(n547), .B(n424), .ZN(n362) );
  XNOR2_X1 U662 ( .A(n528), .B(n424), .ZN(n351) );
  XNOR2_X1 U663 ( .A(n580), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U664 ( .A(n580), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U665 ( .A(n580), .B(n418), .ZN(n384) );
  XNOR2_X1 U666 ( .A(n522), .B(n419), .ZN(n385) );
  XNOR2_X1 U667 ( .A(n522), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U668 ( .A(n580), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U669 ( .A(n522), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U670 ( .A(n583), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U671 ( .A(n583), .B(n418), .ZN(n369) );
  XNOR2_X1 U672 ( .A(n583), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U673 ( .A(n583), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U674 ( .A(n547), .B(n423), .ZN(n361) );
  XNOR2_X1 U675 ( .A(n547), .B(n422), .ZN(n360) );
  XNOR2_X1 U676 ( .A(n527), .B(n423), .ZN(n350) );
  XNOR2_X1 U677 ( .A(n527), .B(n422), .ZN(n349) );
  XNOR2_X1 U678 ( .A(n547), .B(n421), .ZN(n359) );
  XNOR2_X1 U679 ( .A(n527), .B(n421), .ZN(n348) );
  XNOR2_X1 U680 ( .A(n547), .B(n420), .ZN(n358) );
  XNOR2_X1 U681 ( .A(n528), .B(n420), .ZN(n347) );
  XNOR2_X1 U682 ( .A(n547), .B(n419), .ZN(n357) );
  XNOR2_X1 U683 ( .A(n528), .B(n419), .ZN(n346) );
  XNOR2_X1 U684 ( .A(n547), .B(n418), .ZN(n356) );
  XNOR2_X1 U685 ( .A(n547), .B(b[8]), .ZN(n355) );
  XNOR2_X1 U686 ( .A(n577), .B(b[15]), .ZN(n393) );
  BUF_X1 U687 ( .A(n43), .Z(n574) );
  NAND2_X1 U688 ( .A1(n328), .A2(n314), .ZN(n119) );
  OAI22_X1 U689 ( .A1(n558), .A2(n407), .B1(n406), .B2(n544), .ZN(n328) );
  NAND2_X1 U690 ( .A1(n228), .A2(n231), .ZN(n106) );
  NAND2_X1 U691 ( .A1(n572), .A2(n103), .ZN(n55) );
  INV_X1 U692 ( .A(n103), .ZN(n101) );
  NAND2_X1 U693 ( .A1(n224), .A2(n227), .ZN(n103) );
  XNOR2_X1 U694 ( .A(n55), .B(n526), .ZN(product[6]) );
  OAI21_X1 U695 ( .B1(n105), .B2(n107), .A(n106), .ZN(n104) );
  NOR2_X1 U696 ( .A1(n234), .A2(n257), .ZN(n113) );
  XOR2_X1 U697 ( .A(n58), .B(n115), .Z(product[3]) );
  NAND2_X1 U698 ( .A1(n151), .A2(n139), .ZN(n62) );
  NOR2_X1 U699 ( .A1(n204), .A2(n211), .ZN(n89) );
  OAI22_X1 U700 ( .A1(n532), .A2(n350), .B1(n349), .B2(n515), .ZN(n275) );
  OAI22_X1 U701 ( .A1(n29), .A2(n348), .B1(n347), .B2(n548), .ZN(n273) );
  OAI22_X1 U702 ( .A1(n29), .A2(n349), .B1(n348), .B2(n548), .ZN(n274) );
  OAI22_X1 U703 ( .A1(n29), .A2(n511), .B1(n353), .B2(n548), .ZN(n254) );
  OAI22_X1 U704 ( .A1(n29), .A2(n351), .B1(n350), .B2(n548), .ZN(n276) );
  OAI22_X1 U705 ( .A1(n532), .A2(n346), .B1(n345), .B2(n515), .ZN(n271) );
  OAI22_X1 U706 ( .A1(n532), .A2(n347), .B1(n346), .B2(n515), .ZN(n272) );
  INV_X1 U707 ( .A(n548), .ZN(n241) );
  OAI22_X1 U708 ( .A1(n29), .A2(n352), .B1(n351), .B2(n548), .ZN(n277) );
  OAI21_X1 U709 ( .B1(n87), .B2(n85), .A(n86), .ZN(n84) );
  INV_X1 U710 ( .A(n88), .ZN(n87) );
  XNOR2_X1 U711 ( .A(n77), .B(n48), .ZN(product[13]) );
  OAI22_X1 U712 ( .A1(n23), .A2(n358), .B1(n357), .B2(n516), .ZN(n282) );
  OAI22_X1 U713 ( .A1(n23), .A2(n356), .B1(n355), .B2(n516), .ZN(n280) );
  OAI22_X1 U714 ( .A1(n23), .A2(n362), .B1(n361), .B2(n516), .ZN(n286) );
  OAI22_X1 U715 ( .A1(n23), .A2(n360), .B1(n359), .B2(n516), .ZN(n284) );
  OAI22_X1 U716 ( .A1(n524), .A2(n361), .B1(n360), .B2(n21), .ZN(n285) );
  OAI22_X1 U717 ( .A1(n23), .A2(n520), .B1(n364), .B2(n21), .ZN(n255) );
  OAI22_X1 U718 ( .A1(n23), .A2(n357), .B1(n356), .B2(n516), .ZN(n281) );
  OAI22_X1 U719 ( .A1(n524), .A2(n359), .B1(n358), .B2(n21), .ZN(n283) );
  XNOR2_X1 U720 ( .A(n536), .B(n424), .ZN(n375) );
  OAI22_X1 U721 ( .A1(n524), .A2(n363), .B1(n21), .B2(n362), .ZN(n287) );
  XNOR2_X1 U722 ( .A(n536), .B(n423), .ZN(n374) );
  OAI22_X1 U723 ( .A1(n23), .A2(n355), .B1(n354), .B2(n21), .ZN(n279) );
  XNOR2_X1 U724 ( .A(n582), .B(n422), .ZN(n373) );
  XNOR2_X1 U725 ( .A(n582), .B(n421), .ZN(n372) );
  XNOR2_X1 U726 ( .A(n536), .B(n419), .ZN(n370) );
  XNOR2_X1 U727 ( .A(n582), .B(n420), .ZN(n371) );
  XNOR2_X1 U728 ( .A(n576), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U729 ( .A(n576), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U730 ( .A(n576), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U731 ( .A(n576), .B(n418), .ZN(n401) );
  XNOR2_X1 U732 ( .A(n576), .B(n421), .ZN(n404) );
  XNOR2_X1 U733 ( .A(n576), .B(n422), .ZN(n405) );
  XNOR2_X1 U734 ( .A(n576), .B(n420), .ZN(n403) );
  XNOR2_X1 U735 ( .A(n576), .B(n419), .ZN(n402) );
  XNOR2_X1 U736 ( .A(n576), .B(n573), .ZN(n408) );
  XNOR2_X1 U737 ( .A(n576), .B(n423), .ZN(n406) );
  XNOR2_X1 U738 ( .A(n576), .B(n424), .ZN(n407) );
  INV_X1 U739 ( .A(n523), .ZN(n577) );
  OR2_X1 U740 ( .A1(n573), .A2(n523), .ZN(n409) );
  INV_X2 U741 ( .A(n578), .ZN(n576) );
  OAI22_X1 U742 ( .A1(n514), .A2(n370), .B1(n369), .B2(n16), .ZN(n293) );
  OAI22_X1 U743 ( .A1(n514), .A2(n367), .B1(n366), .B2(n16), .ZN(n290) );
  OAI22_X1 U744 ( .A1(n514), .A2(n375), .B1(n374), .B2(n16), .ZN(n298) );
  OAI22_X1 U745 ( .A1(n514), .A2(n373), .B1(n372), .B2(n16), .ZN(n296) );
  OAI22_X1 U746 ( .A1(n514), .A2(n376), .B1(n375), .B2(n16), .ZN(n299) );
  OAI22_X1 U747 ( .A1(n514), .A2(n491), .B1(n377), .B2(n16), .ZN(n256) );
  OAI22_X1 U748 ( .A1(n18), .A2(n372), .B1(n371), .B2(n16), .ZN(n295) );
  OAI22_X1 U749 ( .A1(n514), .A2(n368), .B1(n367), .B2(n16), .ZN(n291) );
  OAI22_X1 U750 ( .A1(n18), .A2(n369), .B1(n368), .B2(n16), .ZN(n292) );
  OAI22_X1 U751 ( .A1(n18), .A2(n371), .B1(n370), .B2(n16), .ZN(n294) );
  OAI22_X1 U752 ( .A1(n18), .A2(n374), .B1(n373), .B2(n16), .ZN(n297) );
  OAI22_X1 U753 ( .A1(n514), .A2(n366), .B1(n365), .B2(n16), .ZN(n289) );
  XNOR2_X1 U754 ( .A(n579), .B(n420), .ZN(n386) );
  XNOR2_X1 U755 ( .A(n579), .B(n573), .ZN(n391) );
  XNOR2_X1 U756 ( .A(n579), .B(n424), .ZN(n390) );
  XNOR2_X1 U757 ( .A(n579), .B(n422), .ZN(n388) );
  XNOR2_X1 U758 ( .A(n579), .B(n423), .ZN(n389) );
  XNOR2_X1 U759 ( .A(n579), .B(n421), .ZN(n387) );
  XNOR2_X1 U760 ( .A(n84), .B(n50), .ZN(product[11]) );
  OAI21_X1 U761 ( .B1(n64), .B2(n503), .A(n65), .ZN(n63) );
  OAI21_X1 U762 ( .B1(n560), .B2(n78), .A(n79), .ZN(n77) );
  OAI21_X1 U763 ( .B1(n501), .B2(n560), .A(n72), .ZN(n70) );
  XOR2_X1 U764 ( .A(n45), .B(n49), .Z(product[12]) );
  XOR2_X1 U765 ( .A(n56), .B(n107), .Z(product[5]) );
  INV_X1 U766 ( .A(n122), .ZN(n120) );
  NAND2_X1 U767 ( .A1(n329), .A2(n258), .ZN(n122) );
  INV_X1 U768 ( .A(n111), .ZN(n109) );
  OAI22_X1 U769 ( .A1(n558), .A2(n578), .B1(n409), .B2(n544), .ZN(n258) );
  OAI22_X1 U770 ( .A1(n12), .A2(n379), .B1(n378), .B2(n507), .ZN(n301) );
  OAI22_X1 U771 ( .A1(n530), .A2(n380), .B1(n379), .B2(n507), .ZN(n302) );
  OAI22_X1 U772 ( .A1(n12), .A2(n385), .B1(n384), .B2(n507), .ZN(n307) );
  OAI22_X1 U773 ( .A1(n12), .A2(n382), .B1(n381), .B2(n507), .ZN(n304) );
  OAI22_X1 U774 ( .A1(n12), .A2(n381), .B1(n380), .B2(n507), .ZN(n303) );
  NAND2_X1 U775 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U776 ( .A1(n550), .A2(n383), .B1(n382), .B2(n571), .ZN(n305) );
  OAI22_X1 U777 ( .A1(n550), .A2(n384), .B1(n383), .B2(n571), .ZN(n306) );
  OAI22_X1 U778 ( .A1(n530), .A2(n386), .B1(n385), .B2(n507), .ZN(n308) );
  OAI22_X1 U779 ( .A1(n530), .A2(n387), .B1(n386), .B2(n507), .ZN(n309) );
  OAI22_X1 U780 ( .A1(n530), .A2(n581), .B1(n392), .B2(n571), .ZN(n257) );
  OAI22_X1 U781 ( .A1(n389), .A2(n550), .B1(n388), .B2(n9), .ZN(n311) );
  OAI22_X1 U782 ( .A1(n388), .A2(n12), .B1(n387), .B2(n507), .ZN(n310) );
  OAI22_X1 U783 ( .A1(n530), .A2(n390), .B1(n389), .B2(n507), .ZN(n312) );
  INV_X1 U784 ( .A(n507), .ZN(n247) );
  OAI22_X1 U785 ( .A1(n530), .A2(n391), .B1(n390), .B2(n507), .ZN(n313) );
  INV_X1 U786 ( .A(n581), .ZN(n580) );
  INV_X1 U787 ( .A(n584), .ZN(n582) );
  INV_X1 U788 ( .A(n584), .ZN(n583) );
  INV_X1 U789 ( .A(n31), .ZN(n590) );
  INV_X1 U790 ( .A(n36), .ZN(n592) );
  INV_X1 U791 ( .A(n594), .ZN(n593) );
  INV_X1 U792 ( .A(n40), .ZN(n594) );
  XOR2_X1 U793 ( .A(n259), .B(n251), .Z(n148) );
  XOR2_X1 U794 ( .A(n289), .B(n279), .Z(n146) );
  XOR2_X1 U795 ( .A(n159), .B(n150), .Z(n142) );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_3_DW01_add_2 ( A, B, CI, 
        SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n5, n8, n9, n10, n11, n12, n13, n14, n15, n16, n19, n20, n22,
         n24, n25, n26, n27, n28, n29, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n42, n44, n45, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n65, n67, n68, n69, n70, n71, n73, n75,
         n76, n77, n78, n79, n81, n83, n84, n86, n88, n90, n91, n94, n95, n96,
         n98, n100, n157, n158, n159, n160, n161, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180;

  NOR2_X1 U122 ( .A1(A[8]), .A2(B[8]), .ZN(n157) );
  NOR2_X1 U123 ( .A1(A[8]), .A2(B[8]), .ZN(n158) );
  NOR2_X1 U124 ( .A1(A[8]), .A2(B[8]), .ZN(n54) );
  AOI21_X1 U125 ( .B1(n52), .B2(n60), .A(n53), .ZN(n159) );
  INV_X1 U126 ( .A(n91), .ZN(n160) );
  XNOR2_X1 U127 ( .A(n37), .B(n161), .ZN(SUM[11]) );
  AND2_X1 U128 ( .A1(n91), .A2(n36), .ZN(n161) );
  AND2_X1 U129 ( .A1(n174), .A2(n86), .ZN(SUM[0]) );
  OR2_X1 U130 ( .A1(A[15]), .A2(B[15]), .ZN(n163) );
  XNOR2_X1 U131 ( .A(n45), .B(n164), .ZN(SUM[10]) );
  AND2_X1 U132 ( .A1(n177), .A2(n44), .ZN(n164) );
  NOR2_X1 U133 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  CLKBUF_X1 U134 ( .A(n171), .Z(n165) );
  NOR2_X1 U135 ( .A1(A[12]), .A2(B[12]), .ZN(n171) );
  AND2_X1 U136 ( .A1(A[9]), .A2(B[9]), .ZN(n166) );
  OR2_X1 U137 ( .A1(A[13]), .A2(B[13]), .ZN(n167) );
  XNOR2_X1 U138 ( .A(n173), .B(n168), .ZN(SUM[13]) );
  AND2_X1 U139 ( .A1(n167), .A2(n29), .ZN(n168) );
  NOR2_X1 U140 ( .A1(n171), .A2(n35), .ZN(n169) );
  NOR2_X1 U141 ( .A1(A[14]), .A2(B[14]), .ZN(n170) );
  AOI21_X1 U142 ( .B1(n38), .B2(n169), .A(n31), .ZN(n172) );
  AOI21_X1 U143 ( .B1(n38), .B2(n169), .A(n31), .ZN(n173) );
  OR2_X1 U144 ( .A1(A[0]), .A2(B[0]), .ZN(n174) );
  INV_X1 U145 ( .A(n60), .ZN(n59) );
  INV_X1 U146 ( .A(n159), .ZN(n50) );
  INV_X1 U147 ( .A(n38), .ZN(n37) );
  AOI21_X1 U148 ( .B1(n52), .B2(n60), .A(n53), .ZN(n51) );
  INV_X1 U149 ( .A(n67), .ZN(n65) );
  AOI21_X1 U150 ( .B1(n176), .B2(n84), .A(n81), .ZN(n79) );
  INV_X1 U151 ( .A(n83), .ZN(n81) );
  OAI21_X1 U152 ( .B1(n79), .B2(n77), .A(n78), .ZN(n76) );
  AOI21_X1 U153 ( .B1(n175), .B2(n76), .A(n73), .ZN(n71) );
  INV_X1 U154 ( .A(n75), .ZN(n73) );
  AOI21_X1 U155 ( .B1(n50), .B2(n178), .A(n166), .ZN(n45) );
  NAND2_X1 U156 ( .A1(n94), .A2(n55), .ZN(n9) );
  INV_X1 U157 ( .A(n86), .ZN(n84) );
  OAI21_X1 U158 ( .B1(n59), .B2(n57), .A(n58), .ZN(n56) );
  NAND2_X1 U159 ( .A1(n95), .A2(n58), .ZN(n10) );
  INV_X1 U160 ( .A(n57), .ZN(n95) );
  NAND2_X1 U161 ( .A1(n179), .A2(n67), .ZN(n12) );
  NAND2_X1 U162 ( .A1(n100), .A2(n78), .ZN(n15) );
  INV_X1 U163 ( .A(n77), .ZN(n100) );
  NAND2_X1 U164 ( .A1(n98), .A2(n70), .ZN(n13) );
  INV_X1 U165 ( .A(n69), .ZN(n98) );
  NAND2_X1 U166 ( .A1(n176), .A2(n83), .ZN(n16) );
  NAND2_X1 U167 ( .A1(n175), .A2(n75), .ZN(n14) );
  NAND2_X1 U168 ( .A1(n96), .A2(n62), .ZN(n11) );
  INV_X1 U169 ( .A(n61), .ZN(n96) );
  XOR2_X1 U170 ( .A(n13), .B(n71), .Z(SUM[4]) );
  XOR2_X1 U171 ( .A(n15), .B(n79), .Z(SUM[2]) );
  NAND2_X1 U172 ( .A1(n88), .A2(n26), .ZN(n3) );
  NOR2_X1 U173 ( .A1(A[7]), .A2(B[7]), .ZN(n57) );
  NOR2_X1 U174 ( .A1(A[12]), .A2(B[12]), .ZN(n32) );
  NOR2_X1 U175 ( .A1(A[14]), .A2(B[14]), .ZN(n25) );
  NOR2_X1 U176 ( .A1(A[2]), .A2(B[2]), .ZN(n77) );
  NAND2_X1 U177 ( .A1(n90), .A2(n33), .ZN(n5) );
  NAND2_X1 U178 ( .A1(A[13]), .A2(B[13]), .ZN(n29) );
  OR2_X1 U179 ( .A1(A[3]), .A2(B[3]), .ZN(n175) );
  OR2_X1 U180 ( .A1(A[1]), .A2(B[1]), .ZN(n176) );
  OR2_X1 U181 ( .A1(A[10]), .A2(B[10]), .ZN(n177) );
  NAND2_X1 U182 ( .A1(n163), .A2(n19), .ZN(n2) );
  OR2_X1 U183 ( .A1(A[9]), .A2(B[9]), .ZN(n178) );
  NAND2_X1 U184 ( .A1(A[14]), .A2(B[14]), .ZN(n26) );
  XNOR2_X1 U185 ( .A(n56), .B(n9), .ZN(SUM[8]) );
  XNOR2_X1 U186 ( .A(n14), .B(n76), .ZN(SUM[3]) );
  NOR2_X1 U187 ( .A1(A[4]), .A2(B[4]), .ZN(n69) );
  NOR2_X1 U188 ( .A1(A[6]), .A2(B[6]), .ZN(n61) );
  NAND2_X1 U189 ( .A1(A[7]), .A2(B[7]), .ZN(n58) );
  NAND2_X1 U190 ( .A1(A[2]), .A2(B[2]), .ZN(n78) );
  NAND2_X1 U191 ( .A1(A[1]), .A2(B[1]), .ZN(n83) );
  NAND2_X1 U192 ( .A1(A[0]), .A2(B[0]), .ZN(n86) );
  NAND2_X1 U193 ( .A1(A[4]), .A2(B[4]), .ZN(n70) );
  NAND2_X1 U194 ( .A1(A[6]), .A2(B[6]), .ZN(n62) );
  OR2_X1 U195 ( .A1(A[5]), .A2(B[5]), .ZN(n179) );
  NAND2_X1 U196 ( .A1(A[3]), .A2(B[3]), .ZN(n75) );
  NAND2_X1 U197 ( .A1(A[12]), .A2(B[12]), .ZN(n33) );
  NAND2_X1 U198 ( .A1(A[9]), .A2(B[9]), .ZN(n49) );
  XNOR2_X1 U199 ( .A(n50), .B(n8), .ZN(SUM[9]) );
  XOR2_X1 U200 ( .A(n59), .B(n10), .Z(SUM[7]) );
  XNOR2_X1 U201 ( .A(n16), .B(n84), .ZN(SUM[1]) );
  NAND2_X1 U202 ( .A1(A[5]), .A2(B[5]), .ZN(n67) );
  OR2_X1 U203 ( .A1(n25), .A2(n28), .ZN(n180) );
  NAND2_X1 U204 ( .A1(n178), .A2(n49), .ZN(n8) );
  INV_X1 U205 ( .A(n158), .ZN(n94) );
  NOR2_X1 U206 ( .A1(n157), .A2(n57), .ZN(n52) );
  OAI21_X1 U207 ( .B1(n54), .B2(n58), .A(n55), .ZN(n53) );
  NAND2_X1 U208 ( .A1(A[8]), .A2(B[8]), .ZN(n55) );
  XOR2_X1 U209 ( .A(n11), .B(n63), .Z(SUM[6]) );
  OAI21_X1 U210 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  AOI21_X1 U211 ( .B1(n179), .B2(n68), .A(n65), .ZN(n63) );
  XNOR2_X1 U212 ( .A(n12), .B(n68), .ZN(SUM[5]) );
  NAND2_X1 U213 ( .A1(A[11]), .A2(B[11]), .ZN(n36) );
  INV_X1 U214 ( .A(n24), .ZN(n22) );
  INV_X1 U215 ( .A(n25), .ZN(n88) );
  OAI21_X1 U216 ( .B1(n170), .B2(n29), .A(n26), .ZN(n24) );
  OAI21_X1 U217 ( .B1(n71), .B2(n69), .A(n70), .ZN(n68) );
  INV_X1 U218 ( .A(n44), .ZN(n42) );
  INV_X1 U219 ( .A(n165), .ZN(n90) );
  OAI21_X1 U220 ( .B1(n32), .B2(n36), .A(n33), .ZN(n31) );
  NAND2_X1 U221 ( .A1(A[15]), .A2(B[15]), .ZN(n19) );
  XNOR2_X1 U222 ( .A(n27), .B(n3), .ZN(SUM[14]) );
  INV_X1 U223 ( .A(n35), .ZN(n91) );
  OAI21_X1 U224 ( .B1(n37), .B2(n160), .A(n36), .ZN(n34) );
  NOR2_X1 U225 ( .A1(A[11]), .A2(B[11]), .ZN(n35) );
  NAND2_X1 U226 ( .A1(n177), .A2(n178), .ZN(n39) );
  AOI21_X1 U227 ( .B1(n177), .B2(n166), .A(n42), .ZN(n40) );
  XNOR2_X1 U228 ( .A(n34), .B(n5), .ZN(SUM[12]) );
  XNOR2_X1 U229 ( .A(n20), .B(n2), .ZN(SUM[15]) );
  OAI21_X1 U230 ( .B1(n172), .B2(n28), .A(n29), .ZN(n27) );
  NAND2_X1 U231 ( .A1(A[10]), .A2(B[10]), .ZN(n44) );
  OAI21_X1 U232 ( .B1(n173), .B2(n180), .A(n22), .ZN(n20) );
  OAI21_X1 U233 ( .B1(n39), .B2(n51), .A(n40), .ZN(n38) );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_3 ( clk, clear_acc, 
        data_out_x, data_out, data_out_w, data_out_b, wr_en_y, m_valid, 
        m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [4:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
         N39, N40, N41, N42, N43, N44, n1, n2, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n85, n102, n111, n112, n113, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n18), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n222), .CK(clk), .Q(n22) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n223), .CK(clk), .Q(n23) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n224), .CK(clk), .Q(n24) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n225), .CK(clk), .Q(n25) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n226), .CK(clk), .Q(n26) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n227), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n228), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n229), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n230), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n231), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n232), .CK(clk), .Q(n34) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n233), .CK(clk), .Q(n35) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n234), .CK(clk), .Q(n36) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n235), .CK(clk), .Q(n37) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n236), .CK(clk), .Q(n38) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n237), .CK(clk), .Q(n40) );
  DFF_X1 \f_reg[0]  ( .D(n102), .CK(clk), .Q(f[0]), .QN(n210) );
  DFF_X1 \f_reg[1]  ( .D(n85), .CK(clk), .Q(f[1]), .QN(n211) );
  DFF_X1 \f_reg[2]  ( .D(n83), .CK(clk), .Q(f[2]), .QN(n212) );
  DFF_X1 \f_reg[3]  ( .D(n82), .CK(clk), .Q(f[3]), .QN(n213) );
  DFF_X1 \f_reg[7]  ( .D(n78), .CK(clk), .Q(f[7]), .QN(n214) );
  DFF_X1 \f_reg[8]  ( .D(n77), .CK(clk), .Q(f[8]), .QN(n215) );
  DFF_X1 \f_reg[9]  ( .D(n76), .CK(clk), .Q(f[9]), .QN(n216) );
  DFF_X1 \f_reg[10]  ( .D(n75), .CK(clk), .Q(n50), .QN(n217) );
  DFF_X1 \f_reg[11]  ( .D(n74), .CK(clk), .Q(n48), .QN(n218) );
  DFF_X1 \f_reg[12]  ( .D(n1), .CK(clk), .Q(n47), .QN(n219) );
  DFF_X1 \f_reg[13]  ( .D(n73), .CK(clk), .Q(n45), .QN(n220) );
  DFF_X1 \f_reg[14]  ( .D(n4), .CK(clk), .Q(n44), .QN(n221) );
  DFF_X1 \f_reg[15]  ( .D(n2), .CK(clk), .Q(f[15]), .QN(n70) );
  DFF_X1 \data_out_reg[15]  ( .D(n112), .CK(clk), .Q(data_out[15]), .QN(n193)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n113), .CK(clk), .Q(data_out[14]), .QN(n192)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n164), .CK(clk), .Q(data_out[13]), .QN(n191)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n165), .CK(clk), .Q(data_out[12]), .QN(n190)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n166), .CK(clk), .Q(data_out[11]), .QN(n189)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n167), .CK(clk), .Q(data_out[10]), .QN(n188)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n168), .CK(clk), .Q(data_out[9]), .QN(n187) );
  DFF_X1 \data_out_reg[8]  ( .D(n169), .CK(clk), .Q(data_out[8]), .QN(n186) );
  DFF_X1 \data_out_reg[7]  ( .D(n170), .CK(clk), .Q(data_out[7]), .QN(n185) );
  DFF_X1 \data_out_reg[6]  ( .D(n171), .CK(clk), .Q(data_out[6]), .QN(n184) );
  DFF_X1 \data_out_reg[5]  ( .D(n172), .CK(clk), .Q(data_out[5]), .QN(n183) );
  DFF_X1 \data_out_reg[4]  ( .D(n173), .CK(clk), .Q(data_out[4]), .QN(n182) );
  DFF_X1 \data_out_reg[3]  ( .D(n174), .CK(clk), .Q(data_out[3]), .QN(n181) );
  DFF_X1 \data_out_reg[2]  ( .D(n175), .CK(clk), .Q(data_out[2]), .QN(n180) );
  DFF_X1 \data_out_reg[1]  ( .D(n176), .CK(clk), .Q(data_out[1]), .QN(n179) );
  DFF_X1 \data_out_reg[0]  ( .D(n177), .CK(clk), .Q(data_out[0]), .QN(n178) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_3_DW_mult_tc_1 mult_2021 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_3_DW01_add_2 add_2022 ( .A({n200, 
        n199, n198, n197, n196, n195, n209, n208, n207, n206, n205, n204, n203, 
        n202, n201, n194}), .B({f[15], n44, n45, n47, n48, n50, f[9:0]}), .CI(
        1'b0), .SUM(adder) );
  DFF_X1 \f_reg[4]  ( .D(n81), .CK(clk), .Q(f[4]), .QN(n63) );
  DFF_X1 \f_reg[5]  ( .D(n80), .CK(clk), .Q(f[5]), .QN(n64) );
  DFF_X1 \f_reg[6]  ( .D(n79), .CK(clk), .Q(f[6]), .QN(n65) );
  DFF_X2 delay_reg ( .D(n111), .CK(clk), .Q(n5), .QN(n238) );
  MUX2_X1 U3 ( .A(N39), .B(n27), .S(n5), .Z(n195) );
  MUX2_X2 U4 ( .A(n29), .B(N37), .S(n238), .Z(n208) );
  AND2_X1 U5 ( .A1(n43), .A2(n19), .ZN(n16) );
  MUX2_X2 U6 ( .A(n32), .B(N36), .S(n238), .Z(n207) );
  MUX2_X2 U8 ( .A(N43), .B(n23), .S(n5), .Z(n199) );
  NAND3_X1 U9 ( .A1(n8), .A2(n7), .A3(n9), .ZN(n1) );
  MUX2_X1 U10 ( .A(n28), .B(N38), .S(n238), .Z(n209) );
  MUX2_X2 U11 ( .A(n25), .B(N41), .S(n238), .Z(n197) );
  MUX2_X2 U12 ( .A(n24), .B(N42), .S(n238), .Z(n198) );
  NAND3_X1 U13 ( .A1(n11), .A2(n10), .A3(n12), .ZN(n2) );
  NAND3_X1 U14 ( .A1(n14), .A2(n13), .A3(n15), .ZN(n4) );
  CLKBUF_X1 U15 ( .A(N43), .Z(n6) );
  NAND2_X1 U16 ( .A1(data_out_b[12]), .A2(n18), .ZN(n7) );
  NAND2_X1 U17 ( .A1(adder[12]), .A2(n16), .ZN(n8) );
  NAND2_X1 U18 ( .A1(n61), .A2(n47), .ZN(n9) );
  NAND2_X1 U19 ( .A1(data_out_b[15]), .A2(n18), .ZN(n10) );
  NAND2_X1 U20 ( .A1(adder[15]), .A2(n16), .ZN(n11) );
  NAND2_X1 U21 ( .A1(n61), .A2(f[15]), .ZN(n12) );
  NAND2_X1 U22 ( .A1(data_out_b[14]), .A2(n18), .ZN(n13) );
  NAND2_X1 U23 ( .A1(adder[14]), .A2(n16), .ZN(n14) );
  NAND2_X1 U24 ( .A1(n61), .A2(n44), .ZN(n15) );
  INV_X1 U25 ( .A(n19), .ZN(n18) );
  NAND2_X1 U26 ( .A1(n111), .A2(n17), .ZN(n240) );
  INV_X1 U27 ( .A(n43), .ZN(n61) );
  INV_X1 U28 ( .A(clear_acc), .ZN(n19) );
  OAI22_X1 U29 ( .A1(n181), .A2(n240), .B1(n213), .B2(n239), .ZN(n174) );
  OAI22_X1 U30 ( .A1(n182), .A2(n240), .B1(n63), .B2(n239), .ZN(n173) );
  OAI22_X1 U31 ( .A1(n183), .A2(n240), .B1(n64), .B2(n239), .ZN(n172) );
  OAI22_X1 U32 ( .A1(n184), .A2(n240), .B1(n65), .B2(n239), .ZN(n171) );
  OAI22_X1 U33 ( .A1(n185), .A2(n240), .B1(n214), .B2(n239), .ZN(n170) );
  OAI22_X1 U34 ( .A1(n186), .A2(n240), .B1(n215), .B2(n239), .ZN(n169) );
  OAI22_X1 U35 ( .A1(n187), .A2(n240), .B1(n216), .B2(n239), .ZN(n168) );
  MUX2_X1 U36 ( .A(n36), .B(N32), .S(n238), .Z(n203) );
  INV_X1 U37 ( .A(n21), .ZN(n39) );
  INV_X1 U38 ( .A(wr_en_y), .ZN(n17) );
  INV_X1 U39 ( .A(m_ready), .ZN(n20) );
  NAND2_X1 U40 ( .A1(m_valid), .A2(n20), .ZN(n41) );
  OAI21_X1 U41 ( .B1(sel[4]), .B2(n72), .A(n41), .ZN(n111) );
  NAND2_X1 U42 ( .A1(clear_acc_delay), .A2(n238), .ZN(n21) );
  MUX2_X1 U43 ( .A(n22), .B(N44), .S(n39), .Z(n222) );
  MUX2_X1 U44 ( .A(n22), .B(N44), .S(n238), .Z(n200) );
  MUX2_X1 U45 ( .A(n23), .B(n6), .S(n39), .Z(n223) );
  MUX2_X1 U46 ( .A(n24), .B(N42), .S(n39), .Z(n224) );
  MUX2_X1 U47 ( .A(n25), .B(N41), .S(n39), .Z(n225) );
  MUX2_X1 U48 ( .A(n26), .B(N40), .S(n39), .Z(n226) );
  MUX2_X1 U49 ( .A(n26), .B(N40), .S(n238), .Z(n196) );
  MUX2_X1 U50 ( .A(n27), .B(N39), .S(n39), .Z(n227) );
  MUX2_X1 U51 ( .A(n28), .B(N38), .S(n39), .Z(n228) );
  MUX2_X1 U52 ( .A(n29), .B(N37), .S(n39), .Z(n229) );
  MUX2_X1 U53 ( .A(n32), .B(N36), .S(n39), .Z(n230) );
  MUX2_X1 U54 ( .A(n33), .B(N35), .S(n39), .Z(n231) );
  MUX2_X1 U55 ( .A(n33), .B(N35), .S(n238), .Z(n206) );
  MUX2_X1 U56 ( .A(n34), .B(N34), .S(n39), .Z(n232) );
  MUX2_X1 U57 ( .A(n34), .B(N34), .S(n238), .Z(n205) );
  MUX2_X1 U58 ( .A(n35), .B(N33), .S(n39), .Z(n233) );
  MUX2_X1 U59 ( .A(n35), .B(N33), .S(n238), .Z(n204) );
  MUX2_X1 U60 ( .A(n36), .B(N32), .S(n39), .Z(n234) );
  MUX2_X1 U61 ( .A(n37), .B(N31), .S(n39), .Z(n235) );
  MUX2_X1 U62 ( .A(n37), .B(N31), .S(n238), .Z(n202) );
  MUX2_X1 U63 ( .A(n38), .B(N30), .S(n39), .Z(n236) );
  MUX2_X1 U64 ( .A(n38), .B(N30), .S(n238), .Z(n201) );
  MUX2_X1 U65 ( .A(n40), .B(N29), .S(n39), .Z(n237) );
  MUX2_X1 U66 ( .A(n40), .B(N29), .S(n238), .Z(n194) );
  INV_X1 U67 ( .A(n41), .ZN(n42) );
  OAI21_X1 U68 ( .B1(n42), .B2(n5), .A(n19), .ZN(n43) );
  AOI222_X1 U69 ( .A1(data_out_b[13]), .A2(n18), .B1(adder[13]), .B2(n16), 
        .C1(n61), .C2(n45), .ZN(n46) );
  INV_X1 U70 ( .A(n46), .ZN(n73) );
  AOI222_X1 U71 ( .A1(data_out_b[11]), .A2(n18), .B1(adder[11]), .B2(n16), 
        .C1(n61), .C2(n48), .ZN(n49) );
  INV_X1 U72 ( .A(n49), .ZN(n74) );
  AOI222_X1 U73 ( .A1(data_out_b[10]), .A2(n18), .B1(adder[10]), .B2(n16), 
        .C1(n61), .C2(n50), .ZN(n51) );
  INV_X1 U74 ( .A(n51), .ZN(n75) );
  AOI222_X1 U75 ( .A1(data_out_b[8]), .A2(n18), .B1(adder[8]), .B2(n16), .C1(
        n61), .C2(f[8]), .ZN(n52) );
  INV_X1 U76 ( .A(n52), .ZN(n77) );
  AOI222_X1 U77 ( .A1(data_out_b[7]), .A2(n18), .B1(adder[7]), .B2(n16), .C1(
        n61), .C2(f[7]), .ZN(n53) );
  INV_X1 U78 ( .A(n53), .ZN(n78) );
  AOI222_X1 U79 ( .A1(data_out_b[6]), .A2(n18), .B1(adder[6]), .B2(n16), .C1(
        n61), .C2(f[6]), .ZN(n54) );
  INV_X1 U80 ( .A(n54), .ZN(n79) );
  AOI222_X1 U81 ( .A1(data_out_b[5]), .A2(n18), .B1(adder[5]), .B2(n16), .C1(
        n61), .C2(f[5]), .ZN(n55) );
  INV_X1 U82 ( .A(n55), .ZN(n80) );
  AOI222_X1 U83 ( .A1(data_out_b[4]), .A2(n18), .B1(adder[4]), .B2(n16), .C1(
        n61), .C2(f[4]), .ZN(n56) );
  INV_X1 U84 ( .A(n56), .ZN(n81) );
  AOI222_X1 U85 ( .A1(data_out_b[3]), .A2(n18), .B1(adder[3]), .B2(n16), .C1(
        n61), .C2(f[3]), .ZN(n57) );
  INV_X1 U86 ( .A(n57), .ZN(n82) );
  AOI222_X1 U87 ( .A1(data_out_b[2]), .A2(n18), .B1(adder[2]), .B2(n16), .C1(
        n61), .C2(f[2]), .ZN(n58) );
  INV_X1 U88 ( .A(n58), .ZN(n83) );
  AOI222_X1 U89 ( .A1(data_out_b[1]), .A2(n18), .B1(adder[1]), .B2(n16), .C1(
        n61), .C2(f[1]), .ZN(n59) );
  INV_X1 U90 ( .A(n59), .ZN(n85) );
  AOI222_X1 U91 ( .A1(data_out_b[0]), .A2(n18), .B1(adder[0]), .B2(n16), .C1(
        n61), .C2(f[0]), .ZN(n60) );
  INV_X1 U92 ( .A(n60), .ZN(n102) );
  AOI222_X1 U93 ( .A1(data_out_b[9]), .A2(n18), .B1(adder[9]), .B2(n16), .C1(
        n61), .C2(f[9]), .ZN(n62) );
  INV_X1 U94 ( .A(n62), .ZN(n76) );
  NOR4_X1 U95 ( .A1(n48), .A2(n47), .A3(n45), .A4(n44), .ZN(n69) );
  NOR4_X1 U96 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n50), .ZN(n68) );
  NAND4_X1 U97 ( .A1(n65), .A2(n64), .A3(n63), .A4(n213), .ZN(n66) );
  NOR4_X1 U98 ( .A1(n66), .A2(f[0]), .A3(f[1]), .A4(f[2]), .ZN(n67) );
  NAND3_X1 U99 ( .A1(n69), .A2(n68), .A3(n67), .ZN(n71) );
  NAND3_X1 U100 ( .A1(wr_en_y), .A2(n71), .A3(n70), .ZN(n239) );
  OAI22_X1 U101 ( .A1(n178), .A2(n240), .B1(n210), .B2(n239), .ZN(n177) );
  OAI22_X1 U102 ( .A1(n179), .A2(n240), .B1(n211), .B2(n239), .ZN(n176) );
  OAI22_X1 U103 ( .A1(n180), .A2(n240), .B1(n212), .B2(n239), .ZN(n175) );
  OAI22_X1 U104 ( .A1(n188), .A2(n240), .B1(n217), .B2(n239), .ZN(n167) );
  OAI22_X1 U105 ( .A1(n189), .A2(n240), .B1(n218), .B2(n239), .ZN(n166) );
  OAI22_X1 U106 ( .A1(n190), .A2(n240), .B1(n219), .B2(n239), .ZN(n165) );
  OAI22_X1 U107 ( .A1(n191), .A2(n240), .B1(n220), .B2(n239), .ZN(n164) );
  OAI22_X1 U108 ( .A1(n192), .A2(n240), .B1(n221), .B2(n239), .ZN(n113) );
  OAI22_X1 U109 ( .A1(n193), .A2(n240), .B1(n70), .B2(n239), .ZN(n112) );
  AND4_X1 U110 ( .A1(sel[3]), .A2(sel[2]), .A3(sel[1]), .A4(sel[0]), .ZN(n72)
         );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_2_DW_mult_tc_1 ( a, b, 
        product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n9, n12, n13, n16, n18, n19, n21, n23, n25, n27, n29, n31,
         n32, n34, n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n50,
         n53, n54, n55, n56, n57, n58, n59, n62, n63, n64, n65, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n93, n95, n96, n97, n98, n99, n101,
         n103, n104, n105, n106, n107, n111, n112, n113, n114, n115, n117,
         n119, n120, n122, n125, n135, n139, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n247, n249, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n418, n419,
         n420, n421, n422, n423, n424, n426, n427, n429, n433, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U148 ( .A(n265), .B(n144), .Z(n145) );
  XOR2_X1 U150 ( .A(n271), .B(n146), .Z(n147) );
  XOR2_X1 U152 ( .A(n301), .B(n148), .Z(n149) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U162 ( .A(n170), .B(n172), .CI(n179), .CO(n165), .S(n166) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n263), .CI(n291), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n317), .B(n252), .CO(n173), .S(n174) );
  FA_X1 U167 ( .A(n180), .B(n187), .CI(n178), .CO(n175), .S(n176) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U169 ( .A(n193), .B(n282), .CI(n191), .CO(n179), .S(n180) );
  FA_X1 U170 ( .A(n268), .B(n292), .CI(n274), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U172 ( .A(n197), .B(n190), .CI(n188), .CO(n185), .S(n186) );
  FA_X1 U173 ( .A(n199), .B(n201), .CI(n192), .CO(n187), .S(n188) );
  FA_X1 U174 ( .A(n275), .B(n293), .CI(n194), .CO(n189), .S(n190) );
  FA_X1 U175 ( .A(n283), .B(n253), .CI(n305), .CO(n191), .S(n192) );
  HA_X1 U176 ( .A(n319), .B(n269), .CO(n193), .S(n194) );
  FA_X1 U177 ( .A(n205), .B(n200), .CI(n198), .CO(n195), .S(n196) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U179 ( .A(n284), .B(n294), .CI(n276), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n320), .B(n270), .CI(n306), .CO(n201), .S(n202) );
  FA_X1 U181 ( .A(n208), .B(n213), .CI(n206), .CO(n203), .S(n204) );
  FA_X1 U182 ( .A(n215), .B(n307), .CI(n210), .CO(n205), .S(n206) );
  FA_X1 U183 ( .A(n295), .B(n285), .CI(n254), .CO(n207), .S(n208) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U185 ( .A(n216), .B(n219), .CI(n214), .CO(n211), .S(n212) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n322), .B(n278), .CI(n308), .CO(n215), .S(n216) );
  FA_X1 U188 ( .A(n225), .B(n222), .CI(n220), .CO(n217), .S(n218) );
  FA_X1 U189 ( .A(n309), .B(n255), .CI(n297), .CO(n219), .S(n220) );
  HA_X1 U190 ( .A(n287), .B(n323), .CO(n221), .S(n222) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  HA_X1 U194 ( .A(n311), .B(n325), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n326), .B(n300), .CI(n312), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  XNOR2_X1 U414 ( .A(n586), .B(a[6]), .ZN(n490) );
  CLKBUF_X1 U415 ( .A(n226), .Z(n491) );
  INV_X1 U416 ( .A(n1), .ZN(n492) );
  INV_X1 U417 ( .A(n490), .ZN(n21) );
  BUF_X1 U418 ( .A(n106), .Z(n497) );
  BUF_X1 U419 ( .A(n12), .Z(n539) );
  AND2_X1 U420 ( .A1(n578), .A2(n517), .ZN(n288) );
  INV_X1 U421 ( .A(n530), .ZN(n37) );
  OR2_X1 U422 ( .A1(n329), .A2(n258), .ZN(n493) );
  BUF_X1 U423 ( .A(n96), .Z(n542) );
  XOR2_X1 U424 ( .A(n594), .B(a[14]), .Z(n41) );
  INV_X1 U425 ( .A(n507), .ZN(n494) );
  XNOR2_X1 U426 ( .A(n590), .B(a[8]), .ZN(n429) );
  INV_X1 U427 ( .A(n561), .ZN(n495) );
  OR2_X1 U428 ( .A1(n218), .A2(n223), .ZN(n496) );
  INV_X1 U429 ( .A(n561), .ZN(n16) );
  AND2_X1 U430 ( .A1(n232), .A2(n233), .ZN(n498) );
  BUF_X1 U431 ( .A(n104), .Z(n511) );
  INV_X1 U432 ( .A(n552), .ZN(n499) );
  INV_X1 U433 ( .A(n552), .ZN(n27) );
  CLKBUF_X1 U434 ( .A(n508), .Z(n500) );
  XNOR2_X1 U435 ( .A(n554), .B(n501), .ZN(product[9]) );
  AND2_X1 U436 ( .A1(n515), .A2(n90), .ZN(n501) );
  BUF_X1 U437 ( .A(n88), .Z(n502) );
  CLKBUF_X1 U438 ( .A(n83), .Z(n503) );
  CLKBUF_X1 U439 ( .A(n186), .Z(n504) );
  XNOR2_X1 U440 ( .A(n505), .B(n226), .ZN(n224) );
  XNOR2_X1 U441 ( .A(n229), .B(n298), .ZN(n505) );
  OR2_X1 U442 ( .A1(n504), .A2(n195), .ZN(n506) );
  INV_X1 U443 ( .A(n590), .ZN(n507) );
  BUF_X1 U444 ( .A(n12), .Z(n508) );
  BUF_X1 U445 ( .A(n12), .Z(n540) );
  OR2_X1 U446 ( .A1(n196), .A2(n203), .ZN(n509) );
  XNOR2_X1 U447 ( .A(n45), .B(n510), .ZN(product[12]) );
  AND2_X1 U448 ( .A1(n523), .A2(n79), .ZN(n510) );
  AOI21_X1 U449 ( .B1(n570), .B2(n112), .A(n498), .ZN(n512) );
  AOI21_X1 U450 ( .B1(n96), .B2(n567), .A(n93), .ZN(n513) );
  AOI21_X1 U451 ( .B1(n96), .B2(n567), .A(n93), .ZN(n91) );
  INV_X1 U452 ( .A(n7), .ZN(n584) );
  INV_X2 U453 ( .A(n594), .ZN(n593) );
  AOI21_X1 U454 ( .B1(n571), .B2(n511), .A(n101), .ZN(n514) );
  OR2_X1 U455 ( .A1(n204), .A2(n211), .ZN(n515) );
  OR2_X1 U456 ( .A1(n228), .A2(n231), .ZN(n516) );
  INV_X1 U457 ( .A(n21), .ZN(n517) );
  CLKBUF_X1 U458 ( .A(n86), .Z(n518) );
  INV_X1 U459 ( .A(n584), .ZN(n519) );
  INV_X1 U460 ( .A(n584), .ZN(n520) );
  INV_X1 U461 ( .A(n584), .ZN(n583) );
  BUF_X2 U462 ( .A(n526), .Z(n521) );
  BUF_X1 U463 ( .A(n324), .Z(n522) );
  XNOR2_X1 U464 ( .A(n584), .B(a[2]), .ZN(n565) );
  OR2_X1 U465 ( .A1(n176), .A2(n185), .ZN(n523) );
  NOR2_X1 U466 ( .A1(n186), .A2(n195), .ZN(n524) );
  NOR2_X1 U467 ( .A1(n186), .A2(n195), .ZN(n82) );
  INV_X1 U468 ( .A(n587), .ZN(n525) );
  XOR2_X1 U469 ( .A(n492), .B(a[2]), .Z(n526) );
  CLKBUF_X1 U470 ( .A(n521), .Z(n527) );
  INV_X1 U471 ( .A(n520), .ZN(n528) );
  OAI21_X1 U472 ( .B1(n513), .B2(n89), .A(n90), .ZN(n529) );
  XNOR2_X1 U473 ( .A(n592), .B(a[12]), .ZN(n530) );
  INV_X1 U474 ( .A(n592), .ZN(n591) );
  CLKBUF_X1 U475 ( .A(n553), .Z(n538) );
  INV_X1 U476 ( .A(n586), .ZN(n531) );
  OAI21_X1 U477 ( .B1(n524), .B2(n86), .A(n83), .ZN(n532) );
  INV_X1 U478 ( .A(n590), .ZN(n589) );
  INV_X1 U479 ( .A(n580), .ZN(n533) );
  INV_X2 U480 ( .A(n492), .ZN(n581) );
  CLKBUF_X1 U481 ( .A(n85), .Z(n534) );
  XNOR2_X1 U482 ( .A(n166), .B(n535), .ZN(n164) );
  XNOR2_X1 U483 ( .A(n168), .B(n177), .ZN(n535) );
  INV_X1 U484 ( .A(n247), .ZN(n536) );
  INV_X1 U485 ( .A(n582), .ZN(n580) );
  NAND2_X2 U486 ( .A1(n429), .A2(n27), .ZN(n29) );
  OR2_X2 U487 ( .A1(n537), .A2(n564), .ZN(n23) );
  XOR2_X1 U488 ( .A(n588), .B(a[6]), .Z(n537) );
  BUF_X2 U489 ( .A(n526), .Z(n575) );
  XOR2_X1 U490 ( .A(n592), .B(a[10]), .Z(n546) );
  NAND2_X1 U491 ( .A1(n9), .A2(n565), .ZN(n12) );
  XNOR2_X1 U492 ( .A(n529), .B(n541), .ZN(product[10]) );
  NAND2_X1 U493 ( .A1(n86), .A2(n509), .ZN(n541) );
  NAND2_X1 U494 ( .A1(n166), .A2(n168), .ZN(n543) );
  NAND2_X1 U495 ( .A1(n166), .A2(n177), .ZN(n544) );
  NAND2_X1 U496 ( .A1(n168), .A2(n177), .ZN(n545) );
  NAND3_X1 U497 ( .A1(n543), .A2(n544), .A3(n545), .ZN(n163) );
  OR2_X2 U498 ( .A1(n546), .A2(n551), .ZN(n34) );
  NOR2_X2 U499 ( .A1(n164), .A2(n175), .ZN(n75) );
  INV_X1 U500 ( .A(n551), .ZN(n32) );
  OR2_X1 U501 ( .A1(n547), .A2(n561), .ZN(n18) );
  XNOR2_X1 U502 ( .A(n13), .B(a[4]), .ZN(n547) );
  OR2_X1 U503 ( .A1(n547), .A2(n561), .ZN(n548) );
  OR2_X1 U504 ( .A1(n547), .A2(n561), .ZN(n549) );
  XNOR2_X1 U505 ( .A(n550), .B(n310), .ZN(n226) );
  XNOR2_X1 U506 ( .A(n324), .B(n288), .ZN(n550) );
  INV_X1 U507 ( .A(n19), .ZN(n588) );
  XNOR2_X1 U508 ( .A(n590), .B(a[10]), .ZN(n551) );
  XNOR2_X1 U509 ( .A(n588), .B(a[8]), .ZN(n552) );
  XOR2_X1 U510 ( .A(n582), .B(a[2]), .Z(n9) );
  AOI21_X1 U511 ( .B1(n529), .B2(n80), .A(n81), .ZN(n553) );
  AOI21_X1 U512 ( .B1(n502), .B2(n80), .A(n532), .ZN(n45) );
  CLKBUF_X1 U513 ( .A(n513), .Z(n554) );
  NAND2_X1 U514 ( .A1(n522), .A2(n288), .ZN(n555) );
  NAND2_X1 U515 ( .A1(n522), .A2(n310), .ZN(n556) );
  NAND2_X1 U516 ( .A1(n288), .A2(n310), .ZN(n557) );
  NAND3_X1 U517 ( .A1(n555), .A2(n556), .A3(n557), .ZN(n225) );
  NAND2_X1 U518 ( .A1(n229), .A2(n298), .ZN(n558) );
  NAND2_X1 U519 ( .A1(n229), .A2(n491), .ZN(n559) );
  NAND2_X1 U520 ( .A1(n298), .A2(n491), .ZN(n560) );
  NAND3_X1 U521 ( .A1(n558), .A2(n559), .A3(n560), .ZN(n223) );
  XNOR2_X1 U522 ( .A(n582), .B(n249), .ZN(n433) );
  INV_X2 U523 ( .A(n249), .ZN(n579) );
  XNOR2_X1 U524 ( .A(n584), .B(a[4]), .ZN(n561) );
  INV_X2 U525 ( .A(n588), .ZN(n587) );
  NAND2_X1 U526 ( .A1(n433), .A2(n579), .ZN(n562) );
  NAND2_X1 U527 ( .A1(n433), .A2(n579), .ZN(n563) );
  XNOR2_X1 U528 ( .A(n586), .B(a[6]), .ZN(n564) );
  BUF_X1 U529 ( .A(n43), .Z(n577) );
  AOI21_X1 U530 ( .B1(n566), .B2(n74), .A(n67), .ZN(n65) );
  INV_X1 U531 ( .A(n69), .ZN(n67) );
  NAND2_X1 U532 ( .A1(n566), .A2(n69), .ZN(n47) );
  INV_X1 U533 ( .A(n73), .ZN(n71) );
  NAND2_X1 U534 ( .A1(n73), .A2(n566), .ZN(n64) );
  INV_X1 U535 ( .A(n74), .ZN(n72) );
  INV_X1 U536 ( .A(n95), .ZN(n93) );
  NOR2_X1 U537 ( .A1(n524), .A2(n85), .ZN(n80) );
  OAI21_X1 U538 ( .B1(n82), .B2(n86), .A(n83), .ZN(n81) );
  NAND2_X1 U539 ( .A1(n506), .A2(n503), .ZN(n50) );
  OR2_X1 U540 ( .A1(n152), .A2(n163), .ZN(n566) );
  OAI21_X1 U541 ( .B1(n75), .B2(n79), .A(n76), .ZN(n74) );
  NAND2_X1 U542 ( .A1(n125), .A2(n76), .ZN(n48) );
  INV_X1 U543 ( .A(n75), .ZN(n125) );
  NOR2_X1 U544 ( .A1(n75), .A2(n78), .ZN(n73) );
  NAND2_X1 U545 ( .A1(n152), .A2(n163), .ZN(n69) );
  NAND2_X1 U546 ( .A1(n567), .A2(n95), .ZN(n53) );
  NAND2_X1 U547 ( .A1(n516), .A2(n497), .ZN(n56) );
  NAND2_X1 U548 ( .A1(n496), .A2(n98), .ZN(n54) );
  AOI21_X1 U549 ( .B1(n568), .B2(n120), .A(n117), .ZN(n115) );
  INV_X1 U550 ( .A(n119), .ZN(n117) );
  NOR2_X1 U551 ( .A1(n196), .A2(n203), .ZN(n85) );
  NOR2_X1 U552 ( .A1(n176), .A2(n185), .ZN(n78) );
  NAND2_X1 U553 ( .A1(n570), .A2(n111), .ZN(n57) );
  XOR2_X1 U554 ( .A(n58), .B(n115), .Z(product[3]) );
  XNOR2_X1 U555 ( .A(n59), .B(n120), .ZN(product[2]) );
  NAND2_X1 U556 ( .A1(n568), .A2(n119), .ZN(n59) );
  NAND2_X1 U557 ( .A1(n176), .A2(n185), .ZN(n79) );
  NAND2_X1 U558 ( .A1(n196), .A2(n203), .ZN(n86) );
  NAND2_X1 U559 ( .A1(n164), .A2(n175), .ZN(n76) );
  NAND2_X1 U560 ( .A1(n186), .A2(n195), .ZN(n83) );
  NAND2_X1 U561 ( .A1(n212), .A2(n217), .ZN(n95) );
  OR2_X1 U562 ( .A1(n212), .A2(n217), .ZN(n567) );
  NAND2_X1 U563 ( .A1(n204), .A2(n211), .ZN(n90) );
  NAND2_X1 U564 ( .A1(n569), .A2(n62), .ZN(n46) );
  OR2_X1 U565 ( .A1(n328), .A2(n314), .ZN(n568) );
  OR2_X1 U566 ( .A1(n151), .A2(n139), .ZN(n569) );
  NAND2_X1 U567 ( .A1(n328), .A2(n314), .ZN(n119) );
  NOR2_X1 U568 ( .A1(n218), .A2(n223), .ZN(n97) );
  NAND2_X1 U569 ( .A1(n218), .A2(n223), .ZN(n98) );
  OR2_X1 U570 ( .A1(n232), .A2(n233), .ZN(n570) );
  INV_X1 U571 ( .A(n41), .ZN(n235) );
  OR2_X1 U572 ( .A1(n224), .A2(n227), .ZN(n571) );
  AND2_X1 U573 ( .A1(n493), .A2(n122), .ZN(product[1]) );
  OAI22_X1 U574 ( .A1(n563), .A2(n407), .B1(n406), .B2(n579), .ZN(n328) );
  OR2_X1 U575 ( .A1(n577), .A2(n528), .ZN(n392) );
  NAND2_X1 U576 ( .A1(n433), .A2(n579), .ZN(n6) );
  OAI22_X1 U577 ( .A1(n6), .A2(n400), .B1(n399), .B2(n579), .ZN(n321) );
  XNOR2_X1 U578 ( .A(n507), .B(n577), .ZN(n352) );
  OAI22_X1 U579 ( .A1(n563), .A2(n408), .B1(n407), .B2(n579), .ZN(n329) );
  XNOR2_X1 U580 ( .A(n155), .B(n573), .ZN(n139) );
  XNOR2_X1 U581 ( .A(n153), .B(n141), .ZN(n573) );
  XNOR2_X1 U582 ( .A(n157), .B(n574), .ZN(n141) );
  XNOR2_X1 U583 ( .A(n145), .B(n143), .ZN(n574) );
  OAI22_X1 U584 ( .A1(n562), .A2(n396), .B1(n395), .B2(n579), .ZN(n317) );
  OAI22_X1 U585 ( .A1(n39), .A2(n594), .B1(n337), .B2(n37), .ZN(n252) );
  OR2_X1 U586 ( .A1(n577), .A2(n594), .ZN(n337) );
  OAI22_X1 U587 ( .A1(n562), .A2(n398), .B1(n397), .B2(n579), .ZN(n319) );
  XNOR2_X1 U588 ( .A(n591), .B(n577), .ZN(n343) );
  OAI22_X1 U589 ( .A1(n563), .A2(n404), .B1(n403), .B2(n579), .ZN(n325) );
  OAI22_X1 U590 ( .A1(n42), .A2(n596), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U591 ( .A1(n577), .A2(n596), .ZN(n332) );
  AND2_X1 U592 ( .A1(n578), .A2(n561), .ZN(n300) );
  OAI22_X1 U593 ( .A1(n562), .A2(n405), .B1(n404), .B2(n579), .ZN(n326) );
  XOR2_X1 U594 ( .A(n315), .B(n261), .Z(n150) );
  OAI22_X1 U595 ( .A1(n6), .A2(n394), .B1(n393), .B2(n579), .ZN(n315) );
  OAI22_X1 U596 ( .A1(n6), .A2(n406), .B1(n405), .B2(n579), .ZN(n327) );
  XNOR2_X1 U597 ( .A(n520), .B(n577), .ZN(n391) );
  XNOR2_X1 U598 ( .A(n593), .B(n577), .ZN(n336) );
  AND2_X1 U599 ( .A1(n578), .A2(n247), .ZN(n314) );
  NAND2_X1 U600 ( .A1(n427), .A2(n37), .ZN(n39) );
  XOR2_X1 U601 ( .A(n593), .B(a[12]), .Z(n427) );
  AND2_X1 U602 ( .A1(n578), .A2(n552), .ZN(n278) );
  OAI22_X1 U603 ( .A1(n563), .A2(n401), .B1(n400), .B2(n579), .ZN(n322) );
  OAI22_X1 U604 ( .A1(n39), .A2(n336), .B1(n37), .B2(n335), .ZN(n263) );
  XNOR2_X1 U605 ( .A(n585), .B(n577), .ZN(n376) );
  OAI22_X1 U606 ( .A1(n6), .A2(n397), .B1(n396), .B2(n579), .ZN(n318) );
  AND2_X1 U607 ( .A1(n578), .A2(n530), .ZN(n264) );
  OAI22_X1 U608 ( .A1(n6), .A2(n403), .B1(n402), .B2(n579), .ZN(n324) );
  AND2_X1 U609 ( .A1(n578), .A2(n551), .ZN(n270) );
  OAI22_X1 U610 ( .A1(n562), .A2(n399), .B1(n398), .B2(n579), .ZN(n320) );
  AND2_X1 U611 ( .A1(n578), .A2(n235), .ZN(n260) );
  OAI22_X1 U612 ( .A1(n563), .A2(n395), .B1(n394), .B2(n579), .ZN(n316) );
  OAI22_X1 U613 ( .A1(n39), .A2(n335), .B1(n37), .B2(n334), .ZN(n262) );
  INV_X1 U614 ( .A(n25), .ZN(n590) );
  NAND2_X1 U615 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U616 ( .A(n595), .B(a[14]), .Z(n426) );
  INV_X1 U617 ( .A(n13), .ZN(n586) );
  OAI22_X1 U618 ( .A1(n6), .A2(n402), .B1(n401), .B2(n579), .ZN(n323) );
  XNOR2_X1 U619 ( .A(n587), .B(n577), .ZN(n363) );
  AND2_X1 U620 ( .A1(n578), .A2(n249), .ZN(product[0]) );
  OR2_X1 U621 ( .A1(n577), .A2(n525), .ZN(n364) );
  OR2_X1 U622 ( .A1(n577), .A2(n592), .ZN(n344) );
  OR2_X1 U623 ( .A1(n577), .A2(n494), .ZN(n353) );
  OR2_X1 U624 ( .A1(n577), .A2(n586), .ZN(n377) );
  XNOR2_X1 U625 ( .A(n587), .B(b[9]), .ZN(n354) );
  OAI22_X1 U626 ( .A1(n39), .A2(n334), .B1(n37), .B2(n333), .ZN(n261) );
  XNOR2_X1 U627 ( .A(n593), .B(n422), .ZN(n333) );
  XNOR2_X1 U628 ( .A(n585), .B(b[11]), .ZN(n365) );
  XNOR2_X1 U629 ( .A(n593), .B(n424), .ZN(n335) );
  XNOR2_X1 U630 ( .A(n593), .B(n423), .ZN(n334) );
  OAI22_X1 U631 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U632 ( .A(n595), .B(n424), .ZN(n330) );
  XNOR2_X1 U633 ( .A(n595), .B(n577), .ZN(n331) );
  XNOR2_X1 U634 ( .A(n581), .B(b[11]), .ZN(n397) );
  XNOR2_X1 U635 ( .A(n581), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U636 ( .A(n581), .B(b[13]), .ZN(n395) );
  XNOR2_X1 U637 ( .A(n581), .B(b[14]), .ZN(n394) );
  XNOR2_X1 U638 ( .A(n507), .B(n418), .ZN(n345) );
  XNOR2_X1 U639 ( .A(n591), .B(n420), .ZN(n338) );
  XNOR2_X1 U640 ( .A(n519), .B(b[13]), .ZN(n378) );
  XNOR2_X1 U641 ( .A(n591), .B(n424), .ZN(n342) );
  XNOR2_X1 U642 ( .A(n587), .B(n424), .ZN(n362) );
  XNOR2_X1 U643 ( .A(n589), .B(n424), .ZN(n351) );
  XNOR2_X1 U644 ( .A(n591), .B(n423), .ZN(n341) );
  XNOR2_X1 U645 ( .A(n591), .B(n422), .ZN(n340) );
  XNOR2_X1 U646 ( .A(n591), .B(n421), .ZN(n339) );
  XNOR2_X1 U647 ( .A(n520), .B(n418), .ZN(n384) );
  XNOR2_X1 U648 ( .A(n519), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U649 ( .A(n583), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U650 ( .A(n519), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U651 ( .A(n519), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U652 ( .A(n520), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U653 ( .A(n520), .B(n419), .ZN(n385) );
  XNOR2_X1 U654 ( .A(n587), .B(n423), .ZN(n361) );
  XNOR2_X1 U655 ( .A(n507), .B(n423), .ZN(n350) );
  XNOR2_X1 U656 ( .A(n585), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U657 ( .A(n585), .B(n418), .ZN(n369) );
  XNOR2_X1 U658 ( .A(n585), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U659 ( .A(n585), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U660 ( .A(n587), .B(n422), .ZN(n360) );
  XNOR2_X1 U661 ( .A(n589), .B(n422), .ZN(n349) );
  XNOR2_X1 U662 ( .A(n587), .B(n421), .ZN(n359) );
  XNOR2_X1 U663 ( .A(n519), .B(n421), .ZN(n387) );
  XNOR2_X1 U664 ( .A(n589), .B(n421), .ZN(n348) );
  XNOR2_X1 U665 ( .A(n587), .B(n420), .ZN(n358) );
  XNOR2_X1 U666 ( .A(n507), .B(n420), .ZN(n347) );
  XNOR2_X1 U667 ( .A(n587), .B(n418), .ZN(n356) );
  XNOR2_X1 U668 ( .A(n587), .B(n419), .ZN(n357) );
  XNOR2_X1 U669 ( .A(n589), .B(n419), .ZN(n346) );
  XNOR2_X1 U670 ( .A(n587), .B(b[8]), .ZN(n355) );
  XNOR2_X1 U671 ( .A(n581), .B(b[15]), .ZN(n393) );
  BUF_X1 U672 ( .A(n43), .Z(n578) );
  OAI22_X1 U673 ( .A1(n34), .A2(n339), .B1(n338), .B2(n32), .ZN(n265) );
  OAI22_X1 U674 ( .A1(n34), .A2(n341), .B1(n340), .B2(n32), .ZN(n267) );
  OAI22_X1 U675 ( .A1(n34), .A2(n340), .B1(n339), .B2(n32), .ZN(n266) );
  OAI22_X1 U676 ( .A1(n34), .A2(n342), .B1(n341), .B2(n32), .ZN(n268) );
  OAI22_X1 U677 ( .A1(n34), .A2(n343), .B1(n342), .B2(n32), .ZN(n269) );
  OAI22_X1 U678 ( .A1(n34), .A2(n592), .B1(n344), .B2(n32), .ZN(n253) );
  NAND2_X1 U679 ( .A1(n228), .A2(n231), .ZN(n106) );
  NOR2_X1 U680 ( .A1(n228), .A2(n231), .ZN(n105) );
  XNOR2_X1 U681 ( .A(n583), .B(n423), .ZN(n389) );
  XNOR2_X1 U682 ( .A(n583), .B(n422), .ZN(n388) );
  XNOR2_X1 U683 ( .A(n519), .B(n424), .ZN(n390) );
  XNOR2_X1 U684 ( .A(n520), .B(n420), .ZN(n386) );
  XNOR2_X1 U685 ( .A(n77), .B(n48), .ZN(product[13]) );
  OAI21_X1 U686 ( .B1(n113), .B2(n115), .A(n114), .ZN(n576) );
  OAI21_X1 U687 ( .B1(n113), .B2(n115), .A(n114), .ZN(n112) );
  NOR2_X1 U688 ( .A1(n234), .A2(n257), .ZN(n113) );
  NAND2_X1 U689 ( .A1(n224), .A2(n227), .ZN(n103) );
  NOR2_X1 U690 ( .A1(n204), .A2(n211), .ZN(n89) );
  OAI22_X1 U691 ( .A1(n29), .A2(n350), .B1(n349), .B2(n499), .ZN(n275) );
  OAI22_X1 U692 ( .A1(n29), .A2(n346), .B1(n345), .B2(n499), .ZN(n271) );
  OAI22_X1 U693 ( .A1(n29), .A2(n347), .B1(n346), .B2(n499), .ZN(n272) );
  OAI22_X1 U694 ( .A1(n29), .A2(n348), .B1(n347), .B2(n499), .ZN(n273) );
  OAI22_X1 U695 ( .A1(n29), .A2(n349), .B1(n348), .B2(n499), .ZN(n274) );
  OAI22_X1 U696 ( .A1(n29), .A2(n351), .B1(n350), .B2(n499), .ZN(n276) );
  OAI22_X1 U697 ( .A1(n29), .A2(n494), .B1(n353), .B2(n499), .ZN(n254) );
  OAI22_X1 U698 ( .A1(n29), .A2(n352), .B1(n351), .B2(n499), .ZN(n277) );
  XNOR2_X1 U699 ( .A(n63), .B(n46), .ZN(product[15]) );
  NAND2_X1 U700 ( .A1(n571), .A2(n103), .ZN(n55) );
  INV_X1 U701 ( .A(n103), .ZN(n101) );
  XNOR2_X1 U702 ( .A(n84), .B(n50), .ZN(product[11]) );
  NAND2_X1 U703 ( .A1(n232), .A2(n233), .ZN(n111) );
  XNOR2_X1 U704 ( .A(n55), .B(n511), .ZN(product[6]) );
  INV_X1 U705 ( .A(n113), .ZN(n135) );
  OR2_X1 U706 ( .A1(n577), .A2(n533), .ZN(n409) );
  INV_X1 U707 ( .A(n1), .ZN(n582) );
  OAI21_X1 U708 ( .B1(n64), .B2(n538), .A(n65), .ZN(n63) );
  OAI21_X1 U709 ( .B1(n105), .B2(n107), .A(n106), .ZN(n104) );
  OAI22_X1 U710 ( .A1(n23), .A2(n358), .B1(n21), .B2(n357), .ZN(n282) );
  OAI22_X1 U711 ( .A1(n23), .A2(n356), .B1(n355), .B2(n21), .ZN(n280) );
  OAI22_X1 U712 ( .A1(n23), .A2(n360), .B1(n21), .B2(n359), .ZN(n284) );
  OAI22_X1 U713 ( .A1(n23), .A2(n357), .B1(n356), .B2(n21), .ZN(n281) );
  OAI22_X1 U714 ( .A1(n23), .A2(n362), .B1(n21), .B2(n361), .ZN(n286) );
  OAI22_X1 U715 ( .A1(n23), .A2(n355), .B1(n21), .B2(n354), .ZN(n279) );
  OAI22_X1 U716 ( .A1(n23), .A2(n361), .B1(n21), .B2(n360), .ZN(n285) );
  OAI22_X1 U717 ( .A1(n23), .A2(n525), .B1(n364), .B2(n21), .ZN(n255) );
  OAI22_X1 U718 ( .A1(n23), .A2(n359), .B1(n21), .B2(n358), .ZN(n283) );
  XNOR2_X1 U719 ( .A(n531), .B(n424), .ZN(n375) );
  OAI22_X1 U720 ( .A1(n23), .A2(n363), .B1(n362), .B2(n21), .ZN(n287) );
  XNOR2_X1 U721 ( .A(n531), .B(n419), .ZN(n370) );
  XNOR2_X1 U722 ( .A(n531), .B(n420), .ZN(n371) );
  XNOR2_X1 U723 ( .A(n531), .B(n421), .ZN(n372) );
  XNOR2_X1 U724 ( .A(n531), .B(n423), .ZN(n374) );
  XNOR2_X1 U725 ( .A(n531), .B(n422), .ZN(n373) );
  XNOR2_X1 U726 ( .A(n542), .B(n53), .ZN(product[8]) );
  AOI21_X1 U727 ( .B1(n104), .B2(n571), .A(n101), .ZN(n99) );
  OAI21_X1 U728 ( .B1(n99), .B2(n97), .A(n98), .ZN(n96) );
  NAND2_X1 U729 ( .A1(n151), .A2(n139), .ZN(n62) );
  OAI22_X1 U730 ( .A1(n549), .A2(n370), .B1(n369), .B2(n495), .ZN(n293) );
  OAI22_X1 U731 ( .A1(n548), .A2(n367), .B1(n366), .B2(n495), .ZN(n290) );
  OAI22_X1 U732 ( .A1(n548), .A2(n375), .B1(n374), .B2(n495), .ZN(n298) );
  OAI22_X1 U733 ( .A1(n549), .A2(n368), .B1(n367), .B2(n495), .ZN(n291) );
  OAI22_X1 U734 ( .A1(n548), .A2(n369), .B1(n368), .B2(n16), .ZN(n292) );
  OAI22_X1 U735 ( .A1(n549), .A2(n586), .B1(n377), .B2(n495), .ZN(n256) );
  OAI22_X1 U736 ( .A1(n548), .A2(n376), .B1(n375), .B2(n495), .ZN(n299) );
  OAI22_X1 U737 ( .A1(n549), .A2(n373), .B1(n372), .B2(n16), .ZN(n296) );
  OAI22_X1 U738 ( .A1(n18), .A2(n371), .B1(n370), .B2(n16), .ZN(n294) );
  OAI22_X1 U739 ( .A1(n549), .A2(n372), .B1(n371), .B2(n16), .ZN(n295) );
  OAI22_X1 U740 ( .A1(n18), .A2(n374), .B1(n373), .B2(n16), .ZN(n297) );
  OAI22_X1 U741 ( .A1(n548), .A2(n366), .B1(n365), .B2(n16), .ZN(n289) );
  OAI21_X1 U742 ( .B1(n87), .B2(n534), .A(n518), .ZN(n84) );
  XOR2_X1 U743 ( .A(n56), .B(n512), .Z(product[5]) );
  AOI21_X1 U744 ( .B1(n570), .B2(n112), .A(n498), .ZN(n107) );
  OAI21_X1 U745 ( .B1(n91), .B2(n89), .A(n90), .ZN(n88) );
  OAI21_X1 U746 ( .B1(n553), .B2(n78), .A(n79), .ZN(n77) );
  XNOR2_X1 U747 ( .A(n57), .B(n576), .ZN(product[4]) );
  INV_X1 U748 ( .A(n88), .ZN(n87) );
  NAND2_X1 U749 ( .A1(n135), .A2(n114), .ZN(n58) );
  XNOR2_X1 U750 ( .A(n581), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U751 ( .A(n581), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U752 ( .A(n580), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U753 ( .A(n580), .B(n418), .ZN(n401) );
  XNOR2_X1 U754 ( .A(n580), .B(n420), .ZN(n403) );
  XNOR2_X1 U755 ( .A(n580), .B(n419), .ZN(n402) );
  XNOR2_X1 U756 ( .A(n580), .B(n421), .ZN(n404) );
  XNOR2_X1 U757 ( .A(n581), .B(n422), .ZN(n405) );
  XNOR2_X1 U758 ( .A(n581), .B(n424), .ZN(n407) );
  XNOR2_X1 U759 ( .A(n581), .B(n423), .ZN(n406) );
  XNOR2_X1 U760 ( .A(n581), .B(n577), .ZN(n408) );
  XNOR2_X1 U761 ( .A(n70), .B(n47), .ZN(product[14]) );
  OAI21_X1 U762 ( .B1(n71), .B2(n553), .A(n72), .ZN(n70) );
  INV_X1 U763 ( .A(n122), .ZN(n120) );
  NAND2_X1 U764 ( .A1(n329), .A2(n258), .ZN(n122) );
  OAI22_X1 U765 ( .A1(n562), .A2(n533), .B1(n409), .B2(n579), .ZN(n258) );
  XOR2_X1 U766 ( .A(n514), .B(n54), .Z(product[7]) );
  OAI22_X1 U767 ( .A1(n379), .A2(n539), .B1(n378), .B2(n536), .ZN(n301) );
  OAI22_X1 U768 ( .A1(n508), .A2(n380), .B1(n379), .B2(n527), .ZN(n302) );
  OAI22_X1 U769 ( .A1(n508), .A2(n385), .B1(n384), .B2(n527), .ZN(n307) );
  OAI22_X1 U770 ( .A1(n508), .A2(n382), .B1(n381), .B2(n521), .ZN(n304) );
  OAI22_X1 U771 ( .A1(n539), .A2(n381), .B1(n380), .B2(n521), .ZN(n303) );
  NAND2_X1 U772 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U773 ( .A1(n540), .A2(n383), .B1(n382), .B2(n521), .ZN(n305) );
  OAI22_X1 U774 ( .A1(n540), .A2(n384), .B1(n383), .B2(n575), .ZN(n306) );
  OAI22_X1 U775 ( .A1(n539), .A2(n386), .B1(n385), .B2(n575), .ZN(n308) );
  OAI22_X1 U776 ( .A1(n508), .A2(n387), .B1(n386), .B2(n521), .ZN(n309) );
  OAI22_X1 U777 ( .A1(n500), .A2(n528), .B1(n392), .B2(n536), .ZN(n257) );
  OAI22_X1 U778 ( .A1(n540), .A2(n389), .B1(n388), .B2(n575), .ZN(n311) );
  OAI22_X1 U779 ( .A1(n539), .A2(n388), .B1(n387), .B2(n575), .ZN(n310) );
  OAI22_X1 U780 ( .A1(n539), .A2(n390), .B1(n389), .B2(n521), .ZN(n312) );
  INV_X1 U781 ( .A(n575), .ZN(n247) );
  OAI22_X1 U782 ( .A1(n508), .A2(n391), .B1(n390), .B2(n575), .ZN(n313) );
  INV_X1 U783 ( .A(n586), .ZN(n585) );
  INV_X1 U784 ( .A(n31), .ZN(n592) );
  INV_X1 U785 ( .A(n36), .ZN(n594) );
  INV_X1 U786 ( .A(n596), .ZN(n595) );
  INV_X1 U787 ( .A(n40), .ZN(n596) );
  XOR2_X1 U788 ( .A(n259), .B(n251), .Z(n148) );
  XOR2_X1 U789 ( .A(n289), .B(n279), .Z(n146) );
  XOR2_X1 U790 ( .A(n149), .B(n147), .Z(n144) );
  XOR2_X1 U791 ( .A(n159), .B(n150), .Z(n142) );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_2_DW01_add_2 ( A, B, CI, 
        SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n8, n9, n10, n11, n12, n13, n14, n15, n16, n19, n20,
         n22, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n44, n45, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n65, n67, n68, n69, n70, n71, n73,
         n75, n76, n77, n78, n79, n81, n83, n84, n86, n88, n89, n90, n95, n96,
         n98, n100, n157, n158, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182;

  AOI21_X2 U122 ( .B1(n181), .B2(n68), .A(n65), .ZN(n63) );
  NOR2_X1 U123 ( .A1(A[8]), .A2(B[8]), .ZN(n157) );
  XNOR2_X1 U124 ( .A(n165), .B(n158), .ZN(SUM[11]) );
  AND2_X1 U125 ( .A1(n164), .A2(n36), .ZN(n158) );
  BUF_X1 U126 ( .A(n37), .Z(n165) );
  AND2_X1 U127 ( .A1(n176), .A2(n86), .ZN(SUM[0]) );
  OR2_X1 U128 ( .A1(A[15]), .A2(B[15]), .ZN(n160) );
  AND2_X1 U129 ( .A1(A[10]), .A2(B[10]), .ZN(n167) );
  INV_X1 U130 ( .A(n167), .ZN(n44) );
  NOR2_X1 U131 ( .A1(A[8]), .A2(B[8]), .ZN(n54) );
  OR2_X1 U132 ( .A1(A[8]), .A2(B[8]), .ZN(n161) );
  XNOR2_X1 U133 ( .A(n45), .B(n162), .ZN(SUM[10]) );
  AND2_X1 U134 ( .A1(n178), .A2(n44), .ZN(n162) );
  CLKBUF_X1 U135 ( .A(n29), .Z(n163) );
  OR2_X1 U136 ( .A1(A[11]), .A2(B[11]), .ZN(n164) );
  AOI21_X1 U137 ( .B1(n52), .B2(n60), .A(n53), .ZN(n166) );
  AOI21_X1 U138 ( .B1(n52), .B2(n60), .A(n53), .ZN(n51) );
  OR2_X2 U139 ( .A1(A[10]), .A2(B[10]), .ZN(n178) );
  AND2_X1 U140 ( .A1(A[9]), .A2(B[9]), .ZN(n168) );
  NOR2_X1 U141 ( .A1(A[12]), .A2(B[12]), .ZN(n169) );
  NOR2_X1 U142 ( .A1(A[12]), .A2(B[12]), .ZN(n32) );
  NOR2_X1 U143 ( .A1(A[14]), .A2(B[14]), .ZN(n170) );
  NOR2_X1 U144 ( .A1(A[14]), .A2(B[14]), .ZN(n25) );
  AOI21_X1 U145 ( .B1(n178), .B2(n168), .A(n167), .ZN(n171) );
  OAI21_X1 U146 ( .B1(n32), .B2(n36), .A(n33), .ZN(n172) );
  OAI21_X1 U147 ( .B1(n39), .B2(n166), .A(n40), .ZN(n173) );
  AOI21_X1 U148 ( .B1(n173), .B2(n30), .A(n172), .ZN(n174) );
  AOI21_X1 U149 ( .B1(n173), .B2(n30), .A(n31), .ZN(n175) );
  OR2_X1 U150 ( .A1(A[0]), .A2(B[0]), .ZN(n176) );
  INV_X1 U151 ( .A(n60), .ZN(n59) );
  INV_X1 U152 ( .A(n51), .ZN(n50) );
  OAI21_X1 U153 ( .B1(n71), .B2(n69), .A(n70), .ZN(n68) );
  AOI21_X1 U154 ( .B1(n182), .B2(n76), .A(n73), .ZN(n71) );
  INV_X1 U155 ( .A(n75), .ZN(n73) );
  AOI21_X1 U156 ( .B1(n180), .B2(n84), .A(n81), .ZN(n79) );
  INV_X1 U157 ( .A(n83), .ZN(n81) );
  INV_X1 U158 ( .A(n67), .ZN(n65) );
  OR2_X1 U159 ( .A1(n170), .A2(n28), .ZN(n177) );
  OAI21_X1 U160 ( .B1(n79), .B2(n77), .A(n78), .ZN(n76) );
  AOI21_X1 U161 ( .B1(n50), .B2(n179), .A(n168), .ZN(n45) );
  NAND2_X1 U162 ( .A1(n161), .A2(n55), .ZN(n9) );
  INV_X1 U163 ( .A(n86), .ZN(n84) );
  OAI21_X1 U164 ( .B1(n59), .B2(n57), .A(n58), .ZN(n56) );
  INV_X1 U165 ( .A(n28), .ZN(n89) );
  NAND2_X1 U166 ( .A1(n182), .A2(n75), .ZN(n14) );
  NAND2_X1 U167 ( .A1(n95), .A2(n58), .ZN(n10) );
  INV_X1 U168 ( .A(n57), .ZN(n95) );
  NAND2_X1 U169 ( .A1(n179), .A2(n49), .ZN(n8) );
  NAND2_X1 U170 ( .A1(n100), .A2(n78), .ZN(n15) );
  INV_X1 U171 ( .A(n77), .ZN(n100) );
  NAND2_X1 U172 ( .A1(n181), .A2(n67), .ZN(n12) );
  NAND2_X1 U173 ( .A1(n180), .A2(n83), .ZN(n16) );
  NAND2_X1 U174 ( .A1(n98), .A2(n70), .ZN(n13) );
  INV_X1 U175 ( .A(n69), .ZN(n98) );
  NAND2_X1 U176 ( .A1(n96), .A2(n62), .ZN(n11) );
  INV_X1 U177 ( .A(n61), .ZN(n96) );
  XNOR2_X1 U178 ( .A(n34), .B(n5), .ZN(SUM[12]) );
  NAND2_X1 U179 ( .A1(n90), .A2(n33), .ZN(n5) );
  XNOR2_X1 U180 ( .A(n50), .B(n8), .ZN(SUM[9]) );
  XOR2_X1 U181 ( .A(n59), .B(n10), .Z(SUM[7]) );
  XNOR2_X1 U182 ( .A(n14), .B(n76), .ZN(SUM[3]) );
  XOR2_X1 U183 ( .A(n15), .B(n79), .Z(SUM[2]) );
  NOR2_X1 U184 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  NOR2_X1 U185 ( .A1(A[11]), .A2(B[11]), .ZN(n35) );
  NOR2_X1 U186 ( .A1(A[7]), .A2(B[7]), .ZN(n57) );
  OR2_X1 U187 ( .A1(A[9]), .A2(B[9]), .ZN(n179) );
  NOR2_X1 U188 ( .A1(A[2]), .A2(B[2]), .ZN(n77) );
  NAND2_X1 U189 ( .A1(n88), .A2(n26), .ZN(n3) );
  NAND2_X1 U190 ( .A1(A[11]), .A2(B[11]), .ZN(n36) );
  OR2_X1 U191 ( .A1(A[1]), .A2(B[1]), .ZN(n180) );
  NOR2_X1 U192 ( .A1(A[4]), .A2(B[4]), .ZN(n69) );
  NAND2_X1 U193 ( .A1(A[12]), .A2(B[12]), .ZN(n33) );
  XNOR2_X1 U194 ( .A(n56), .B(n9), .ZN(SUM[8]) );
  XNOR2_X1 U195 ( .A(n16), .B(n84), .ZN(SUM[1]) );
  NOR2_X1 U196 ( .A1(A[6]), .A2(B[6]), .ZN(n61) );
  NAND2_X1 U197 ( .A1(A[7]), .A2(B[7]), .ZN(n58) );
  OR2_X1 U198 ( .A1(A[5]), .A2(B[5]), .ZN(n181) );
  NAND2_X1 U199 ( .A1(A[2]), .A2(B[2]), .ZN(n78) );
  OR2_X1 U200 ( .A1(A[3]), .A2(B[3]), .ZN(n182) );
  NAND2_X1 U201 ( .A1(A[15]), .A2(B[15]), .ZN(n19) );
  NAND2_X1 U202 ( .A1(A[9]), .A2(B[9]), .ZN(n49) );
  NAND2_X1 U203 ( .A1(A[5]), .A2(B[5]), .ZN(n67) );
  NAND2_X1 U204 ( .A1(A[1]), .A2(B[1]), .ZN(n83) );
  NAND2_X1 U205 ( .A1(A[0]), .A2(B[0]), .ZN(n86) );
  NAND2_X1 U206 ( .A1(A[4]), .A2(B[4]), .ZN(n70) );
  NAND2_X1 U207 ( .A1(A[6]), .A2(B[6]), .ZN(n62) );
  XNOR2_X1 U208 ( .A(n12), .B(n68), .ZN(SUM[5]) );
  NAND2_X1 U209 ( .A1(n89), .A2(n29), .ZN(n4) );
  NAND2_X1 U210 ( .A1(A[13]), .A2(B[13]), .ZN(n29) );
  XOR2_X1 U211 ( .A(n13), .B(n71), .Z(SUM[4]) );
  XOR2_X1 U212 ( .A(n11), .B(n63), .Z(SUM[6]) );
  OAI21_X1 U213 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  XNOR2_X1 U214 ( .A(n20), .B(n2), .ZN(SUM[15]) );
  NAND2_X1 U215 ( .A1(n160), .A2(n19), .ZN(n2) );
  INV_X1 U216 ( .A(n170), .ZN(n88) );
  OAI21_X1 U217 ( .B1(n25), .B2(n29), .A(n26), .ZN(n24) );
  NAND2_X1 U218 ( .A1(A[14]), .A2(B[14]), .ZN(n26) );
  OAI21_X1 U219 ( .B1(n37), .B2(n35), .A(n36), .ZN(n34) );
  OAI21_X1 U220 ( .B1(n169), .B2(n36), .A(n33), .ZN(n31) );
  NOR2_X1 U221 ( .A1(n32), .A2(n35), .ZN(n30) );
  INV_X1 U222 ( .A(n169), .ZN(n90) );
  NAND2_X1 U223 ( .A1(A[3]), .A2(B[3]), .ZN(n75) );
  INV_X1 U224 ( .A(n38), .ZN(n37) );
  NAND2_X1 U225 ( .A1(n178), .A2(n179), .ZN(n39) );
  OAI21_X1 U226 ( .B1(n39), .B2(n166), .A(n171), .ZN(n38) );
  AOI21_X1 U227 ( .B1(n178), .B2(n168), .A(n167), .ZN(n40) );
  NOR2_X1 U228 ( .A1(n157), .A2(n57), .ZN(n52) );
  OAI21_X1 U229 ( .B1(n54), .B2(n58), .A(n55), .ZN(n53) );
  NAND2_X1 U230 ( .A1(A[8]), .A2(B[8]), .ZN(n55) );
  INV_X1 U231 ( .A(n24), .ZN(n22) );
  XNOR2_X1 U232 ( .A(n27), .B(n3), .ZN(SUM[14]) );
  XOR2_X1 U233 ( .A(n174), .B(n4), .Z(SUM[13]) );
  OAI21_X1 U234 ( .B1(n175), .B2(n28), .A(n163), .ZN(n27) );
  OAI21_X1 U235 ( .B1(n174), .B2(n177), .A(n22), .ZN(n20) );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_2 ( clk, clear_acc, 
        data_out_x, data_out, data_out_w, data_out_b, wr_en_y, m_valid, 
        m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [4:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
         N39, N40, N41, N42, N43, N44, n1, n2, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n85, n102, n111, n112, n113, n114, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n13), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n215), .CK(clk), .Q(n17) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n216), .CK(clk), .Q(n18) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n217), .CK(clk), .Q(n19) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n218), .CK(clk), .Q(n20) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n219), .CK(clk), .Q(n21) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n220), .CK(clk), .Q(n22) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n221), .CK(clk), .Q(n23) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n222), .CK(clk), .Q(n24) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n223), .CK(clk), .Q(n25) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n224), .CK(clk), .Q(n26) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n225), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n226), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n227), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n228), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n229), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n230), .CK(clk), .Q(n35) );
  DFF_X1 \f_reg[0]  ( .D(n83), .CK(clk), .Q(f[0]), .QN(n204) );
  DFF_X1 \f_reg[1]  ( .D(n82), .CK(clk), .Q(f[1]), .QN(n205) );
  DFF_X1 \f_reg[2]  ( .D(n81), .CK(clk), .Q(f[2]), .QN(n206) );
  DFF_X1 \f_reg[8]  ( .D(n75), .CK(clk), .Q(f[8]), .QN(n208) );
  DFF_X1 \f_reg[9]  ( .D(n74), .CK(clk), .Q(f[9]), .QN(n209) );
  DFF_X1 \f_reg[10]  ( .D(n73), .CK(clk), .Q(n46), .QN(n210) );
  DFF_X1 \f_reg[11]  ( .D(n72), .CK(clk), .Q(n44), .QN(n211) );
  DFF_X1 \f_reg[12]  ( .D(n71), .CK(clk), .Q(n42), .QN(n212) );
  DFF_X1 \f_reg[13]  ( .D(n70), .CK(clk), .Q(n40), .QN(n213) );
  DFF_X1 \f_reg[14]  ( .D(n1), .CK(clk), .Q(n39), .QN(n214) );
  DFF_X1 \f_reg[15]  ( .D(n2), .CK(clk), .Q(f[15]), .QN(n67) );
  DFF_X1 \data_out_reg[4]  ( .D(n167), .CK(clk), .Q(data_out[4]), .QN(n176) );
  DFF_X1 \data_out_reg[3]  ( .D(n168), .CK(clk), .Q(data_out[3]), .QN(n175) );
  DFF_X1 \data_out_reg[2]  ( .D(n169), .CK(clk), .Q(data_out[2]), .QN(n174) );
  DFF_X1 \data_out_reg[1]  ( .D(n170), .CK(clk), .Q(data_out[1]), .QN(n173) );
  DFF_X1 \data_out_reg[0]  ( .D(n171), .CK(clk), .Q(data_out[0]), .QN(n172) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_2_DW_mult_tc_1 mult_2021 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_2_DW01_add_2 add_2022 ( .A({n194, 
        n193, n192, n191, n190, n189, n203, n202, n201, n200, n199, n198, n197, 
        n196, n195, n188}), .B({f[15], n39, n40, n42, n44, n46, f[9:0]}), .CI(
        1'b0), .SUM(adder) );
  DFF_X1 \data_out_reg[15]  ( .D(n102), .CK(clk), .Q(data_out[15]), .QN(n187)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n111), .CK(clk), .Q(data_out[14]), .QN(n186)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n112), .CK(clk), .Q(data_out[13]), .QN(n185)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n113), .CK(clk), .Q(data_out[12]), .QN(n184)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n114), .CK(clk), .Q(data_out[11]), .QN(n183)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n161), .CK(clk), .Q(data_out[10]), .QN(n182)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n162), .CK(clk), .Q(data_out[9]), .QN(n181) );
  DFF_X1 \data_out_reg[8]  ( .D(n163), .CK(clk), .Q(data_out[8]), .QN(n180) );
  DFF_X1 \data_out_reg[7]  ( .D(n164), .CK(clk), .Q(data_out[7]), .QN(n179) );
  DFF_X1 \data_out_reg[6]  ( .D(n165), .CK(clk), .Q(data_out[6]), .QN(n178) );
  DFF_X1 \data_out_reg[5]  ( .D(n166), .CK(clk), .Q(data_out[5]), .QN(n177) );
  DFF_X1 \f_reg[3]  ( .D(n80), .CK(clk), .Q(f[3]), .QN(n59) );
  DFF_X1 \f_reg[4]  ( .D(n79), .CK(clk), .Q(f[4]), .QN(n60) );
  DFF_X1 \f_reg[5]  ( .D(n78), .CK(clk), .Q(f[5]), .QN(n61) );
  DFF_X1 \f_reg[6]  ( .D(n77), .CK(clk), .Q(f[6]), .QN(n62) );
  DFF_X1 \f_reg[7]  ( .D(n76), .CK(clk), .Q(f[7]), .QN(n207) );
  DFF_X2 delay_reg ( .D(n85), .CK(clk), .Q(n4), .QN(n231) );
  MUX2_X2 U3 ( .A(N39), .B(n22), .S(n4), .Z(n189) );
  AND2_X1 U4 ( .A1(n38), .A2(n14), .ZN(n11) );
  NAND3_X1 U5 ( .A1(n9), .A2(n8), .A3(n10), .ZN(n1) );
  MUX2_X2 U6 ( .A(n21), .B(N40), .S(n231), .Z(n190) );
  NAND3_X1 U8 ( .A1(n5), .A2(n6), .A3(n7), .ZN(n2) );
  MUX2_X2 U9 ( .A(n19), .B(N42), .S(n231), .Z(n192) );
  MUX2_X2 U10 ( .A(n23), .B(N38), .S(n231), .Z(n203) );
  MUX2_X2 U11 ( .A(n24), .B(N37), .S(n231), .Z(n202) );
  MUX2_X2 U12 ( .A(n20), .B(N41), .S(n231), .Z(n191) );
  MUX2_X2 U13 ( .A(n18), .B(N43), .S(n231), .Z(n193) );
  NAND2_X1 U14 ( .A1(data_out_b[15]), .A2(n13), .ZN(n5) );
  NAND2_X1 U15 ( .A1(adder[15]), .A2(n11), .ZN(n6) );
  NAND2_X1 U16 ( .A1(n57), .A2(f[15]), .ZN(n7) );
  NAND2_X1 U17 ( .A1(data_out_b[14]), .A2(n13), .ZN(n8) );
  NAND2_X1 U18 ( .A1(adder[14]), .A2(n11), .ZN(n9) );
  NAND2_X1 U19 ( .A1(n57), .A2(n39), .ZN(n10) );
  INV_X1 U20 ( .A(n14), .ZN(n13) );
  NAND2_X1 U21 ( .A1(n85), .A2(n12), .ZN(n233) );
  INV_X1 U22 ( .A(n38), .ZN(n57) );
  INV_X1 U23 ( .A(clear_acc), .ZN(n14) );
  OAI22_X1 U24 ( .A1(n175), .A2(n233), .B1(n59), .B2(n232), .ZN(n168) );
  OAI22_X1 U25 ( .A1(n176), .A2(n233), .B1(n60), .B2(n232), .ZN(n167) );
  OAI22_X1 U26 ( .A1(n177), .A2(n233), .B1(n61), .B2(n232), .ZN(n166) );
  OAI22_X1 U27 ( .A1(n178), .A2(n233), .B1(n62), .B2(n232), .ZN(n165) );
  OAI22_X1 U28 ( .A1(n179), .A2(n233), .B1(n207), .B2(n232), .ZN(n164) );
  OAI22_X1 U29 ( .A1(n180), .A2(n233), .B1(n208), .B2(n232), .ZN(n163) );
  OAI22_X1 U30 ( .A1(n181), .A2(n233), .B1(n209), .B2(n232), .ZN(n162) );
  INV_X1 U31 ( .A(n16), .ZN(n34) );
  MUX2_X1 U32 ( .A(n29), .B(N32), .S(n231), .Z(n197) );
  INV_X1 U33 ( .A(wr_en_y), .ZN(n12) );
  INV_X1 U34 ( .A(m_ready), .ZN(n15) );
  NAND2_X1 U35 ( .A1(m_valid), .A2(n15), .ZN(n36) );
  OAI21_X1 U36 ( .B1(sel[4]), .B2(n69), .A(n36), .ZN(n85) );
  NAND2_X1 U37 ( .A1(clear_acc_delay), .A2(n231), .ZN(n16) );
  MUX2_X1 U38 ( .A(n17), .B(N44), .S(n34), .Z(n215) );
  MUX2_X1 U39 ( .A(n17), .B(N44), .S(n231), .Z(n194) );
  MUX2_X1 U40 ( .A(n18), .B(N43), .S(n34), .Z(n216) );
  MUX2_X1 U41 ( .A(n19), .B(N42), .S(n34), .Z(n217) );
  MUX2_X1 U42 ( .A(n20), .B(N41), .S(n34), .Z(n218) );
  MUX2_X1 U43 ( .A(n21), .B(N40), .S(n34), .Z(n219) );
  MUX2_X1 U44 ( .A(n22), .B(N39), .S(n34), .Z(n220) );
  MUX2_X1 U45 ( .A(n23), .B(N38), .S(n34), .Z(n221) );
  MUX2_X1 U46 ( .A(n24), .B(N37), .S(n34), .Z(n222) );
  MUX2_X1 U47 ( .A(n25), .B(N36), .S(n34), .Z(n223) );
  MUX2_X1 U48 ( .A(n25), .B(N36), .S(n231), .Z(n201) );
  MUX2_X1 U49 ( .A(n26), .B(N35), .S(n34), .Z(n224) );
  MUX2_X1 U50 ( .A(n26), .B(N35), .S(n231), .Z(n200) );
  MUX2_X1 U51 ( .A(n27), .B(N34), .S(n34), .Z(n225) );
  MUX2_X1 U52 ( .A(n27), .B(N34), .S(n231), .Z(n199) );
  MUX2_X1 U53 ( .A(n28), .B(N33), .S(n34), .Z(n226) );
  MUX2_X1 U54 ( .A(n28), .B(N33), .S(n231), .Z(n198) );
  MUX2_X1 U55 ( .A(n29), .B(N32), .S(n34), .Z(n227) );
  MUX2_X1 U56 ( .A(n32), .B(N31), .S(n34), .Z(n228) );
  MUX2_X1 U57 ( .A(n32), .B(N31), .S(n231), .Z(n196) );
  MUX2_X1 U58 ( .A(n33), .B(N30), .S(n34), .Z(n229) );
  MUX2_X1 U59 ( .A(n33), .B(N30), .S(n231), .Z(n195) );
  MUX2_X1 U60 ( .A(n35), .B(N29), .S(n34), .Z(n230) );
  MUX2_X1 U61 ( .A(n35), .B(N29), .S(n231), .Z(n188) );
  INV_X1 U62 ( .A(n36), .ZN(n37) );
  OAI21_X1 U63 ( .B1(n37), .B2(n4), .A(n14), .ZN(n38) );
  AOI222_X1 U64 ( .A1(data_out_b[13]), .A2(n13), .B1(adder[13]), .B2(n11), 
        .C1(n57), .C2(n40), .ZN(n41) );
  INV_X1 U65 ( .A(n41), .ZN(n70) );
  AOI222_X1 U66 ( .A1(data_out_b[12]), .A2(n13), .B1(adder[12]), .B2(n11), 
        .C1(n57), .C2(n42), .ZN(n43) );
  INV_X1 U67 ( .A(n43), .ZN(n71) );
  AOI222_X1 U68 ( .A1(data_out_b[11]), .A2(n13), .B1(adder[11]), .B2(n11), 
        .C1(n57), .C2(n44), .ZN(n45) );
  INV_X1 U69 ( .A(n45), .ZN(n72) );
  AOI222_X1 U70 ( .A1(data_out_b[10]), .A2(n13), .B1(adder[10]), .B2(n11), 
        .C1(n57), .C2(n46), .ZN(n47) );
  INV_X1 U71 ( .A(n47), .ZN(n73) );
  AOI222_X1 U72 ( .A1(data_out_b[8]), .A2(n13), .B1(adder[8]), .B2(n11), .C1(
        n57), .C2(f[8]), .ZN(n48) );
  INV_X1 U73 ( .A(n48), .ZN(n75) );
  AOI222_X1 U74 ( .A1(data_out_b[7]), .A2(n13), .B1(adder[7]), .B2(n11), .C1(
        n57), .C2(f[7]), .ZN(n49) );
  INV_X1 U75 ( .A(n49), .ZN(n76) );
  AOI222_X1 U76 ( .A1(data_out_b[6]), .A2(n13), .B1(adder[6]), .B2(n11), .C1(
        n57), .C2(f[6]), .ZN(n50) );
  INV_X1 U77 ( .A(n50), .ZN(n77) );
  AOI222_X1 U78 ( .A1(data_out_b[5]), .A2(n13), .B1(adder[5]), .B2(n11), .C1(
        n57), .C2(f[5]), .ZN(n51) );
  INV_X1 U79 ( .A(n51), .ZN(n78) );
  AOI222_X1 U80 ( .A1(data_out_b[4]), .A2(n13), .B1(adder[4]), .B2(n11), .C1(
        n57), .C2(f[4]), .ZN(n52) );
  INV_X1 U81 ( .A(n52), .ZN(n79) );
  AOI222_X1 U82 ( .A1(data_out_b[3]), .A2(n13), .B1(adder[3]), .B2(n11), .C1(
        n57), .C2(f[3]), .ZN(n53) );
  INV_X1 U83 ( .A(n53), .ZN(n80) );
  AOI222_X1 U84 ( .A1(data_out_b[2]), .A2(n13), .B1(adder[2]), .B2(n11), .C1(
        n57), .C2(f[2]), .ZN(n54) );
  INV_X1 U85 ( .A(n54), .ZN(n81) );
  AOI222_X1 U86 ( .A1(data_out_b[1]), .A2(n13), .B1(adder[1]), .B2(n11), .C1(
        n57), .C2(f[1]), .ZN(n55) );
  INV_X1 U87 ( .A(n55), .ZN(n82) );
  AOI222_X1 U88 ( .A1(data_out_b[0]), .A2(n13), .B1(adder[0]), .B2(n11), .C1(
        n57), .C2(f[0]), .ZN(n56) );
  INV_X1 U89 ( .A(n56), .ZN(n83) );
  AOI222_X1 U90 ( .A1(data_out_b[9]), .A2(n13), .B1(adder[9]), .B2(n11), .C1(
        n57), .C2(f[9]), .ZN(n58) );
  INV_X1 U91 ( .A(n58), .ZN(n74) );
  NOR4_X1 U92 ( .A1(n44), .A2(n42), .A3(n40), .A4(n39), .ZN(n66) );
  NOR4_X1 U93 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n46), .ZN(n65) );
  NAND4_X1 U94 ( .A1(n62), .A2(n61), .A3(n60), .A4(n59), .ZN(n63) );
  NOR4_X1 U95 ( .A1(n63), .A2(f[0]), .A3(f[1]), .A4(f[2]), .ZN(n64) );
  NAND3_X1 U96 ( .A1(n66), .A2(n65), .A3(n64), .ZN(n68) );
  NAND3_X1 U97 ( .A1(wr_en_y), .A2(n68), .A3(n67), .ZN(n232) );
  OAI22_X1 U98 ( .A1(n172), .A2(n233), .B1(n204), .B2(n232), .ZN(n171) );
  OAI22_X1 U99 ( .A1(n173), .A2(n233), .B1(n205), .B2(n232), .ZN(n170) );
  OAI22_X1 U100 ( .A1(n174), .A2(n233), .B1(n206), .B2(n232), .ZN(n169) );
  OAI22_X1 U101 ( .A1(n182), .A2(n233), .B1(n210), .B2(n232), .ZN(n161) );
  OAI22_X1 U102 ( .A1(n183), .A2(n233), .B1(n211), .B2(n232), .ZN(n114) );
  OAI22_X1 U103 ( .A1(n184), .A2(n233), .B1(n212), .B2(n232), .ZN(n113) );
  OAI22_X1 U104 ( .A1(n185), .A2(n233), .B1(n213), .B2(n232), .ZN(n112) );
  OAI22_X1 U105 ( .A1(n186), .A2(n233), .B1(n214), .B2(n232), .ZN(n111) );
  OAI22_X1 U106 ( .A1(n187), .A2(n233), .B1(n67), .B2(n232), .ZN(n102) );
  AND4_X1 U107 ( .A1(sel[3]), .A2(sel[2]), .A3(sel[1]), .A4(sel[0]), .ZN(n69)
         );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_1_DW_mult_tc_1 ( a, b, 
        product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n6, n7, n9, n12, n13, n16, n18, n19, n23, n25, n27, n29, n31, n32,
         n34, n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n50, n53,
         n55, n56, n57, n58, n59, n62, n63, n64, n65, n67, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n93, n95, n96, n97, n98, n99, n103, n104,
         n105, n106, n107, n109, n111, n112, n113, n114, n115, n117, n119,
         n120, n122, n125, n128, n135, n139, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n247, n249, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n418, n419, n420,
         n421, n422, n423, n424, n426, n427, n428, n429, n432, n433, n490,
         n491, n492, n493, n494, n495, n496, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n36 = a[13];
  assign n40 = a[15];
  assign n43 = b[0];
  assign n249 = a[0];
  assign n418 = b[7];
  assign n419 = b[6];
  assign n420 = b[5];
  assign n421 = b[4];
  assign n422 = b[3];
  assign n423 = b[2];
  assign n424 = b[1];

  XOR2_X1 U146 ( .A(n161), .B(n142), .Z(n143) );
  XOR2_X1 U148 ( .A(n265), .B(n144), .Z(n145) );
  XOR2_X1 U150 ( .A(n271), .B(n146), .Z(n147) );
  XOR2_X1 U152 ( .A(n301), .B(n148), .Z(n149) );
  FA_X1 U155 ( .A(n156), .B(n165), .CI(n154), .CO(n151), .S(n152) );
  FA_X1 U156 ( .A(n158), .B(n160), .CI(n167), .CO(n153), .S(n154) );
  FA_X1 U157 ( .A(n169), .B(n171), .CI(n162), .CO(n155), .S(n156) );
  FA_X1 U158 ( .A(n280), .B(n290), .CI(n173), .CO(n157), .S(n158) );
  FA_X1 U159 ( .A(n266), .B(n302), .CI(n272), .CO(n159), .S(n160) );
  FA_X1 U160 ( .A(n262), .B(n260), .CI(n316), .CO(n161), .S(n162) );
  FA_X1 U162 ( .A(n170), .B(n172), .CI(n179), .CO(n165), .S(n166) );
  FA_X1 U163 ( .A(n183), .B(n174), .CI(n181), .CO(n167), .S(n168) );
  FA_X1 U164 ( .A(n267), .B(n281), .CI(n273), .CO(n169), .S(n170) );
  FA_X1 U165 ( .A(n303), .B(n263), .CI(n291), .CO(n171), .S(n172) );
  HA_X1 U166 ( .A(n317), .B(n252), .CO(n173), .S(n174) );
  FA_X1 U167 ( .A(n180), .B(n187), .CI(n178), .CO(n175), .S(n176) );
  FA_X1 U168 ( .A(n182), .B(n184), .CI(n189), .CO(n177), .S(n178) );
  FA_X1 U169 ( .A(n193), .B(n282), .CI(n191), .CO(n179), .S(n180) );
  FA_X1 U170 ( .A(n268), .B(n292), .CI(n274), .CO(n181), .S(n182) );
  FA_X1 U171 ( .A(n318), .B(n264), .CI(n304), .CO(n183), .S(n184) );
  FA_X1 U172 ( .A(n197), .B(n190), .CI(n188), .CO(n185), .S(n186) );
  FA_X1 U173 ( .A(n199), .B(n201), .CI(n192), .CO(n187), .S(n188) );
  FA_X1 U174 ( .A(n275), .B(n293), .CI(n194), .CO(n189), .S(n190) );
  FA_X1 U175 ( .A(n283), .B(n253), .CI(n305), .CO(n191), .S(n192) );
  HA_X1 U176 ( .A(n269), .B(n319), .CO(n193), .S(n194) );
  FA_X1 U177 ( .A(n205), .B(n200), .CI(n198), .CO(n195), .S(n196) );
  FA_X1 U178 ( .A(n207), .B(n209), .CI(n202), .CO(n197), .S(n198) );
  FA_X1 U179 ( .A(n294), .B(n284), .CI(n276), .CO(n199), .S(n200) );
  FA_X1 U180 ( .A(n306), .B(n270), .CI(n320), .CO(n201), .S(n202) );
  FA_X1 U181 ( .A(n208), .B(n213), .CI(n206), .CO(n203), .S(n204) );
  FA_X1 U182 ( .A(n215), .B(n307), .CI(n210), .CO(n205), .S(n206) );
  FA_X1 U183 ( .A(n295), .B(n285), .CI(n254), .CO(n207), .S(n208) );
  HA_X1 U184 ( .A(n277), .B(n321), .CO(n209), .S(n210) );
  FA_X1 U185 ( .A(n216), .B(n219), .CI(n214), .CO(n211), .S(n212) );
  FA_X1 U186 ( .A(n286), .B(n296), .CI(n221), .CO(n213), .S(n214) );
  FA_X1 U187 ( .A(n322), .B(n278), .CI(n308), .CO(n215), .S(n216) );
  FA_X1 U188 ( .A(n225), .B(n222), .CI(n220), .CO(n217), .S(n218) );
  FA_X1 U189 ( .A(n255), .B(n297), .CI(n309), .CO(n219), .S(n220) );
  HA_X1 U190 ( .A(n323), .B(n287), .CO(n221), .S(n222) );
  FA_X1 U191 ( .A(n229), .B(n298), .CI(n226), .CO(n223), .S(n224) );
  FA_X1 U192 ( .A(n324), .B(n288), .CI(n310), .CO(n225), .S(n226) );
  FA_X1 U193 ( .A(n256), .B(n299), .CI(n230), .CO(n227), .S(n228) );
  HA_X1 U194 ( .A(n325), .B(n311), .CO(n229), .S(n230) );
  FA_X1 U195 ( .A(n312), .B(n300), .CI(n326), .CO(n231), .S(n232) );
  HA_X1 U196 ( .A(n313), .B(n327), .CO(n233), .S(n234) );
  XNOR2_X1 U414 ( .A(n582), .B(a[12]), .ZN(n490) );
  INV_X4 U415 ( .A(n490), .ZN(n531) );
  INV_X1 U416 ( .A(n128), .ZN(n491) );
  INV_X1 U417 ( .A(n568), .ZN(n492) );
  XOR2_X1 U418 ( .A(n177), .B(n168), .Z(n493) );
  XOR2_X1 U419 ( .A(n166), .B(n493), .Z(n164) );
  NAND2_X1 U420 ( .A1(n166), .A2(n177), .ZN(n494) );
  NAND2_X1 U421 ( .A1(n166), .A2(n168), .ZN(n495) );
  NAND2_X1 U422 ( .A1(n177), .A2(n168), .ZN(n496) );
  NAND3_X1 U423 ( .A1(n494), .A2(n495), .A3(n496), .ZN(n163) );
  OR2_X2 U424 ( .A1(n152), .A2(n163), .ZN(n555) );
  INV_X1 U425 ( .A(n506), .ZN(n41) );
  AND2_X1 U426 ( .A1(n498), .A2(n122), .ZN(product[1]) );
  OR2_X1 U427 ( .A1(n329), .A2(n258), .ZN(n498) );
  OR2_X1 U428 ( .A1(n186), .A2(n195), .ZN(n499) );
  OR2_X1 U429 ( .A1(n218), .A2(n223), .ZN(n500) );
  CLKBUF_X1 U430 ( .A(n224), .Z(n501) );
  XNOR2_X1 U431 ( .A(n507), .B(n502), .ZN(product[7]) );
  AND2_X1 U432 ( .A1(n500), .A2(n98), .ZN(n502) );
  CLKBUF_X1 U433 ( .A(n95), .Z(n503) );
  BUF_X1 U434 ( .A(n9), .Z(n512) );
  BUF_X1 U435 ( .A(n9), .Z(n563) );
  BUF_X1 U436 ( .A(n384), .Z(n504) );
  CLKBUF_X1 U437 ( .A(n104), .Z(n505) );
  XNOR2_X1 U438 ( .A(n584), .B(a[14]), .ZN(n506) );
  AOI21_X1 U439 ( .B1(n547), .B2(n505), .A(n548), .ZN(n507) );
  XNOR2_X1 U440 ( .A(n508), .B(n543), .ZN(product[9]) );
  AND2_X1 U441 ( .A1(n526), .A2(n90), .ZN(n508) );
  BUF_X1 U442 ( .A(n546), .Z(n509) );
  BUF_X2 U443 ( .A(n569), .Z(n528) );
  INV_X1 U444 ( .A(n541), .ZN(n510) );
  BUF_X1 U445 ( .A(n9), .Z(n511) );
  BUF_X1 U446 ( .A(n579), .Z(n513) );
  BUF_X1 U447 ( .A(n579), .Z(n514) );
  INV_X1 U448 ( .A(n580), .ZN(n579) );
  XOR2_X1 U449 ( .A(n492), .B(b[11]), .Z(n397) );
  XNOR2_X1 U450 ( .A(n45), .B(n515), .ZN(product[12]) );
  AND2_X1 U451 ( .A1(n540), .A2(n79), .ZN(n515) );
  NOR2_X1 U452 ( .A1(n186), .A2(n195), .ZN(n516) );
  NOR2_X1 U453 ( .A1(n186), .A2(n195), .ZN(n82) );
  INV_X1 U454 ( .A(n13), .ZN(n576) );
  NOR2_X1 U455 ( .A1(n164), .A2(n175), .ZN(n517) );
  INV_X1 U456 ( .A(n551), .ZN(n518) );
  INV_X1 U457 ( .A(n551), .ZN(n519) );
  NOR2_X1 U458 ( .A1(n164), .A2(n175), .ZN(n75) );
  INV_X2 U459 ( .A(n582), .ZN(n581) );
  OR2_X2 U460 ( .A1(n520), .A2(n521), .ZN(n23) );
  XOR2_X1 U461 ( .A(n578), .B(a[6]), .Z(n520) );
  XNOR2_X1 U462 ( .A(n576), .B(a[6]), .ZN(n521) );
  BUF_X1 U463 ( .A(n530), .Z(n525) );
  INV_X1 U464 ( .A(n544), .ZN(n522) );
  INV_X1 U465 ( .A(n544), .ZN(n523) );
  INV_X1 U466 ( .A(n544), .ZN(n27) );
  INV_X2 U467 ( .A(n573), .ZN(n572) );
  XOR2_X1 U468 ( .A(n576), .B(a[4]), .Z(n536) );
  INV_X1 U469 ( .A(n577), .ZN(n524) );
  OR2_X1 U470 ( .A1(n204), .A2(n211), .ZN(n526) );
  XNOR2_X1 U471 ( .A(n582), .B(a[10]), .ZN(n428) );
  CLKBUF_X1 U472 ( .A(n569), .Z(n527) );
  BUF_X2 U473 ( .A(n569), .Z(n529) );
  INV_X1 U474 ( .A(n570), .ZN(n569) );
  XOR2_X1 U475 ( .A(n570), .B(a[2]), .Z(n530) );
  INV_X1 U476 ( .A(n568), .ZN(n532) );
  NAND2_X1 U477 ( .A1(n428), .A2(n32), .ZN(n533) );
  CLKBUF_X1 U478 ( .A(n554), .Z(n534) );
  XOR2_X1 U479 ( .A(n570), .B(a[2]), .Z(n9) );
  OR2_X1 U480 ( .A1(n228), .A2(n231), .ZN(n535) );
  INV_X1 U481 ( .A(n541), .ZN(n32) );
  OR2_X1 U482 ( .A1(n536), .A2(n509), .ZN(n18) );
  OR2_X1 U483 ( .A1(n536), .A2(n546), .ZN(n537) );
  OR2_X1 U484 ( .A1(n536), .A2(n546), .ZN(n538) );
  XNOR2_X1 U485 ( .A(n570), .B(n249), .ZN(n433) );
  XNOR2_X1 U486 ( .A(n88), .B(n539), .ZN(product[10]) );
  NAND2_X1 U487 ( .A1(n128), .A2(n86), .ZN(n539) );
  OR2_X1 U488 ( .A1(n176), .A2(n185), .ZN(n540) );
  XNOR2_X1 U489 ( .A(n580), .B(a[10]), .ZN(n541) );
  INV_X2 U490 ( .A(n249), .ZN(n567) );
  CLKBUF_X1 U491 ( .A(n96), .Z(n542) );
  CLKBUF_X1 U492 ( .A(n91), .Z(n543) );
  INV_X1 U493 ( .A(n19), .ZN(n578) );
  INV_X2 U494 ( .A(n546), .ZN(n16) );
  XNOR2_X1 U495 ( .A(n578), .B(a[8]), .ZN(n544) );
  XNOR2_X1 U496 ( .A(n573), .B(a[2]), .ZN(n432) );
  INV_X1 U497 ( .A(n573), .ZN(n571) );
  OAI21_X1 U498 ( .B1(n89), .B2(n91), .A(n90), .ZN(n545) );
  OAI21_X1 U499 ( .B1(n91), .B2(n89), .A(n90), .ZN(n88) );
  XNOR2_X1 U500 ( .A(n573), .B(a[4]), .ZN(n546) );
  INV_X1 U501 ( .A(n570), .ZN(n568) );
  CLKBUF_X1 U502 ( .A(n560), .Z(n547) );
  INV_X2 U503 ( .A(n578), .ZN(n577) );
  NAND2_X2 U504 ( .A1(n429), .A2(n27), .ZN(n29) );
  AND2_X1 U505 ( .A1(n224), .A2(n227), .ZN(n548) );
  NAND2_X1 U506 ( .A1(n433), .A2(n567), .ZN(n549) );
  NAND2_X1 U507 ( .A1(n433), .A2(n567), .ZN(n550) );
  XNOR2_X1 U508 ( .A(n576), .B(a[6]), .ZN(n551) );
  NAND2_X1 U509 ( .A1(n530), .A2(n432), .ZN(n552) );
  NAND2_X1 U510 ( .A1(n432), .A2(n9), .ZN(n553) );
  AOI21_X1 U511 ( .B1(n545), .B2(n80), .A(n81), .ZN(n554) );
  BUF_X1 U512 ( .A(n43), .Z(n565) );
  NAND2_X1 U513 ( .A1(n555), .A2(n69), .ZN(n47) );
  INV_X1 U514 ( .A(n73), .ZN(n71) );
  INV_X1 U515 ( .A(n69), .ZN(n67) );
  INV_X1 U516 ( .A(n74), .ZN(n72) );
  NAND2_X1 U517 ( .A1(n73), .A2(n555), .ZN(n64) );
  INV_X1 U518 ( .A(n95), .ZN(n93) );
  AOI21_X1 U519 ( .B1(n80), .B2(n545), .A(n81), .ZN(n45) );
  NOR2_X1 U520 ( .A1(n82), .A2(n85), .ZN(n80) );
  OAI21_X1 U521 ( .B1(n516), .B2(n86), .A(n83), .ZN(n81) );
  NAND2_X1 U522 ( .A1(n125), .A2(n76), .ZN(n48) );
  INV_X1 U523 ( .A(n517), .ZN(n125) );
  INV_X1 U524 ( .A(n85), .ZN(n128) );
  NAND2_X1 U525 ( .A1(n556), .A2(n503), .ZN(n53) );
  OAI21_X1 U526 ( .B1(n75), .B2(n79), .A(n76), .ZN(n74) );
  NAND2_X1 U527 ( .A1(n499), .A2(n83), .ZN(n50) );
  NOR2_X1 U528 ( .A1(n517), .A2(n78), .ZN(n73) );
  NAND2_X1 U529 ( .A1(n152), .A2(n163), .ZN(n69) );
  OAI21_X1 U530 ( .B1(n113), .B2(n115), .A(n114), .ZN(n112) );
  NAND2_X1 U531 ( .A1(n535), .A2(n106), .ZN(n56) );
  AOI21_X1 U532 ( .B1(n558), .B2(n120), .A(n117), .ZN(n115) );
  INV_X1 U533 ( .A(n119), .ZN(n117) );
  NOR2_X1 U534 ( .A1(n176), .A2(n185), .ZN(n78) );
  NOR2_X1 U535 ( .A1(n196), .A2(n203), .ZN(n85) );
  NAND2_X1 U536 ( .A1(n560), .A2(n103), .ZN(n55) );
  XOR2_X1 U537 ( .A(n58), .B(n115), .Z(product[3]) );
  NAND2_X1 U538 ( .A1(n135), .A2(n114), .ZN(n58) );
  INV_X1 U539 ( .A(n113), .ZN(n135) );
  XNOR2_X1 U540 ( .A(n63), .B(n46), .ZN(product[15]) );
  NAND2_X1 U541 ( .A1(n559), .A2(n62), .ZN(n46) );
  AOI21_X1 U542 ( .B1(n74), .B2(n555), .A(n67), .ZN(n65) );
  XNOR2_X1 U543 ( .A(n59), .B(n120), .ZN(product[2]) );
  NAND2_X1 U544 ( .A1(n558), .A2(n119), .ZN(n59) );
  XNOR2_X1 U545 ( .A(n57), .B(n112), .ZN(product[4]) );
  NAND2_X1 U546 ( .A1(n557), .A2(n111), .ZN(n57) );
  NAND2_X1 U547 ( .A1(n176), .A2(n185), .ZN(n79) );
  NAND2_X1 U548 ( .A1(n186), .A2(n195), .ZN(n83) );
  NAND2_X1 U549 ( .A1(n164), .A2(n175), .ZN(n76) );
  NAND2_X1 U550 ( .A1(n196), .A2(n203), .ZN(n86) );
  NAND2_X1 U551 ( .A1(n212), .A2(n217), .ZN(n95) );
  NAND2_X1 U552 ( .A1(n204), .A2(n211), .ZN(n90) );
  OR2_X1 U553 ( .A1(n212), .A2(n217), .ZN(n556) );
  OR2_X1 U554 ( .A1(n232), .A2(n233), .ZN(n557) );
  OR2_X1 U555 ( .A1(n328), .A2(n314), .ZN(n558) );
  NOR2_X1 U556 ( .A1(n234), .A2(n257), .ZN(n113) );
  OR2_X1 U557 ( .A1(n151), .A2(n139), .ZN(n559) );
  NAND2_X1 U558 ( .A1(n328), .A2(n314), .ZN(n119) );
  NOR2_X1 U559 ( .A1(n228), .A2(n231), .ZN(n105) );
  NAND2_X1 U560 ( .A1(n228), .A2(n231), .ZN(n106) );
  NAND2_X1 U561 ( .A1(n232), .A2(n233), .ZN(n111) );
  OR2_X1 U562 ( .A1(n224), .A2(n227), .ZN(n560) );
  NAND2_X1 U563 ( .A1(n501), .A2(n227), .ZN(n103) );
  NAND2_X1 U564 ( .A1(n218), .A2(n223), .ZN(n98) );
  XNOR2_X1 U565 ( .A(n581), .B(a[12]), .ZN(n37) );
  OR2_X1 U566 ( .A1(n565), .A2(n573), .ZN(n392) );
  OAI22_X1 U567 ( .A1(n549), .A2(n406), .B1(n405), .B2(n567), .ZN(n327) );
  OAI22_X1 U568 ( .A1(n550), .A2(n407), .B1(n406), .B2(n567), .ZN(n328) );
  OAI22_X1 U569 ( .A1(n549), .A2(n408), .B1(n407), .B2(n567), .ZN(n329) );
  NAND2_X1 U570 ( .A1(n530), .A2(n432), .ZN(n12) );
  NAND2_X1 U571 ( .A1(n433), .A2(n567), .ZN(n6) );
  XNOR2_X1 U572 ( .A(n575), .B(n565), .ZN(n376) );
  AND2_X1 U573 ( .A1(n566), .A2(n509), .ZN(n300) );
  OAI22_X1 U574 ( .A1(n6), .A2(n405), .B1(n404), .B2(n567), .ZN(n326) );
  OAI22_X1 U575 ( .A1(n550), .A2(n400), .B1(n399), .B2(n567), .ZN(n321) );
  XNOR2_X1 U576 ( .A(n514), .B(n565), .ZN(n352) );
  OAI22_X1 U577 ( .A1(n42), .A2(n586), .B1(n332), .B2(n41), .ZN(n251) );
  OR2_X1 U578 ( .A1(n565), .A2(n586), .ZN(n332) );
  OAI22_X1 U579 ( .A1(n404), .A2(n6), .B1(n403), .B2(n567), .ZN(n325) );
  OAI22_X1 U580 ( .A1(n549), .A2(n398), .B1(n397), .B2(n567), .ZN(n319) );
  XNOR2_X1 U581 ( .A(n581), .B(n565), .ZN(n343) );
  XOR2_X1 U582 ( .A(n579), .B(a[8]), .Z(n429) );
  XOR2_X1 U583 ( .A(n315), .B(n261), .Z(n150) );
  OAI22_X1 U584 ( .A1(n550), .A2(n394), .B1(n393), .B2(n567), .ZN(n315) );
  XNOR2_X1 U585 ( .A(n155), .B(n561), .ZN(n139) );
  XNOR2_X1 U586 ( .A(n153), .B(n141), .ZN(n561) );
  XNOR2_X1 U587 ( .A(n157), .B(n562), .ZN(n141) );
  XNOR2_X1 U588 ( .A(n145), .B(n143), .ZN(n562) );
  XNOR2_X1 U589 ( .A(n583), .B(n565), .ZN(n336) );
  NAND2_X1 U590 ( .A1(n427), .A2(n37), .ZN(n39) );
  XOR2_X1 U591 ( .A(n583), .B(a[12]), .Z(n427) );
  OAI22_X1 U592 ( .A1(n39), .A2(n336), .B1(n531), .B2(n335), .ZN(n263) );
  AND2_X1 U593 ( .A1(n566), .A2(n551), .ZN(n288) );
  OAI22_X1 U594 ( .A1(n6), .A2(n403), .B1(n402), .B2(n567), .ZN(n324) );
  AND2_X1 U595 ( .A1(n566), .A2(n541), .ZN(n270) );
  OAI22_X1 U596 ( .A1(n550), .A2(n399), .B1(n398), .B2(n567), .ZN(n320) );
  AND2_X1 U597 ( .A1(n566), .A2(n506), .ZN(n260) );
  OAI22_X1 U598 ( .A1(n549), .A2(n395), .B1(n394), .B2(n567), .ZN(n316) );
  OAI22_X1 U599 ( .A1(n39), .A2(n335), .B1(n531), .B2(n334), .ZN(n262) );
  INV_X1 U600 ( .A(n25), .ZN(n580) );
  AND2_X1 U601 ( .A1(n566), .A2(n544), .ZN(n278) );
  OAI22_X1 U602 ( .A1(n549), .A2(n401), .B1(n400), .B2(n567), .ZN(n322) );
  NAND2_X1 U603 ( .A1(n426), .A2(n41), .ZN(n42) );
  XOR2_X1 U604 ( .A(n585), .B(a[14]), .Z(n426) );
  INV_X1 U605 ( .A(n7), .ZN(n573) );
  OAI22_X1 U606 ( .A1(n549), .A2(n402), .B1(n401), .B2(n567), .ZN(n323) );
  XNOR2_X1 U607 ( .A(n577), .B(n565), .ZN(n363) );
  OAI22_X1 U608 ( .A1(n549), .A2(n396), .B1(n395), .B2(n567), .ZN(n317) );
  OAI22_X1 U609 ( .A1(n39), .A2(n584), .B1(n337), .B2(n531), .ZN(n252) );
  OR2_X1 U610 ( .A1(n565), .A2(n584), .ZN(n337) );
  AND2_X1 U611 ( .A1(n566), .A2(n247), .ZN(n314) );
  OAI22_X1 U612 ( .A1(n550), .A2(n397), .B1(n396), .B2(n567), .ZN(n318) );
  AND2_X1 U613 ( .A1(n566), .A2(n490), .ZN(n264) );
  AND2_X1 U614 ( .A1(n566), .A2(n249), .ZN(product[0]) );
  OR2_X1 U615 ( .A1(n565), .A2(n582), .ZN(n344) );
  OR2_X1 U616 ( .A1(n565), .A2(n524), .ZN(n364) );
  OR2_X1 U617 ( .A1(n565), .A2(n580), .ZN(n353) );
  OR2_X1 U618 ( .A1(n565), .A2(n576), .ZN(n377) );
  XNOR2_X1 U619 ( .A(n577), .B(b[9]), .ZN(n354) );
  OAI22_X1 U620 ( .A1(n39), .A2(n334), .B1(n531), .B2(n333), .ZN(n261) );
  XNOR2_X1 U621 ( .A(n583), .B(n422), .ZN(n333) );
  XNOR2_X1 U622 ( .A(n575), .B(b[11]), .ZN(n365) );
  XNOR2_X1 U623 ( .A(n583), .B(n424), .ZN(n335) );
  XNOR2_X1 U624 ( .A(n583), .B(n423), .ZN(n334) );
  OAI22_X1 U625 ( .A1(n42), .A2(n331), .B1(n330), .B2(n41), .ZN(n259) );
  XNOR2_X1 U626 ( .A(n585), .B(n424), .ZN(n330) );
  XNOR2_X1 U627 ( .A(n585), .B(n565), .ZN(n331) );
  XNOR2_X1 U628 ( .A(n528), .B(b[12]), .ZN(n396) );
  XNOR2_X1 U629 ( .A(n528), .B(b[13]), .ZN(n395) );
  XNOR2_X1 U630 ( .A(n529), .B(b[14]), .ZN(n394) );
  XNOR2_X1 U631 ( .A(n513), .B(n418), .ZN(n345) );
  XNOR2_X1 U632 ( .A(n581), .B(n420), .ZN(n338) );
  XNOR2_X1 U633 ( .A(n572), .B(b[13]), .ZN(n378) );
  XNOR2_X1 U634 ( .A(n581), .B(n424), .ZN(n342) );
  XNOR2_X1 U635 ( .A(n577), .B(n424), .ZN(n362) );
  XNOR2_X1 U636 ( .A(n513), .B(n424), .ZN(n351) );
  XNOR2_X1 U637 ( .A(n581), .B(n423), .ZN(n341) );
  XNOR2_X1 U638 ( .A(n581), .B(n422), .ZN(n340) );
  XNOR2_X1 U639 ( .A(n581), .B(n421), .ZN(n339) );
  XNOR2_X1 U640 ( .A(n571), .B(b[8]), .ZN(n383) );
  XNOR2_X1 U641 ( .A(n572), .B(b[9]), .ZN(n382) );
  XNOR2_X1 U642 ( .A(n572), .B(n418), .ZN(n384) );
  XNOR2_X1 U643 ( .A(n572), .B(n419), .ZN(n385) );
  XNOR2_X1 U644 ( .A(n572), .B(b[10]), .ZN(n381) );
  XNOR2_X1 U645 ( .A(n572), .B(b[11]), .ZN(n380) );
  XNOR2_X1 U646 ( .A(n572), .B(b[12]), .ZN(n379) );
  XNOR2_X1 U647 ( .A(n577), .B(n422), .ZN(n360) );
  XNOR2_X1 U648 ( .A(n514), .B(n422), .ZN(n349) );
  XNOR2_X1 U649 ( .A(n575), .B(b[10]), .ZN(n366) );
  XNOR2_X1 U650 ( .A(n575), .B(n418), .ZN(n369) );
  XNOR2_X1 U651 ( .A(n575), .B(b[8]), .ZN(n368) );
  XNOR2_X1 U652 ( .A(n575), .B(b[9]), .ZN(n367) );
  XNOR2_X1 U653 ( .A(n577), .B(n423), .ZN(n361) );
  XNOR2_X1 U654 ( .A(n513), .B(n423), .ZN(n350) );
  XNOR2_X1 U655 ( .A(n577), .B(n420), .ZN(n358) );
  XNOR2_X1 U656 ( .A(n513), .B(n420), .ZN(n347) );
  XNOR2_X1 U657 ( .A(n577), .B(n421), .ZN(n359) );
  XNOR2_X1 U658 ( .A(n514), .B(n421), .ZN(n348) );
  XNOR2_X1 U659 ( .A(n577), .B(n418), .ZN(n356) );
  XNOR2_X1 U660 ( .A(n577), .B(n419), .ZN(n357) );
  XNOR2_X1 U661 ( .A(n514), .B(n419), .ZN(n346) );
  XNOR2_X1 U662 ( .A(n577), .B(b[8]), .ZN(n355) );
  XNOR2_X1 U663 ( .A(n528), .B(b[15]), .ZN(n393) );
  BUF_X1 U664 ( .A(n43), .Z(n566) );
  OAI22_X1 U665 ( .A1(n533), .A2(n339), .B1(n338), .B2(n510), .ZN(n265) );
  OAI22_X1 U666 ( .A1(n533), .A2(n340), .B1(n339), .B2(n510), .ZN(n266) );
  OAI22_X1 U667 ( .A1(n533), .A2(n341), .B1(n340), .B2(n510), .ZN(n267) );
  OAI22_X1 U668 ( .A1(n533), .A2(n342), .B1(n341), .B2(n510), .ZN(n268) );
  OAI22_X1 U669 ( .A1(n533), .A2(n343), .B1(n342), .B2(n510), .ZN(n269) );
  OAI22_X1 U670 ( .A1(n34), .A2(n582), .B1(n344), .B2(n510), .ZN(n253) );
  NAND2_X1 U671 ( .A1(n428), .A2(n32), .ZN(n34) );
  NOR2_X1 U672 ( .A1(n218), .A2(n223), .ZN(n97) );
  CLKBUF_X1 U673 ( .A(n107), .Z(n564) );
  AOI21_X1 U674 ( .B1(n557), .B2(n112), .A(n109), .ZN(n107) );
  XNOR2_X1 U675 ( .A(n77), .B(n48), .ZN(product[13]) );
  XNOR2_X1 U676 ( .A(n572), .B(n420), .ZN(n386) );
  XNOR2_X1 U677 ( .A(n571), .B(n422), .ZN(n388) );
  XNOR2_X1 U678 ( .A(n572), .B(n565), .ZN(n391) );
  XNOR2_X1 U679 ( .A(n571), .B(n421), .ZN(n387) );
  XNOR2_X1 U680 ( .A(n571), .B(n423), .ZN(n389) );
  XNOR2_X1 U681 ( .A(n571), .B(n424), .ZN(n390) );
  NOR2_X1 U682 ( .A1(n204), .A2(n211), .ZN(n89) );
  OAI22_X1 U683 ( .A1(n29), .A2(n350), .B1(n349), .B2(n522), .ZN(n275) );
  OAI22_X1 U684 ( .A1(n29), .A2(n346), .B1(n345), .B2(n522), .ZN(n271) );
  OAI22_X1 U685 ( .A1(n29), .A2(n348), .B1(n347), .B2(n523), .ZN(n273) );
  OAI22_X1 U686 ( .A1(n29), .A2(n347), .B1(n346), .B2(n523), .ZN(n272) );
  OAI22_X1 U687 ( .A1(n29), .A2(n351), .B1(n350), .B2(n523), .ZN(n276) );
  OAI22_X1 U688 ( .A1(n29), .A2(n349), .B1(n348), .B2(n522), .ZN(n274) );
  OAI22_X1 U689 ( .A1(n29), .A2(n580), .B1(n353), .B2(n523), .ZN(n254) );
  OAI22_X1 U690 ( .A1(n29), .A2(n352), .B1(n351), .B2(n522), .ZN(n277) );
  OAI21_X1 U691 ( .B1(n87), .B2(n491), .A(n86), .ZN(n84) );
  XNOR2_X1 U692 ( .A(n574), .B(n424), .ZN(n375) );
  XNOR2_X1 U693 ( .A(n574), .B(n419), .ZN(n370) );
  XNOR2_X1 U694 ( .A(n574), .B(n420), .ZN(n371) );
  XNOR2_X1 U695 ( .A(n574), .B(n423), .ZN(n374) );
  XNOR2_X1 U696 ( .A(n574), .B(n422), .ZN(n373) );
  XNOR2_X1 U697 ( .A(n574), .B(n421), .ZN(n372) );
  XNOR2_X1 U698 ( .A(n84), .B(n50), .ZN(product[11]) );
  AOI21_X1 U699 ( .B1(n560), .B2(n104), .A(n548), .ZN(n99) );
  OR2_X1 U700 ( .A1(n565), .A2(n532), .ZN(n409) );
  INV_X1 U701 ( .A(n1), .ZN(n570) );
  OAI22_X1 U702 ( .A1(n23), .A2(n356), .B1(n355), .B2(n518), .ZN(n280) );
  OAI22_X1 U703 ( .A1(n23), .A2(n358), .B1(n357), .B2(n519), .ZN(n282) );
  OAI22_X1 U704 ( .A1(n23), .A2(n362), .B1(n361), .B2(n518), .ZN(n286) );
  OAI22_X1 U705 ( .A1(n23), .A2(n360), .B1(n359), .B2(n519), .ZN(n284) );
  OAI22_X1 U706 ( .A1(n23), .A2(n361), .B1(n360), .B2(n519), .ZN(n285) );
  OAI22_X1 U707 ( .A1(n23), .A2(n524), .B1(n364), .B2(n518), .ZN(n255) );
  OAI22_X1 U708 ( .A1(n23), .A2(n355), .B1(n354), .B2(n519), .ZN(n279) );
  OAI22_X1 U709 ( .A1(n23), .A2(n357), .B1(n356), .B2(n518), .ZN(n281) );
  OAI22_X1 U710 ( .A1(n23), .A2(n363), .B1(n362), .B2(n518), .ZN(n287) );
  OAI22_X1 U711 ( .A1(n23), .A2(n359), .B1(n358), .B2(n519), .ZN(n283) );
  XNOR2_X1 U712 ( .A(n529), .B(b[8]), .ZN(n400) );
  XNOR2_X1 U713 ( .A(n527), .B(b[10]), .ZN(n398) );
  XNOR2_X1 U714 ( .A(n527), .B(b[9]), .ZN(n399) );
  XNOR2_X1 U715 ( .A(n529), .B(n418), .ZN(n401) );
  XNOR2_X1 U716 ( .A(n568), .B(n419), .ZN(n402) );
  XNOR2_X1 U717 ( .A(n568), .B(n420), .ZN(n403) );
  XNOR2_X1 U718 ( .A(n529), .B(n421), .ZN(n404) );
  XNOR2_X1 U719 ( .A(n528), .B(n422), .ZN(n405) );
  XNOR2_X1 U720 ( .A(n542), .B(n53), .ZN(product[8]) );
  OAI21_X1 U721 ( .B1(n99), .B2(n97), .A(n98), .ZN(n96) );
  XNOR2_X1 U722 ( .A(n55), .B(n505), .ZN(product[6]) );
  OAI21_X1 U723 ( .B1(n105), .B2(n107), .A(n106), .ZN(n104) );
  NAND2_X1 U724 ( .A1(n151), .A2(n139), .ZN(n62) );
  OAI22_X1 U725 ( .A1(n537), .A2(n370), .B1(n369), .B2(n16), .ZN(n293) );
  OAI22_X1 U726 ( .A1(n537), .A2(n367), .B1(n366), .B2(n16), .ZN(n290) );
  OAI22_X1 U727 ( .A1(n538), .A2(n375), .B1(n374), .B2(n16), .ZN(n298) );
  OAI22_X1 U728 ( .A1(n18), .A2(n372), .B1(n371), .B2(n16), .ZN(n295) );
  OAI22_X1 U729 ( .A1(n537), .A2(n373), .B1(n372), .B2(n16), .ZN(n296) );
  OAI22_X1 U730 ( .A1(n538), .A2(n374), .B1(n373), .B2(n16), .ZN(n297) );
  OAI22_X1 U731 ( .A1(n538), .A2(n368), .B1(n367), .B2(n16), .ZN(n291) );
  OAI22_X1 U732 ( .A1(n537), .A2(n369), .B1(n368), .B2(n16), .ZN(n292) );
  OAI22_X1 U733 ( .A1(n537), .A2(n576), .B1(n377), .B2(n16), .ZN(n256) );
  OAI22_X1 U734 ( .A1(n18), .A2(n371), .B1(n370), .B2(n16), .ZN(n294) );
  OAI22_X1 U735 ( .A1(n538), .A2(n376), .B1(n375), .B2(n16), .ZN(n299) );
  OAI22_X1 U736 ( .A1(n538), .A2(n366), .B1(n365), .B2(n16), .ZN(n289) );
  XNOR2_X1 U737 ( .A(n528), .B(n424), .ZN(n407) );
  XNOR2_X1 U738 ( .A(n529), .B(n423), .ZN(n406) );
  XNOR2_X1 U739 ( .A(n528), .B(n565), .ZN(n408) );
  INV_X1 U740 ( .A(n88), .ZN(n87) );
  XOR2_X1 U741 ( .A(n56), .B(n564), .Z(product[5]) );
  OAI21_X1 U742 ( .B1(n64), .B2(n534), .A(n65), .ZN(n63) );
  XNOR2_X1 U743 ( .A(n70), .B(n47), .ZN(product[14]) );
  OAI21_X1 U744 ( .B1(n554), .B2(n78), .A(n79), .ZN(n77) );
  OAI21_X1 U745 ( .B1(n554), .B2(n71), .A(n72), .ZN(n70) );
  INV_X1 U746 ( .A(n122), .ZN(n120) );
  NAND2_X1 U747 ( .A1(n329), .A2(n258), .ZN(n122) );
  AOI21_X1 U748 ( .B1(n96), .B2(n556), .A(n93), .ZN(n91) );
  INV_X1 U749 ( .A(n111), .ZN(n109) );
  OAI22_X1 U750 ( .A1(n550), .A2(n532), .B1(n409), .B2(n567), .ZN(n258) );
  OAI22_X1 U751 ( .A1(n552), .A2(n379), .B1(n378), .B2(n511), .ZN(n301) );
  OAI22_X1 U752 ( .A1(n552), .A2(n380), .B1(n379), .B2(n525), .ZN(n302) );
  OAI22_X1 U753 ( .A1(n553), .A2(n385), .B1(n504), .B2(n525), .ZN(n307) );
  OAI22_X1 U754 ( .A1(n552), .A2(n382), .B1(n381), .B2(n525), .ZN(n304) );
  OAI22_X1 U755 ( .A1(n552), .A2(n381), .B1(n380), .B2(n511), .ZN(n303) );
  NAND2_X1 U756 ( .A1(n234), .A2(n257), .ZN(n114) );
  OAI22_X1 U757 ( .A1(n553), .A2(n383), .B1(n382), .B2(n512), .ZN(n305) );
  OAI22_X1 U758 ( .A1(n12), .A2(n384), .B1(n525), .B2(n383), .ZN(n306) );
  OAI22_X1 U759 ( .A1(n553), .A2(n386), .B1(n385), .B2(n512), .ZN(n308) );
  OAI22_X1 U760 ( .A1(n552), .A2(n387), .B1(n386), .B2(n511), .ZN(n309) );
  OAI22_X1 U761 ( .A1(n552), .A2(n573), .B1(n392), .B2(n512), .ZN(n257) );
  OAI22_X1 U762 ( .A1(n12), .A2(n389), .B1(n388), .B2(n563), .ZN(n311) );
  OAI22_X1 U763 ( .A1(n12), .A2(n388), .B1(n387), .B2(n563), .ZN(n310) );
  OAI22_X1 U764 ( .A1(n12), .A2(n390), .B1(n389), .B2(n511), .ZN(n312) );
  INV_X1 U765 ( .A(n512), .ZN(n247) );
  OAI22_X1 U766 ( .A1(n553), .A2(n391), .B1(n390), .B2(n511), .ZN(n313) );
  INV_X1 U767 ( .A(n576), .ZN(n574) );
  INV_X1 U768 ( .A(n576), .ZN(n575) );
  INV_X1 U769 ( .A(n31), .ZN(n582) );
  INV_X1 U770 ( .A(n584), .ZN(n583) );
  INV_X1 U771 ( .A(n36), .ZN(n584) );
  INV_X1 U772 ( .A(n586), .ZN(n585) );
  INV_X1 U773 ( .A(n40), .ZN(n586) );
  XOR2_X1 U774 ( .A(n259), .B(n251), .Z(n148) );
  XOR2_X1 U775 ( .A(n289), .B(n279), .Z(n146) );
  XOR2_X1 U776 ( .A(n149), .B(n147), .Z(n144) );
  XOR2_X1 U777 ( .A(n159), .B(n150), .Z(n142) );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_1_DW01_add_2 ( A, B, CI, 
        SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n5, n8, n9, n10, n11, n12, n13, n14, n15, n16, n19, n20, n22,
         n24, n25, n26, n27, n28, n29, n30, n32, n33, n34, n35, n36, n37, n39,
         n40, n44, n45, n47, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n65, n67, n68, n69, n70, n71, n73, n75, n76,
         n77, n78, n79, n81, n83, n84, n86, n91, n94, n95, n96, n98, n100,
         n157, n158, n159, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180;

  AOI21_X1 U122 ( .B1(n52), .B2(n60), .A(n53), .ZN(n157) );
  XNOR2_X1 U123 ( .A(n37), .B(n158), .ZN(SUM[11]) );
  AND2_X1 U124 ( .A1(n91), .A2(n36), .ZN(n158) );
  OR2_X1 U125 ( .A1(A[12]), .A2(B[12]), .ZN(n159) );
  AND2_X1 U126 ( .A1(n173), .A2(n86), .ZN(SUM[0]) );
  OR2_X1 U127 ( .A1(A[15]), .A2(B[15]), .ZN(n161) );
  NOR2_X1 U128 ( .A1(A[8]), .A2(B[8]), .ZN(n162) );
  NOR2_X1 U129 ( .A1(A[8]), .A2(B[8]), .ZN(n54) );
  XNOR2_X1 U130 ( .A(n45), .B(n163), .ZN(SUM[10]) );
  AND2_X1 U131 ( .A1(n170), .A2(n44), .ZN(n163) );
  OAI21_X1 U132 ( .B1(n39), .B2(n51), .A(n40), .ZN(n164) );
  XNOR2_X1 U133 ( .A(n172), .B(n165), .ZN(SUM[13]) );
  AND2_X1 U134 ( .A1(n166), .A2(n29), .ZN(n165) );
  OR2_X1 U135 ( .A1(A[13]), .A2(B[13]), .ZN(n166) );
  CLKBUF_X1 U136 ( .A(n36), .Z(n167) );
  OR2_X1 U137 ( .A1(A[14]), .A2(B[14]), .ZN(n168) );
  OAI21_X1 U138 ( .B1(n32), .B2(n36), .A(n33), .ZN(n169) );
  NOR2_X2 U139 ( .A1(A[11]), .A2(B[11]), .ZN(n35) );
  NOR2_X2 U140 ( .A1(A[12]), .A2(B[12]), .ZN(n32) );
  OR2_X1 U141 ( .A1(A[10]), .A2(B[10]), .ZN(n170) );
  OR2_X1 U142 ( .A1(A[10]), .A2(B[10]), .ZN(n179) );
  AOI21_X1 U143 ( .B1(n164), .B2(n30), .A(n169), .ZN(n171) );
  AOI21_X1 U144 ( .B1(n164), .B2(n30), .A(n169), .ZN(n172) );
  INV_X1 U145 ( .A(n24), .ZN(n22) );
  OR2_X1 U146 ( .A1(A[0]), .A2(B[0]), .ZN(n173) );
  INV_X1 U147 ( .A(n60), .ZN(n59) );
  AOI21_X1 U148 ( .B1(n176), .B2(n84), .A(n81), .ZN(n79) );
  INV_X1 U149 ( .A(n83), .ZN(n81) );
  AOI21_X1 U150 ( .B1(n177), .B2(n68), .A(n65), .ZN(n63) );
  INV_X1 U151 ( .A(n67), .ZN(n65) );
  AOI21_X1 U152 ( .B1(n178), .B2(n76), .A(n73), .ZN(n71) );
  INV_X1 U153 ( .A(n75), .ZN(n73) );
  OR2_X1 U154 ( .A1(n25), .A2(n28), .ZN(n174) );
  OAI21_X1 U155 ( .B1(n79), .B2(n77), .A(n78), .ZN(n76) );
  AOI21_X1 U156 ( .B1(n50), .B2(n175), .A(n47), .ZN(n45) );
  INV_X1 U157 ( .A(n86), .ZN(n84) );
  OAI21_X1 U158 ( .B1(n59), .B2(n57), .A(n58), .ZN(n56) );
  NOR2_X1 U159 ( .A1(n162), .A2(n57), .ZN(n52) );
  OAI21_X1 U160 ( .B1(n54), .B2(n58), .A(n55), .ZN(n53) );
  INV_X1 U161 ( .A(n49), .ZN(n47) );
  NAND2_X1 U162 ( .A1(n95), .A2(n58), .ZN(n10) );
  INV_X1 U163 ( .A(n57), .ZN(n95) );
  NAND2_X1 U164 ( .A1(n94), .A2(n55), .ZN(n9) );
  INV_X1 U165 ( .A(n162), .ZN(n94) );
  INV_X1 U166 ( .A(n35), .ZN(n91) );
  NAND2_X1 U167 ( .A1(n175), .A2(n49), .ZN(n8) );
  NAND2_X1 U168 ( .A1(n100), .A2(n78), .ZN(n15) );
  INV_X1 U169 ( .A(n77), .ZN(n100) );
  NAND2_X1 U170 ( .A1(n177), .A2(n67), .ZN(n12) );
  NAND2_X1 U171 ( .A1(n176), .A2(n83), .ZN(n16) );
  NAND2_X1 U172 ( .A1(n178), .A2(n75), .ZN(n14) );
  NAND2_X1 U173 ( .A1(n96), .A2(n62), .ZN(n11) );
  INV_X1 U174 ( .A(n61), .ZN(n96) );
  NAND2_X1 U175 ( .A1(n98), .A2(n70), .ZN(n13) );
  INV_X1 U176 ( .A(n69), .ZN(n98) );
  XNOR2_X1 U177 ( .A(n50), .B(n8), .ZN(SUM[9]) );
  XNOR2_X1 U178 ( .A(n56), .B(n9), .ZN(SUM[8]) );
  XOR2_X1 U179 ( .A(n59), .B(n10), .Z(SUM[7]) );
  XNOR2_X1 U180 ( .A(n14), .B(n76), .ZN(SUM[3]) );
  NOR2_X1 U181 ( .A1(A[7]), .A2(B[7]), .ZN(n57) );
  NOR2_X1 U182 ( .A1(A[13]), .A2(B[13]), .ZN(n28) );
  NOR2_X1 U183 ( .A1(A[14]), .A2(B[14]), .ZN(n25) );
  OR2_X1 U184 ( .A1(A[9]), .A2(B[9]), .ZN(n175) );
  NOR2_X1 U185 ( .A1(A[2]), .A2(B[2]), .ZN(n77) );
  NAND2_X1 U186 ( .A1(A[11]), .A2(B[11]), .ZN(n36) );
  OR2_X1 U187 ( .A1(A[1]), .A2(B[1]), .ZN(n176) );
  NAND2_X1 U188 ( .A1(A[7]), .A2(B[7]), .ZN(n58) );
  NAND2_X1 U189 ( .A1(A[3]), .A2(B[3]), .ZN(n75) );
  XNOR2_X1 U190 ( .A(n12), .B(n68), .ZN(SUM[5]) );
  XNOR2_X1 U191 ( .A(n27), .B(n3), .ZN(SUM[14]) );
  NAND2_X1 U192 ( .A1(n168), .A2(n26), .ZN(n3) );
  NOR2_X1 U193 ( .A1(A[6]), .A2(B[6]), .ZN(n61) );
  NOR2_X1 U194 ( .A1(A[4]), .A2(B[4]), .ZN(n69) );
  OR2_X1 U195 ( .A1(A[5]), .A2(B[5]), .ZN(n177) );
  OR2_X1 U196 ( .A1(A[3]), .A2(B[3]), .ZN(n178) );
  NAND2_X1 U197 ( .A1(A[8]), .A2(B[8]), .ZN(n55) );
  NAND2_X1 U198 ( .A1(A[2]), .A2(B[2]), .ZN(n78) );
  NAND2_X1 U199 ( .A1(A[9]), .A2(B[9]), .ZN(n49) );
  NAND2_X1 U200 ( .A1(A[1]), .A2(B[1]), .ZN(n83) );
  NAND2_X1 U201 ( .A1(A[5]), .A2(B[5]), .ZN(n67) );
  NAND2_X1 U202 ( .A1(A[0]), .A2(B[0]), .ZN(n86) );
  NAND2_X1 U203 ( .A1(A[4]), .A2(B[4]), .ZN(n70) );
  NAND2_X1 U204 ( .A1(A[6]), .A2(B[6]), .ZN(n62) );
  XOR2_X1 U205 ( .A(n15), .B(n79), .Z(SUM[2]) );
  XNOR2_X1 U206 ( .A(n16), .B(n84), .ZN(SUM[1]) );
  NAND2_X1 U207 ( .A1(n161), .A2(n19), .ZN(n2) );
  NAND2_X1 U208 ( .A1(n159), .A2(n33), .ZN(n5) );
  INV_X1 U209 ( .A(n180), .ZN(n44) );
  AND2_X1 U210 ( .A1(A[10]), .A2(B[10]), .ZN(n180) );
  OAI21_X1 U211 ( .B1(n37), .B2(n35), .A(n167), .ZN(n34) );
  NAND2_X1 U212 ( .A1(A[13]), .A2(B[13]), .ZN(n29) );
  NAND2_X1 U213 ( .A1(A[12]), .A2(B[12]), .ZN(n33) );
  NAND2_X1 U214 ( .A1(A[15]), .A2(B[15]), .ZN(n19) );
  XOR2_X1 U215 ( .A(n13), .B(n71), .Z(SUM[4]) );
  OAI21_X1 U216 ( .B1(n71), .B2(n69), .A(n70), .ZN(n68) );
  INV_X1 U217 ( .A(n157), .ZN(n50) );
  AOI21_X1 U218 ( .B1(n52), .B2(n60), .A(n53), .ZN(n51) );
  OAI21_X1 U219 ( .B1(n25), .B2(n29), .A(n26), .ZN(n24) );
  NAND2_X1 U220 ( .A1(A[14]), .A2(B[14]), .ZN(n26) );
  XOR2_X1 U221 ( .A(n11), .B(n63), .Z(SUM[6]) );
  OAI21_X1 U222 ( .B1(n63), .B2(n61), .A(n62), .ZN(n60) );
  NAND2_X1 U223 ( .A1(n170), .A2(n175), .ZN(n39) );
  AOI21_X1 U224 ( .B1(n179), .B2(n47), .A(n180), .ZN(n40) );
  INV_X1 U225 ( .A(n164), .ZN(n37) );
  XNOR2_X1 U226 ( .A(n34), .B(n5), .ZN(SUM[12]) );
  XNOR2_X1 U227 ( .A(n20), .B(n2), .ZN(SUM[15]) );
  OAI21_X1 U228 ( .B1(n171), .B2(n28), .A(n29), .ZN(n27) );
  NOR2_X1 U229 ( .A1(n32), .A2(n35), .ZN(n30) );
  OAI21_X1 U230 ( .B1(n172), .B2(n174), .A(n22), .ZN(n20) );
endmodule


module layer3_16_12_16_16_datapath_M16_N12_T16_P16_1 ( clk, clear_acc, 
        data_out_x, data_out, data_out_w, data_out_b, wr_en_y, m_valid, 
        m_ready, sel );
  input [15:0] data_out_x;
  output [15:0] data_out;
  input [15:0] data_out_w;
  input [15:0] data_out_b;
  input [4:0] sel;
  input clk, clear_acc, wr_en_y, m_valid, m_ready;
  wire   clear_acc_delay, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
         N39, N40, N41, N42, N43, N44, n1, n2, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n85, n102, n111, n112, n113, n114, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244;
  wire   [15:0] f;
  wire   [15:0] adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF_X1 clear_acc_delay_reg ( .D(n21), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \mul_out_save_reg[15]  ( .D(n226), .CK(clk), .Q(n25) );
  DFF_X1 \mul_out_save_reg[14]  ( .D(n227), .CK(clk), .Q(n26) );
  DFF_X1 \mul_out_save_reg[13]  ( .D(n228), .CK(clk), .Q(n27) );
  DFF_X1 \mul_out_save_reg[12]  ( .D(n229), .CK(clk), .Q(n28) );
  DFF_X1 \mul_out_save_reg[11]  ( .D(n230), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_save_reg[10]  ( .D(n231), .CK(clk), .Q(n32) );
  DFF_X1 \mul_out_save_reg[9]  ( .D(n232), .CK(clk), .Q(n33) );
  DFF_X1 \mul_out_save_reg[8]  ( .D(n233), .CK(clk), .Q(n34) );
  DFF_X1 \mul_out_save_reg[7]  ( .D(n234), .CK(clk), .Q(n35) );
  DFF_X1 \mul_out_save_reg[6]  ( .D(n235), .CK(clk), .Q(n36) );
  DFF_X1 \mul_out_save_reg[5]  ( .D(n236), .CK(clk), .Q(n37) );
  DFF_X1 \mul_out_save_reg[4]  ( .D(n237), .CK(clk), .Q(n38) );
  DFF_X1 \mul_out_save_reg[3]  ( .D(n238), .CK(clk), .Q(n39) );
  DFF_X1 \mul_out_save_reg[2]  ( .D(n239), .CK(clk), .Q(n40) );
  DFF_X1 \mul_out_save_reg[1]  ( .D(n240), .CK(clk), .Q(n41) );
  DFF_X1 \mul_out_save_reg[0]  ( .D(n241), .CK(clk), .Q(n43) );
  DFF_X1 \f_reg[0]  ( .D(n114), .CK(clk), .Q(f[0]), .QN(n215) );
  DFF_X1 \f_reg[1]  ( .D(n113), .CK(clk), .Q(f[1]), .QN(n216) );
  DFF_X1 \f_reg[2]  ( .D(n112), .CK(clk), .Q(f[2]), .QN(n217) );
  DFF_X1 \f_reg[8]  ( .D(n81), .CK(clk), .Q(f[8]), .QN(n219) );
  DFF_X1 \f_reg[9]  ( .D(n80), .CK(clk), .Q(f[9]), .QN(n220) );
  DFF_X1 \f_reg[10]  ( .D(n79), .CK(clk), .Q(n52), .QN(n221) );
  DFF_X1 \f_reg[11]  ( .D(n78), .CK(clk), .Q(n50), .QN(n222) );
  DFF_X1 \f_reg[12]  ( .D(n77), .CK(clk), .Q(n49), .QN(n223) );
  DFF_X1 \f_reg[14]  ( .D(n7), .CK(clk), .Q(n47), .QN(n225) );
  DFF_X1 \f_reg[15]  ( .D(n76), .CK(clk), .Q(f[15]), .QN(n73) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_1_DW_mult_tc_1 mult_2021 ( .a(
        data_out_x), .b(data_out_w), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29}) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_1_DW01_add_2 add_2022 ( .A({n205, 
        n204, n203, n202, n201, n200, n214, n213, n212, n211, n210, n209, n208, 
        n207, n206, n199}), .B({f[15], n47, n48, n49, n50, n52, f[9:0]}), .CI(
        1'b0), .SUM(adder) );
  DFF_X1 delay_reg ( .D(n166), .CK(clk), .Q(n11), .QN(n242) );
  DFF_X1 \data_out_reg[15]  ( .D(n167), .CK(clk), .Q(data_out[15]), .QN(n198)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n168), .CK(clk), .Q(data_out[14]), .QN(n197)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n169), .CK(clk), .Q(data_out[13]), .QN(n196)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n170), .CK(clk), .Q(data_out[12]), .QN(n195)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n171), .CK(clk), .Q(data_out[11]), .QN(n194)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n172), .CK(clk), .Q(data_out[10]), .QN(n193)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n173), .CK(clk), .Q(data_out[9]), .QN(n192) );
  DFF_X1 \data_out_reg[8]  ( .D(n174), .CK(clk), .Q(data_out[8]), .QN(n191) );
  DFF_X1 \data_out_reg[7]  ( .D(n175), .CK(clk), .Q(data_out[7]), .QN(n190) );
  DFF_X1 \data_out_reg[6]  ( .D(n176), .CK(clk), .Q(data_out[6]), .QN(n189) );
  DFF_X1 \data_out_reg[5]  ( .D(n177), .CK(clk), .Q(data_out[5]), .QN(n188) );
  DFF_X1 \data_out_reg[4]  ( .D(n178), .CK(clk), .Q(data_out[4]), .QN(n187) );
  DFF_X1 \data_out_reg[3]  ( .D(n179), .CK(clk), .Q(data_out[3]), .QN(n186) );
  DFF_X1 \data_out_reg[2]  ( .D(n180), .CK(clk), .Q(data_out[2]), .QN(n185) );
  DFF_X1 \data_out_reg[1]  ( .D(n181), .CK(clk), .Q(data_out[1]), .QN(n184) );
  DFF_X1 \data_out_reg[0]  ( .D(n182), .CK(clk), .Q(data_out[0]), .QN(n183) );
  DFF_X1 \f_reg[3]  ( .D(n111), .CK(clk), .Q(f[3]), .QN(n65) );
  DFF_X1 \f_reg[4]  ( .D(n102), .CK(clk), .Q(f[4]), .QN(n66) );
  DFF_X1 \f_reg[5]  ( .D(n85), .CK(clk), .Q(f[5]), .QN(n67) );
  DFF_X1 \f_reg[6]  ( .D(n83), .CK(clk), .Q(f[6]), .QN(n68) );
  DFF_X1 \f_reg[7]  ( .D(n82), .CK(clk), .Q(f[7]), .QN(n218) );
  DFF_X2 \f_reg[13]  ( .D(n1), .CK(clk), .Q(n48), .QN(n224) );
  MUX2_X2 U3 ( .A(N39), .B(n32), .S(n11), .Z(n200) );
  INV_X1 U4 ( .A(n46), .ZN(n63) );
  AND2_X1 U5 ( .A1(n46), .A2(n22), .ZN(n19) );
  AND2_X1 U6 ( .A1(n10), .A2(n8), .ZN(n2) );
  NAND3_X1 U8 ( .A1(n5), .A2(n4), .A3(n6), .ZN(n1) );
  MUX2_X2 U9 ( .A(n35), .B(N36), .S(n242), .Z(n212) );
  MUX2_X2 U10 ( .A(n34), .B(N37), .S(n242), .Z(n213) );
  MUX2_X2 U11 ( .A(n27), .B(N42), .S(n242), .Z(n203) );
  MUX2_X2 U12 ( .A(n26), .B(N43), .S(n242), .Z(n204) );
  NAND2_X1 U13 ( .A1(n9), .A2(n2), .ZN(n77) );
  NAND2_X1 U14 ( .A1(data_out_b[13]), .A2(n21), .ZN(n4) );
  NAND2_X1 U15 ( .A1(adder[13]), .A2(n19), .ZN(n5) );
  NAND2_X1 U16 ( .A1(n63), .A2(n48), .ZN(n6) );
  NAND3_X1 U17 ( .A1(n14), .A2(n13), .A3(n15), .ZN(n7) );
  MUX2_X2 U18 ( .A(n28), .B(N41), .S(n242), .Z(n202) );
  MUX2_X2 U19 ( .A(n29), .B(N40), .S(n242), .Z(n201) );
  NAND2_X1 U20 ( .A1(data_out_b[12]), .A2(n21), .ZN(n8) );
  NAND2_X1 U21 ( .A1(adder[12]), .A2(n19), .ZN(n9) );
  NAND2_X1 U22 ( .A1(n63), .A2(n49), .ZN(n10) );
  AND2_X1 U23 ( .A1(n18), .A2(n16), .ZN(n12) );
  NAND2_X1 U24 ( .A1(n17), .A2(n12), .ZN(n76) );
  NAND2_X1 U25 ( .A1(data_out_b[14]), .A2(n21), .ZN(n13) );
  NAND2_X1 U26 ( .A1(adder[14]), .A2(n19), .ZN(n14) );
  NAND2_X1 U27 ( .A1(n63), .A2(n47), .ZN(n15) );
  NAND2_X1 U28 ( .A1(data_out_b[15]), .A2(n21), .ZN(n16) );
  NAND2_X1 U29 ( .A1(adder[15]), .A2(n19), .ZN(n17) );
  NAND2_X1 U30 ( .A1(n63), .A2(f[15]), .ZN(n18) );
  NAND2_X1 U31 ( .A1(n166), .A2(n20), .ZN(n244) );
  INV_X1 U32 ( .A(clear_acc), .ZN(n22) );
  NAND3_X1 U33 ( .A1(wr_en_y), .A2(n74), .A3(n73), .ZN(n243) );
  INV_X1 U34 ( .A(n24), .ZN(n42) );
  OAI22_X1 U35 ( .A1(n186), .A2(n244), .B1(n65), .B2(n243), .ZN(n179) );
  OAI22_X1 U36 ( .A1(n187), .A2(n244), .B1(n66), .B2(n243), .ZN(n178) );
  OAI22_X1 U37 ( .A1(n188), .A2(n244), .B1(n67), .B2(n243), .ZN(n177) );
  OAI22_X1 U38 ( .A1(n189), .A2(n244), .B1(n68), .B2(n243), .ZN(n176) );
  OAI22_X1 U39 ( .A1(n190), .A2(n244), .B1(n218), .B2(n243), .ZN(n175) );
  OAI22_X1 U40 ( .A1(n191), .A2(n244), .B1(n219), .B2(n243), .ZN(n174) );
  OAI22_X1 U41 ( .A1(n192), .A2(n244), .B1(n220), .B2(n243), .ZN(n173) );
  MUX2_X1 U42 ( .A(n39), .B(N32), .S(n242), .Z(n208) );
  INV_X1 U43 ( .A(wr_en_y), .ZN(n20) );
  INV_X1 U44 ( .A(n22), .ZN(n21) );
  INV_X1 U45 ( .A(m_ready), .ZN(n23) );
  NAND2_X1 U46 ( .A1(m_valid), .A2(n23), .ZN(n44) );
  OAI21_X1 U47 ( .B1(sel[4]), .B2(n75), .A(n44), .ZN(n166) );
  NAND2_X1 U48 ( .A1(clear_acc_delay), .A2(n242), .ZN(n24) );
  MUX2_X1 U49 ( .A(n25), .B(N44), .S(n42), .Z(n226) );
  MUX2_X1 U50 ( .A(n25), .B(N44), .S(n242), .Z(n205) );
  MUX2_X1 U51 ( .A(n26), .B(N43), .S(n42), .Z(n227) );
  MUX2_X1 U52 ( .A(n27), .B(N42), .S(n42), .Z(n228) );
  MUX2_X1 U53 ( .A(n28), .B(N41), .S(n42), .Z(n229) );
  MUX2_X1 U54 ( .A(n29), .B(N40), .S(n42), .Z(n230) );
  MUX2_X1 U55 ( .A(n32), .B(N39), .S(n42), .Z(n231) );
  MUX2_X1 U56 ( .A(n33), .B(N38), .S(n42), .Z(n232) );
  MUX2_X1 U57 ( .A(n33), .B(N38), .S(n242), .Z(n214) );
  MUX2_X1 U58 ( .A(n34), .B(N37), .S(n42), .Z(n233) );
  MUX2_X1 U59 ( .A(n35), .B(N36), .S(n42), .Z(n234) );
  MUX2_X1 U60 ( .A(n36), .B(N35), .S(n42), .Z(n235) );
  MUX2_X1 U61 ( .A(n36), .B(N35), .S(n242), .Z(n211) );
  MUX2_X1 U62 ( .A(n37), .B(N34), .S(n42), .Z(n236) );
  MUX2_X1 U63 ( .A(n37), .B(N34), .S(n242), .Z(n210) );
  MUX2_X1 U64 ( .A(n38), .B(N33), .S(n42), .Z(n237) );
  MUX2_X1 U65 ( .A(n38), .B(N33), .S(n242), .Z(n209) );
  MUX2_X1 U66 ( .A(n39), .B(N32), .S(n42), .Z(n238) );
  MUX2_X1 U67 ( .A(n40), .B(N31), .S(n42), .Z(n239) );
  MUX2_X1 U68 ( .A(n40), .B(N31), .S(n242), .Z(n207) );
  MUX2_X1 U69 ( .A(n41), .B(N30), .S(n42), .Z(n240) );
  MUX2_X1 U70 ( .A(n41), .B(N30), .S(n242), .Z(n206) );
  MUX2_X1 U71 ( .A(n43), .B(N29), .S(n42), .Z(n241) );
  MUX2_X1 U72 ( .A(n43), .B(N29), .S(n242), .Z(n199) );
  INV_X1 U73 ( .A(n44), .ZN(n45) );
  OAI21_X1 U74 ( .B1(n45), .B2(n11), .A(n22), .ZN(n46) );
  AOI222_X1 U75 ( .A1(data_out_b[11]), .A2(n21), .B1(adder[11]), .B2(n19), 
        .C1(n63), .C2(n50), .ZN(n51) );
  INV_X1 U76 ( .A(n51), .ZN(n78) );
  AOI222_X1 U77 ( .A1(data_out_b[10]), .A2(n21), .B1(adder[10]), .B2(n19), 
        .C1(n63), .C2(n52), .ZN(n53) );
  INV_X1 U78 ( .A(n53), .ZN(n79) );
  AOI222_X1 U79 ( .A1(data_out_b[8]), .A2(n21), .B1(adder[8]), .B2(n19), .C1(
        n63), .C2(f[8]), .ZN(n54) );
  INV_X1 U80 ( .A(n54), .ZN(n81) );
  AOI222_X1 U81 ( .A1(data_out_b[7]), .A2(n21), .B1(adder[7]), .B2(n19), .C1(
        n63), .C2(f[7]), .ZN(n55) );
  INV_X1 U82 ( .A(n55), .ZN(n82) );
  AOI222_X1 U83 ( .A1(data_out_b[6]), .A2(n21), .B1(adder[6]), .B2(n19), .C1(
        n63), .C2(f[6]), .ZN(n56) );
  INV_X1 U84 ( .A(n56), .ZN(n83) );
  AOI222_X1 U85 ( .A1(data_out_b[5]), .A2(n21), .B1(adder[5]), .B2(n19), .C1(
        n63), .C2(f[5]), .ZN(n57) );
  INV_X1 U86 ( .A(n57), .ZN(n85) );
  AOI222_X1 U87 ( .A1(data_out_b[4]), .A2(n21), .B1(adder[4]), .B2(n19), .C1(
        n63), .C2(f[4]), .ZN(n58) );
  INV_X1 U88 ( .A(n58), .ZN(n102) );
  AOI222_X1 U89 ( .A1(data_out_b[3]), .A2(n21), .B1(adder[3]), .B2(n19), .C1(
        n63), .C2(f[3]), .ZN(n59) );
  INV_X1 U90 ( .A(n59), .ZN(n111) );
  AOI222_X1 U91 ( .A1(data_out_b[2]), .A2(n21), .B1(adder[2]), .B2(n19), .C1(
        n63), .C2(f[2]), .ZN(n60) );
  INV_X1 U92 ( .A(n60), .ZN(n112) );
  AOI222_X1 U93 ( .A1(data_out_b[1]), .A2(n21), .B1(adder[1]), .B2(n19), .C1(
        n63), .C2(f[1]), .ZN(n61) );
  INV_X1 U94 ( .A(n61), .ZN(n113) );
  AOI222_X1 U95 ( .A1(data_out_b[0]), .A2(n21), .B1(adder[0]), .B2(n19), .C1(
        n63), .C2(f[0]), .ZN(n62) );
  INV_X1 U96 ( .A(n62), .ZN(n114) );
  AOI222_X1 U97 ( .A1(data_out_b[9]), .A2(n21), .B1(adder[9]), .B2(n19), .C1(
        n63), .C2(f[9]), .ZN(n64) );
  INV_X1 U98 ( .A(n64), .ZN(n80) );
  NOR4_X1 U99 ( .A1(n50), .A2(n49), .A3(n48), .A4(n47), .ZN(n72) );
  NOR4_X1 U100 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(n52), .ZN(n71) );
  NAND4_X1 U101 ( .A1(n68), .A2(n67), .A3(n66), .A4(n65), .ZN(n69) );
  NOR4_X1 U102 ( .A1(n69), .A2(f[0]), .A3(f[1]), .A4(f[2]), .ZN(n70) );
  NAND3_X1 U103 ( .A1(n72), .A2(n71), .A3(n70), .ZN(n74) );
  OAI22_X1 U104 ( .A1(n183), .A2(n244), .B1(n215), .B2(n243), .ZN(n182) );
  OAI22_X1 U105 ( .A1(n184), .A2(n244), .B1(n216), .B2(n243), .ZN(n181) );
  OAI22_X1 U106 ( .A1(n185), .A2(n244), .B1(n217), .B2(n243), .ZN(n180) );
  OAI22_X1 U107 ( .A1(n193), .A2(n244), .B1(n221), .B2(n243), .ZN(n172) );
  OAI22_X1 U108 ( .A1(n194), .A2(n244), .B1(n222), .B2(n243), .ZN(n171) );
  OAI22_X1 U109 ( .A1(n195), .A2(n244), .B1(n223), .B2(n243), .ZN(n170) );
  OAI22_X1 U110 ( .A1(n196), .A2(n244), .B1(n224), .B2(n243), .ZN(n169) );
  OAI22_X1 U111 ( .A1(n197), .A2(n244), .B1(n225), .B2(n243), .ZN(n168) );
  OAI22_X1 U112 ( .A1(n198), .A2(n244), .B1(n73), .B2(n243), .ZN(n167) );
  AND4_X1 U113 ( .A1(sel[3]), .A2(sel[2]), .A3(sel[1]), .A4(sel[0]), .ZN(n75)
         );
endmodule


module layer3_16_12_16_16_ctrlpath_M16_N12_T16_P16 ( clk, reset, s_valid, 
        s_ready, m_valid, m_ready, clear_acc, wr_en_x, wr_en_y, sel, addr_x, 
        addr_w_0, addr_b_0, addr_w_1, addr_b_1, addr_w_2, addr_b_2, addr_w_3, 
        addr_b_3, addr_w_4, addr_b_4, addr_w_5, addr_b_5, addr_w_6, addr_b_6, 
        addr_w_7, addr_b_7, addr_w_8, addr_b_8, addr_w_9, addr_b_9, addr_w_10, 
        addr_b_10, addr_w_11, addr_b_11, addr_w_12, addr_b_12, addr_w_13, 
        addr_b_13, addr_w_14, addr_b_14, addr_w_15, addr_b_15 );
  output [4:0] sel;
  output [3:0] addr_x;
  output [3:0] addr_w_0;
  output [0:0] addr_b_0;
  output [3:0] addr_w_1;
  output [0:0] addr_b_1;
  output [3:0] addr_w_2;
  output [0:0] addr_b_2;
  output [3:0] addr_w_3;
  output [0:0] addr_b_3;
  output [3:0] addr_w_4;
  output [0:0] addr_b_4;
  output [3:0] addr_w_5;
  output [0:0] addr_b_5;
  output [3:0] addr_w_6;
  output [0:0] addr_b_6;
  output [3:0] addr_w_7;
  output [0:0] addr_b_7;
  output [3:0] addr_w_8;
  output [0:0] addr_b_8;
  output [3:0] addr_w_9;
  output [0:0] addr_b_9;
  output [3:0] addr_w_10;
  output [0:0] addr_b_10;
  output [3:0] addr_w_11;
  output [0:0] addr_b_11;
  output [3:0] addr_w_12;
  output [0:0] addr_b_12;
  output [3:0] addr_w_13;
  output [0:0] addr_b_13;
  output [3:0] addr_w_14;
  output [0:0] addr_b_14;
  output [3:0] addr_w_15;
  output [0:0] addr_b_15;
  input clk, reset, s_valid, m_ready;
  output s_ready, m_valid, clear_acc, wr_en_x, wr_en_y;
  wire   n132, N11, clear_acc_delay, N221, N222, N223, N224, N243, N244, N245,
         N246, N265, N266, N267, N268, N287, N288, N289, N290, N309, N310,
         N311, N312, N331, N332, N333, N334, N353, N354, N355, N356, N375,
         N376, N377, N378, N397, N398, N399, N400, N419, N420, N421, N422,
         N441, N442, N443, N444, N463, N464, N465, N466, N485, N486, N487,
         N488, N507, N508, N509, N510, N529, N530, N531, N532, N551, N552,
         N553, N554, N569, n55, n151, n152, n153, n155, n156, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n183, n184, n185, n186, n191, n193,
         n194, n195, n196, n197, n198, n200, n201, n202, n203, n205, n206,
         n207, n208, n210, n211, n212, n213, n215, n216, n217, n218, n220,
         n221, n222, n223, n225, n226, n227, n228, n230, n231, n232, n233,
         n235, n236, n237, n238, n240, n241, n242, n243, n245, n246, n247,
         n248, n250, n251, n252, n253, n255, n256, n257, n258, n260, n261,
         n262, n263, n265, n266, n267, n268, n270, n271, n272, n273, n278,
         n279, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n295, n296, n306, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, \r444/GE_LT_GT_LE ,
         \add_2461_S2/carry[3] , \add_2461_S2/carry[2] ,
         \add_2453_S2/carry[3] , \add_2453_S2/carry[2] ,
         \add_2445_S2/carry[3] , \add_2445_S2/carry[2] ,
         \add_2437_S2/carry[3] , \add_2437_S2/carry[2] ,
         \add_2429_S2/carry[3] , \add_2429_S2/carry[2] ,
         \add_2421_S2/carry[3] , \add_2421_S2/carry[2] ,
         \add_2413_S2/carry[3] , \add_2413_S2/carry[2] ,
         \add_2405_S2/carry[3] , \add_2405_S2/carry[2] ,
         \add_2397_S2/carry[3] , \add_2397_S2/carry[2] ,
         \add_2389_S2/carry[3] , \add_2389_S2/carry[2] ,
         \add_2381_S2/carry[3] , \add_2381_S2/carry[2] ,
         \add_2373_S2/carry[3] , \add_2373_S2/carry[2] ,
         \add_2365_S2/carry[3] , \add_2365_S2/carry[2] ,
         \add_2357_S2/carry[3] , \add_2357_S2/carry[2] ,
         \add_2349_S2/carry[3] , \add_2349_S2/carry[2] ,
         \add_2341_S2/carry[3] , \add_2341_S2/carry[2] , n1, n2, n4, n5, n7,
         n8, n9, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131;
  wire   [3:0] state;

  DFF_X1 \state_reg[0]  ( .D(N11), .CK(clk), .Q(state[0]), .QN(n153) );
  DFF_X1 wr_en_y_reg ( .D(n131), .CK(clk), .Q(wr_en_y) );
  DFF_X1 \sel_count_reg[4]  ( .D(n342), .CK(clk), .Q(sel[4]), .QN(n177) );
  DFF_X1 \sel_count_reg[2]  ( .D(n340), .CK(clk), .Q(sel[2]), .QN(n184) );
  DFF_X1 \sel_count_reg[3]  ( .D(n339), .CK(clk), .Q(sel[3]), .QN(n183) );
  DFF_X1 \state_reg[1]  ( .D(n60), .CK(clk), .Q(state[1]), .QN(n152) );
  DFF_X1 \addr_x_reg[2]  ( .D(n336), .CK(clk), .Q(addr_x[2]), .QN(n156) );
  DFF_X1 \addr_x_reg[3]  ( .D(n338), .CK(clk), .Q(addr_x[3]), .QN(n155) );
  DFF_X1 \addr_w2_15_reg[0]  ( .D(n126), .CK(clk), .Q(addr_w_15[0]), .QN(N551)
         );
  DFF_X1 \addr_w2_15_reg[1]  ( .D(n127), .CK(clk), .Q(addr_w_15[1]) );
  DFF_X1 \addr_w2_15_reg[2]  ( .D(n128), .CK(clk), .Q(addr_w_15[2]) );
  DFF_X1 \addr_w2_15_reg[3]  ( .D(n129), .CK(clk), .Q(addr_w_15[3]) );
  DFF_X1 \addr_w2_14_reg[0]  ( .D(n122), .CK(clk), .Q(addr_w_14[0]), .QN(N529)
         );
  DFF_X1 \addr_w2_14_reg[1]  ( .D(n123), .CK(clk), .Q(addr_w_14[1]) );
  DFF_X1 \addr_w2_14_reg[2]  ( .D(n124), .CK(clk), .Q(addr_w_14[2]) );
  DFF_X1 \addr_w2_14_reg[3]  ( .D(n125), .CK(clk), .Q(addr_w_14[3]) );
  DFF_X1 \addr_w2_13_reg[0]  ( .D(n118), .CK(clk), .Q(addr_w_13[0]), .QN(N507)
         );
  DFF_X1 \addr_w2_13_reg[1]  ( .D(n119), .CK(clk), .Q(addr_w_13[1]) );
  DFF_X1 \addr_w2_13_reg[2]  ( .D(n120), .CK(clk), .Q(addr_w_13[2]) );
  DFF_X1 \addr_w2_13_reg[3]  ( .D(n121), .CK(clk), .Q(addr_w_13[3]) );
  DFF_X1 \addr_w2_12_reg[0]  ( .D(n114), .CK(clk), .Q(addr_w_12[0]), .QN(N485)
         );
  DFF_X1 \addr_w2_12_reg[1]  ( .D(n115), .CK(clk), .Q(addr_w_12[1]) );
  DFF_X1 \addr_w2_12_reg[2]  ( .D(n116), .CK(clk), .Q(addr_w_12[2]) );
  DFF_X1 \addr_w2_12_reg[3]  ( .D(n117), .CK(clk), .Q(addr_w_12[3]) );
  DFF_X1 \addr_w2_11_reg[0]  ( .D(n110), .CK(clk), .Q(addr_w_11[0]), .QN(N463)
         );
  DFF_X1 \addr_w2_11_reg[1]  ( .D(n111), .CK(clk), .Q(addr_w_11[1]) );
  DFF_X1 \addr_w2_11_reg[2]  ( .D(n112), .CK(clk), .Q(addr_w_11[2]) );
  DFF_X1 \addr_w2_11_reg[3]  ( .D(n113), .CK(clk), .Q(addr_w_11[3]) );
  DFF_X1 \addr_w2_10_reg[0]  ( .D(n106), .CK(clk), .Q(addr_w_10[0]), .QN(N441)
         );
  DFF_X1 \addr_w2_10_reg[1]  ( .D(n107), .CK(clk), .Q(addr_w_10[1]) );
  DFF_X1 \addr_w2_10_reg[2]  ( .D(n108), .CK(clk), .Q(addr_w_10[2]) );
  DFF_X1 \addr_w2_10_reg[3]  ( .D(n109), .CK(clk), .Q(addr_w_10[3]) );
  DFF_X1 \addr_w2_9_reg[0]  ( .D(n102), .CK(clk), .Q(addr_w_9[0]), .QN(N419)
         );
  DFF_X1 \addr_w2_9_reg[1]  ( .D(n103), .CK(clk), .Q(addr_w_9[1]) );
  DFF_X1 \addr_w2_9_reg[2]  ( .D(n104), .CK(clk), .Q(addr_w_9[2]) );
  DFF_X1 \addr_w2_9_reg[3]  ( .D(n105), .CK(clk), .Q(addr_w_9[3]) );
  DFF_X1 \addr_w2_8_reg[0]  ( .D(n98), .CK(clk), .Q(addr_w_8[0]), .QN(N397) );
  DFF_X1 \addr_w2_8_reg[1]  ( .D(n99), .CK(clk), .Q(addr_w_8[1]) );
  DFF_X1 \addr_w2_8_reg[2]  ( .D(n100), .CK(clk), .Q(addr_w_8[2]) );
  DFF_X1 \addr_w2_8_reg[3]  ( .D(n101), .CK(clk), .Q(addr_w_8[3]) );
  DFF_X1 \addr_w2_7_reg[0]  ( .D(n94), .CK(clk), .Q(addr_w_7[0]), .QN(N375) );
  DFF_X1 \addr_w2_7_reg[1]  ( .D(n95), .CK(clk), .Q(addr_w_7[1]) );
  DFF_X1 \addr_w2_7_reg[2]  ( .D(n96), .CK(clk), .Q(addr_w_7[2]) );
  DFF_X1 \addr_w2_7_reg[3]  ( .D(n97), .CK(clk), .Q(addr_w_7[3]) );
  DFF_X1 \addr_w2_6_reg[0]  ( .D(n90), .CK(clk), .Q(addr_w_6[0]), .QN(N353) );
  DFF_X1 \addr_w2_6_reg[1]  ( .D(n91), .CK(clk), .Q(addr_w_6[1]) );
  DFF_X1 \addr_w2_6_reg[2]  ( .D(n92), .CK(clk), .Q(addr_w_6[2]) );
  DFF_X1 \addr_w2_6_reg[3]  ( .D(n93), .CK(clk), .Q(addr_w_6[3]) );
  DFF_X1 \addr_w2_5_reg[0]  ( .D(n86), .CK(clk), .Q(addr_w_5[0]), .QN(N331) );
  DFF_X1 \addr_w2_5_reg[1]  ( .D(n87), .CK(clk), .Q(addr_w_5[1]) );
  DFF_X1 \addr_w2_5_reg[2]  ( .D(n88), .CK(clk), .Q(addr_w_5[2]) );
  DFF_X1 \addr_w2_5_reg[3]  ( .D(n89), .CK(clk), .Q(addr_w_5[3]) );
  DFF_X1 \addr_w2_4_reg[0]  ( .D(n82), .CK(clk), .Q(addr_w_4[0]), .QN(N309) );
  DFF_X1 \addr_w2_4_reg[1]  ( .D(n83), .CK(clk), .Q(addr_w_4[1]) );
  DFF_X1 \addr_w2_4_reg[2]  ( .D(n84), .CK(clk), .Q(addr_w_4[2]) );
  DFF_X1 \addr_w2_4_reg[3]  ( .D(n85), .CK(clk), .Q(addr_w_4[3]) );
  DFF_X1 \addr_w2_3_reg[0]  ( .D(n78), .CK(clk), .Q(addr_w_3[0]), .QN(N287) );
  DFF_X1 \addr_w2_3_reg[1]  ( .D(n79), .CK(clk), .Q(addr_w_3[1]) );
  DFF_X1 \addr_w2_3_reg[2]  ( .D(n80), .CK(clk), .Q(addr_w_3[2]) );
  DFF_X1 \addr_w2_3_reg[3]  ( .D(n81), .CK(clk), .Q(addr_w_3[3]) );
  DFF_X1 \addr_w2_2_reg[0]  ( .D(n74), .CK(clk), .Q(addr_w_2[0]), .QN(N265) );
  DFF_X1 \addr_w2_2_reg[1]  ( .D(n75), .CK(clk), .Q(addr_w_2[1]) );
  DFF_X1 \addr_w2_2_reg[2]  ( .D(n76), .CK(clk), .Q(addr_w_2[2]) );
  DFF_X1 \addr_w2_2_reg[3]  ( .D(n77), .CK(clk), .Q(addr_w_2[3]) );
  DFF_X1 \addr_w2_1_reg[0]  ( .D(n70), .CK(clk), .Q(addr_w_1[0]), .QN(N243) );
  DFF_X1 \addr_w2_1_reg[1]  ( .D(n71), .CK(clk), .Q(addr_w_1[1]) );
  DFF_X1 \addr_w2_1_reg[2]  ( .D(n72), .CK(clk), .Q(addr_w_1[2]) );
  DFF_X1 \addr_w2_1_reg[3]  ( .D(n73), .CK(clk), .Q(addr_w_1[3]) );
  DFF_X1 \addr_w2_0_reg[0]  ( .D(n66), .CK(clk), .Q(addr_w_0[0]), .QN(N221) );
  DFF_X1 \addr_w2_0_reg[1]  ( .D(n67), .CK(clk), .Q(addr_w_0[1]) );
  DFF_X1 \addr_w2_0_reg[2]  ( .D(n68), .CK(clk), .Q(addr_w_0[2]) );
  DFF_X1 \addr_w2_0_reg[3]  ( .D(n69), .CK(clk), .Q(addr_w_0[3]) );
  NAND3_X1 U267 ( .A1(addr_x[1]), .A2(n156), .A3(n283), .ZN(n282) );
  NAND3_X1 U268 ( .A1(n295), .A2(n62), .A3(wr_en_y), .ZN(n296) );
  HA_X1 \add_2461_S2/U1_1_1  ( .A(addr_w_15[1]), .B(addr_w_15[0]), .CO(
        \add_2461_S2/carry[2] ), .S(N552) );
  HA_X1 \add_2461_S2/U1_1_2  ( .A(addr_w_15[2]), .B(\add_2461_S2/carry[2] ), 
        .CO(\add_2461_S2/carry[3] ), .S(N553) );
  HA_X1 \add_2453_S2/U1_1_1  ( .A(addr_w_14[1]), .B(addr_w_14[0]), .CO(
        \add_2453_S2/carry[2] ), .S(N530) );
  HA_X1 \add_2453_S2/U1_1_2  ( .A(addr_w_14[2]), .B(\add_2453_S2/carry[2] ), 
        .CO(\add_2453_S2/carry[3] ), .S(N531) );
  HA_X1 \add_2445_S2/U1_1_1  ( .A(addr_w_13[1]), .B(addr_w_13[0]), .CO(
        \add_2445_S2/carry[2] ), .S(N508) );
  HA_X1 \add_2445_S2/U1_1_2  ( .A(addr_w_13[2]), .B(\add_2445_S2/carry[2] ), 
        .CO(\add_2445_S2/carry[3] ), .S(N509) );
  HA_X1 \add_2437_S2/U1_1_1  ( .A(addr_w_12[1]), .B(addr_w_12[0]), .CO(
        \add_2437_S2/carry[2] ), .S(N486) );
  HA_X1 \add_2437_S2/U1_1_2  ( .A(addr_w_12[2]), .B(\add_2437_S2/carry[2] ), 
        .CO(\add_2437_S2/carry[3] ), .S(N487) );
  HA_X1 \add_2429_S2/U1_1_1  ( .A(addr_w_11[1]), .B(addr_w_11[0]), .CO(
        \add_2429_S2/carry[2] ), .S(N464) );
  HA_X1 \add_2429_S2/U1_1_2  ( .A(addr_w_11[2]), .B(\add_2429_S2/carry[2] ), 
        .CO(\add_2429_S2/carry[3] ), .S(N465) );
  HA_X1 \add_2421_S2/U1_1_1  ( .A(addr_w_10[1]), .B(addr_w_10[0]), .CO(
        \add_2421_S2/carry[2] ), .S(N442) );
  HA_X1 \add_2421_S2/U1_1_2  ( .A(addr_w_10[2]), .B(\add_2421_S2/carry[2] ), 
        .CO(\add_2421_S2/carry[3] ), .S(N443) );
  HA_X1 \add_2413_S2/U1_1_1  ( .A(addr_w_9[1]), .B(addr_w_9[0]), .CO(
        \add_2413_S2/carry[2] ), .S(N420) );
  HA_X1 \add_2413_S2/U1_1_2  ( .A(addr_w_9[2]), .B(\add_2413_S2/carry[2] ), 
        .CO(\add_2413_S2/carry[3] ), .S(N421) );
  HA_X1 \add_2405_S2/U1_1_1  ( .A(addr_w_8[1]), .B(addr_w_8[0]), .CO(
        \add_2405_S2/carry[2] ), .S(N398) );
  HA_X1 \add_2405_S2/U1_1_2  ( .A(addr_w_8[2]), .B(\add_2405_S2/carry[2] ), 
        .CO(\add_2405_S2/carry[3] ), .S(N399) );
  HA_X1 \add_2397_S2/U1_1_1  ( .A(addr_w_7[1]), .B(addr_w_7[0]), .CO(
        \add_2397_S2/carry[2] ), .S(N376) );
  HA_X1 \add_2397_S2/U1_1_2  ( .A(addr_w_7[2]), .B(\add_2397_S2/carry[2] ), 
        .CO(\add_2397_S2/carry[3] ), .S(N377) );
  HA_X1 \add_2389_S2/U1_1_1  ( .A(addr_w_6[1]), .B(addr_w_6[0]), .CO(
        \add_2389_S2/carry[2] ), .S(N354) );
  HA_X1 \add_2389_S2/U1_1_2  ( .A(addr_w_6[2]), .B(\add_2389_S2/carry[2] ), 
        .CO(\add_2389_S2/carry[3] ), .S(N355) );
  HA_X1 \add_2381_S2/U1_1_1  ( .A(addr_w_5[1]), .B(addr_w_5[0]), .CO(
        \add_2381_S2/carry[2] ), .S(N332) );
  HA_X1 \add_2381_S2/U1_1_2  ( .A(addr_w_5[2]), .B(\add_2381_S2/carry[2] ), 
        .CO(\add_2381_S2/carry[3] ), .S(N333) );
  HA_X1 \add_2373_S2/U1_1_1  ( .A(addr_w_4[1]), .B(addr_w_4[0]), .CO(
        \add_2373_S2/carry[2] ), .S(N310) );
  HA_X1 \add_2373_S2/U1_1_2  ( .A(addr_w_4[2]), .B(\add_2373_S2/carry[2] ), 
        .CO(\add_2373_S2/carry[3] ), .S(N311) );
  HA_X1 \add_2365_S2/U1_1_1  ( .A(addr_w_3[1]), .B(addr_w_3[0]), .CO(
        \add_2365_S2/carry[2] ), .S(N288) );
  HA_X1 \add_2365_S2/U1_1_2  ( .A(addr_w_3[2]), .B(\add_2365_S2/carry[2] ), 
        .CO(\add_2365_S2/carry[3] ), .S(N289) );
  HA_X1 \add_2357_S2/U1_1_1  ( .A(addr_w_2[1]), .B(addr_w_2[0]), .CO(
        \add_2357_S2/carry[2] ), .S(N266) );
  HA_X1 \add_2357_S2/U1_1_2  ( .A(addr_w_2[2]), .B(\add_2357_S2/carry[2] ), 
        .CO(\add_2357_S2/carry[3] ), .S(N267) );
  HA_X1 \add_2349_S2/U1_1_1  ( .A(addr_w_1[1]), .B(addr_w_1[0]), .CO(
        \add_2349_S2/carry[2] ), .S(N244) );
  HA_X1 \add_2349_S2/U1_1_2  ( .A(addr_w_1[2]), .B(\add_2349_S2/carry[2] ), 
        .CO(\add_2349_S2/carry[3] ), .S(N245) );
  HA_X1 \add_2341_S2/U1_1_1  ( .A(addr_w_0[1]), .B(addr_w_0[0]), .CO(
        \add_2341_S2/carry[2] ), .S(N222) );
  HA_X1 \add_2341_S2/U1_1_2  ( .A(addr_w_0[2]), .B(\add_2341_S2/carry[2] ), 
        .CO(\add_2341_S2/carry[3] ), .S(N223) );
  DFF_X1 \sel_count_reg[0]  ( .D(n344), .CK(clk), .Q(sel[0]), .QN(n186) );
  DFF_X1 \sel_count_reg[1]  ( .D(n341), .CK(clk), .Q(n132), .QN(n185) );
  DFF_X1 clear_acc_delay_reg ( .D(n5), .CK(clk), .Q(clear_acc_delay), .QN(n175) );
  DFF_X1 clear_acc_reg ( .D(N569), .CK(clk), .Q(clear_acc), .QN(n55) );
  DFF_X1 \addr_b_15_reg[0]  ( .D(n331), .CK(clk), .Q(addr_b_15[0]), .QN(n174)
         );
  DFF_X1 \addr_b_14_reg[0]  ( .D(n330), .CK(clk), .Q(addr_b_14[0]), .QN(n173)
         );
  DFF_X1 \addr_b_13_reg[0]  ( .D(n329), .CK(clk), .Q(addr_b_13[0]), .QN(n172)
         );
  DFF_X1 \addr_b_12_reg[0]  ( .D(n328), .CK(clk), .Q(addr_b_12[0]), .QN(n171)
         );
  DFF_X1 \addr_b_11_reg[0]  ( .D(n327), .CK(clk), .Q(addr_b_11[0]), .QN(n170)
         );
  DFF_X1 \addr_b_10_reg[0]  ( .D(n326), .CK(clk), .Q(addr_b_10[0]), .QN(n169)
         );
  DFF_X1 \addr_b_9_reg[0]  ( .D(n325), .CK(clk), .Q(addr_b_9[0]), .QN(n168) );
  DFF_X1 \addr_b_8_reg[0]  ( .D(n324), .CK(clk), .Q(addr_b_8[0]), .QN(n167) );
  DFF_X1 \addr_b_7_reg[0]  ( .D(n323), .CK(clk), .Q(addr_b_7[0]), .QN(n166) );
  DFF_X1 \addr_b_6_reg[0]  ( .D(n322), .CK(clk), .Q(addr_b_6[0]), .QN(n165) );
  DFF_X1 \addr_b_5_reg[0]  ( .D(n321), .CK(clk), .Q(addr_b_5[0]), .QN(n164) );
  DFF_X1 \addr_b_4_reg[0]  ( .D(n320), .CK(clk), .Q(addr_b_4[0]), .QN(n163) );
  DFF_X1 \addr_b_3_reg[0]  ( .D(n335), .CK(clk), .Q(addr_b_3[0]), .QN(n162) );
  DFF_X1 \addr_b_2_reg[0]  ( .D(n334), .CK(clk), .Q(addr_b_2[0]), .QN(n161) );
  DFF_X1 \addr_b_1_reg[0]  ( .D(n333), .CK(clk), .Q(addr_b_1[0]), .QN(n160) );
  DFF_X1 \addr_b_0_reg[0]  ( .D(n332), .CK(clk), .Q(addr_b_0[0]), .QN(n159) );
  DFF_X1 \addr_x_reg[0]  ( .D(n337), .CK(clk), .Q(addr_x[0]), .QN(n29) );
  DFF_X1 \addr_x_reg[1]  ( .D(n65), .CK(clk), .Q(addr_x[1]), .QN(n28) );
  DFF_X1 m_valid_reg ( .D(n343), .CK(clk), .Q(m_valid), .QN(n176) );
  SDFF_X1 \state_reg[2]  ( .D(1'b0), .SI(n191), .SE(n62), .CK(clk), .Q(
        state[2]), .QN(n151) );
  NOR4_X1 U3 ( .A1(n61), .A2(n7), .A3(n194), .A4(reset), .ZN(n195) );
  CLKBUF_X1 U4 ( .A(n56), .Z(n1) );
  NAND2_X1 U5 ( .A1(n132), .A2(n2), .ZN(n48) );
  NOR2_X1 U6 ( .A1(n186), .A2(n184), .ZN(n2) );
  NOR2_X1 U8 ( .A1(n55), .A2(n4), .ZN(n5) );
  INV_X1 U9 ( .A(n11), .ZN(n4) );
  INV_X1 U10 ( .A(n185), .ZN(sel[1]) );
  OAI22_X1 U11 ( .A1(n56), .A2(n191), .B1(reset), .B2(n54), .ZN(s_ready) );
  BUF_X1 U12 ( .A(n194), .Z(n17) );
  BUF_X1 U13 ( .A(n194), .Z(n18) );
  NAND4_X1 U14 ( .A1(n290), .A2(n130), .A3(n287), .A4(n62), .ZN(n286) );
  BUF_X1 U15 ( .A(n195), .Z(n14) );
  BUF_X1 U16 ( .A(n195), .Z(n15) );
  BUF_X1 U17 ( .A(n195), .Z(n16) );
  AND2_X1 U18 ( .A1(n8), .A2(n62), .ZN(n194) );
  AND2_X1 U19 ( .A1(n12), .A2(n42), .ZN(n7) );
  OAI21_X1 U20 ( .B1(n47), .B2(n131), .A(n62), .ZN(n56) );
  NOR2_X1 U21 ( .A1(n306), .A2(n7), .ZN(n290) );
  AND3_X1 U22 ( .A1(n11), .A2(n59), .A3(n58), .ZN(n8) );
  AND2_X1 U23 ( .A1(n36), .A2(n62), .ZN(n9) );
  NAND2_X1 U24 ( .A1(n290), .A2(n62), .ZN(N569) );
  OAI211_X2 U25 ( .C1(n153), .C2(n152), .A(n175), .B(n62), .ZN(n278) );
  NAND2_X1 U26 ( .A1(clear_acc_delay), .A2(n62), .ZN(n279) );
  AND3_X1 U27 ( .A1(s_valid), .A2(n53), .A3(n52), .ZN(wr_en_x) );
  NOR2_X1 U28 ( .A1(n287), .A2(n29), .ZN(n283) );
  OAI21_X1 U29 ( .B1(addr_x[0]), .B2(n287), .A(n286), .ZN(n285) );
  OAI22_X1 U30 ( .A1(n278), .A2(n162), .B1(addr_b_3[0]), .B2(n279), .ZN(n335)
         );
  OAI22_X1 U31 ( .A1(n278), .A2(n161), .B1(addr_b_2[0]), .B2(n279), .ZN(n334)
         );
  OAI22_X1 U32 ( .A1(n278), .A2(n160), .B1(addr_b_1[0]), .B2(n279), .ZN(n333)
         );
  OAI22_X1 U33 ( .A1(n278), .A2(n159), .B1(addr_b_0[0]), .B2(n279), .ZN(n332)
         );
  OAI22_X1 U34 ( .A1(n278), .A2(n174), .B1(addr_b_15[0]), .B2(n279), .ZN(n331)
         );
  OAI22_X1 U35 ( .A1(n278), .A2(n173), .B1(addr_b_14[0]), .B2(n279), .ZN(n330)
         );
  OAI22_X1 U36 ( .A1(n278), .A2(n172), .B1(addr_b_13[0]), .B2(n279), .ZN(n329)
         );
  OAI22_X1 U37 ( .A1(n278), .A2(n171), .B1(addr_b_12[0]), .B2(n279), .ZN(n328)
         );
  OAI22_X1 U38 ( .A1(n278), .A2(n170), .B1(addr_b_11[0]), .B2(n279), .ZN(n327)
         );
  OAI22_X1 U39 ( .A1(n278), .A2(n169), .B1(addr_b_10[0]), .B2(n279), .ZN(n326)
         );
  OAI22_X1 U40 ( .A1(n278), .A2(n168), .B1(addr_b_9[0]), .B2(n279), .ZN(n325)
         );
  OAI22_X1 U41 ( .A1(n278), .A2(n167), .B1(addr_b_8[0]), .B2(n279), .ZN(n324)
         );
  OAI22_X1 U42 ( .A1(n278), .A2(n166), .B1(addr_b_7[0]), .B2(n279), .ZN(n323)
         );
  OAI22_X1 U43 ( .A1(n278), .A2(n165), .B1(addr_b_6[0]), .B2(n279), .ZN(n322)
         );
  OAI22_X1 U44 ( .A1(n278), .A2(n164), .B1(addr_b_5[0]), .B2(n279), .ZN(n321)
         );
  OAI22_X1 U45 ( .A1(n278), .A2(n163), .B1(addr_b_4[0]), .B2(n279), .ZN(n320)
         );
  OR2_X1 U46 ( .A1(n183), .A2(n48), .ZN(n40) );
  XOR2_X1 U47 ( .A(sel[0]), .B(n185), .Z(n37) );
  AOI21_X1 U48 ( .B1(n28), .B2(n64), .A(n285), .ZN(n281) );
  OAI22_X1 U49 ( .A1(n29), .A2(n286), .B1(addr_x[0]), .B2(n287), .ZN(n337) );
  OAI21_X1 U50 ( .B1(\r444/GE_LT_GT_LE ), .B2(n291), .A(n62), .ZN(n295) );
  NOR2_X1 U51 ( .A1(n176), .A2(m_ready), .ZN(n291) );
  AND3_X1 U52 ( .A1(n153), .A2(state[2]), .A3(n152), .ZN(n11) );
  AND3_X1 U53 ( .A1(n151), .A2(state[0]), .A3(state[1]), .ZN(n12) );
  AND2_X1 U54 ( .A1(state[1]), .A2(state[2]), .ZN(n13) );
  NAND4_X1 U55 ( .A1(n283), .A2(addr_x[1]), .A3(addr_x[2]), .A4(n155), .ZN(
        n288) );
  OAI21_X1 U56 ( .B1(n287), .B2(addr_x[2]), .A(n281), .ZN(n289) );
  INV_X1 U57 ( .A(n251), .ZN(n84) );
  AOI22_X1 U58 ( .A1(N311), .A2(n17), .B1(addr_w_4[2]), .B2(n15), .ZN(n251) );
  INV_X1 U59 ( .A(n256), .ZN(n80) );
  AOI22_X1 U60 ( .A1(N289), .A2(n17), .B1(addr_w_3[2]), .B2(n15), .ZN(n256) );
  INV_X1 U61 ( .A(n250), .ZN(n85) );
  AOI22_X1 U62 ( .A1(N312), .A2(n17), .B1(addr_w_4[3]), .B2(n15), .ZN(n250) );
  XOR2_X1 U63 ( .A(addr_w_4[3]), .B(\add_2373_S2/carry[3] ), .Z(N312) );
  INV_X1 U64 ( .A(n253), .ZN(n82) );
  AOI22_X1 U65 ( .A1(N309), .A2(n17), .B1(addr_w_4[0]), .B2(n15), .ZN(n253) );
  INV_X1 U66 ( .A(n218), .ZN(n110) );
  AOI22_X1 U67 ( .A1(N463), .A2(n17), .B1(addr_w_11[0]), .B2(n16), .ZN(n218)
         );
  INV_X1 U68 ( .A(n223), .ZN(n106) );
  AOI22_X1 U69 ( .A1(N441), .A2(n17), .B1(addr_w_10[0]), .B2(n14), .ZN(n223)
         );
  INV_X1 U70 ( .A(n213), .ZN(n114) );
  AOI22_X1 U71 ( .A1(N485), .A2(n17), .B1(addr_w_12[0]), .B2(n15), .ZN(n213)
         );
  INV_X1 U72 ( .A(n273), .ZN(n66) );
  AOI22_X1 U73 ( .A1(N221), .A2(n194), .B1(addr_w_0[0]), .B2(n14), .ZN(n273)
         );
  INV_X1 U74 ( .A(n241), .ZN(n92) );
  AOI22_X1 U75 ( .A1(N355), .A2(n18), .B1(addr_w_6[2]), .B2(n16), .ZN(n241) );
  INV_X1 U76 ( .A(n196), .ZN(n128) );
  AOI22_X1 U77 ( .A1(N553), .A2(n18), .B1(addr_w_15[2]), .B2(n14), .ZN(n196)
         );
  INV_X1 U78 ( .A(n200), .ZN(n125) );
  AOI22_X1 U79 ( .A1(N532), .A2(n18), .B1(addr_w_14[3]), .B2(n16), .ZN(n200)
         );
  XOR2_X1 U80 ( .A(addr_w_14[3]), .B(\add_2453_S2/carry[3] ), .Z(N532) );
  INV_X1 U81 ( .A(n235), .ZN(n97) );
  AOI22_X1 U82 ( .A1(N378), .A2(n18), .B1(addr_w_7[3]), .B2(n16), .ZN(n235) );
  XOR2_X1 U83 ( .A(addr_w_7[3]), .B(\add_2397_S2/carry[3] ), .Z(N378) );
  INV_X1 U84 ( .A(n198), .ZN(n126) );
  AOI22_X1 U85 ( .A1(N551), .A2(n18), .B1(addr_w_15[0]), .B2(n15), .ZN(n198)
         );
  INV_X1 U86 ( .A(n243), .ZN(n90) );
  AOI22_X1 U87 ( .A1(N353), .A2(n18), .B1(addr_w_6[0]), .B2(n16), .ZN(n243) );
  INV_X1 U88 ( .A(n222), .ZN(n107) );
  AOI22_X1 U89 ( .A1(N442), .A2(n18), .B1(addr_w_10[1]), .B2(n15), .ZN(n222)
         );
  INV_X1 U90 ( .A(n245), .ZN(n89) );
  AOI22_X1 U91 ( .A1(N334), .A2(n18), .B1(addr_w_5[3]), .B2(n15), .ZN(n245) );
  XOR2_X1 U92 ( .A(addr_w_5[3]), .B(\add_2381_S2/carry[3] ), .Z(N334) );
  INV_X1 U93 ( .A(n238), .ZN(n94) );
  AOI22_X1 U94 ( .A1(N375), .A2(n18), .B1(addr_w_7[0]), .B2(n16), .ZN(n238) );
  INV_X1 U95 ( .A(n203), .ZN(n122) );
  AOI22_X1 U96 ( .A1(N529), .A2(n18), .B1(addr_w_14[0]), .B2(n15), .ZN(n203)
         );
  INV_X1 U97 ( .A(n266), .ZN(n72) );
  AOI22_X1 U98 ( .A1(N245), .A2(n194), .B1(addr_w_1[2]), .B2(n14), .ZN(n266)
         );
  INV_X1 U99 ( .A(n233), .ZN(n98) );
  AOI22_X1 U100 ( .A1(N397), .A2(n18), .B1(addr_w_8[0]), .B2(n16), .ZN(n233)
         );
  INV_X1 U101 ( .A(n271), .ZN(n68) );
  AOI22_X1 U102 ( .A1(N223), .A2(n194), .B1(addr_w_0[2]), .B2(n14), .ZN(n271)
         );
  INV_X1 U103 ( .A(n193), .ZN(n129) );
  AOI22_X1 U104 ( .A1(N554), .A2(n18), .B1(addr_w_15[3]), .B2(n16), .ZN(n193)
         );
  XOR2_X1 U105 ( .A(addr_w_15[3]), .B(\add_2461_S2/carry[3] ), .Z(N554) );
  INV_X1 U106 ( .A(n236), .ZN(n96) );
  AOI22_X1 U107 ( .A1(N377), .A2(n18), .B1(addr_w_7[2]), .B2(n16), .ZN(n236)
         );
  INV_X1 U108 ( .A(n255), .ZN(n81) );
  AOI22_X1 U109 ( .A1(N290), .A2(n17), .B1(addr_w_3[3]), .B2(n15), .ZN(n255)
         );
  XOR2_X1 U110 ( .A(addr_w_3[3]), .B(\add_2365_S2/carry[3] ), .Z(N290) );
  INV_X1 U111 ( .A(n240), .ZN(n93) );
  AOI22_X1 U112 ( .A1(N356), .A2(n18), .B1(addr_w_6[3]), .B2(n16), .ZN(n240)
         );
  XOR2_X1 U113 ( .A(addr_w_6[3]), .B(\add_2389_S2/carry[3] ), .Z(N356) );
  INV_X1 U114 ( .A(n268), .ZN(n70) );
  AOI22_X1 U115 ( .A1(N243), .A2(n194), .B1(addr_w_1[0]), .B2(n14), .ZN(n268)
         );
  INV_X1 U116 ( .A(n215), .ZN(n113) );
  AOI22_X1 U117 ( .A1(N466), .A2(n17), .B1(addr_w_11[3]), .B2(n14), .ZN(n215)
         );
  XOR2_X1 U118 ( .A(addr_w_11[3]), .B(\add_2429_S2/carry[3] ), .Z(N466) );
  INV_X1 U119 ( .A(n217), .ZN(n111) );
  AOI22_X1 U120 ( .A1(N464), .A2(n17), .B1(addr_w_11[1]), .B2(n16), .ZN(n217)
         );
  INV_X1 U121 ( .A(n228), .ZN(n102) );
  AOI22_X1 U122 ( .A1(N419), .A2(n18), .B1(addr_w_9[0]), .B2(n15), .ZN(n228)
         );
  INV_X1 U123 ( .A(n206), .ZN(n120) );
  AOI22_X1 U124 ( .A1(N509), .A2(n17), .B1(addr_w_13[2]), .B2(n14), .ZN(n206)
         );
  INV_X1 U125 ( .A(n247), .ZN(n87) );
  AOI22_X1 U126 ( .A1(N332), .A2(n17), .B1(addr_w_5[1]), .B2(n15), .ZN(n247)
         );
  INV_X1 U127 ( .A(n212), .ZN(n115) );
  AOI22_X1 U128 ( .A1(N486), .A2(n18), .B1(addr_w_12[1]), .B2(n16), .ZN(n212)
         );
  INV_X1 U129 ( .A(n201), .ZN(n124) );
  AOI22_X1 U130 ( .A1(N531), .A2(n17), .B1(addr_w_14[2]), .B2(n14), .ZN(n201)
         );
  INV_X1 U131 ( .A(n261), .ZN(n76) );
  AOI22_X1 U132 ( .A1(N267), .A2(n194), .B1(addr_w_2[2]), .B2(n14), .ZN(n261)
         );
  INV_X1 U133 ( .A(n226), .ZN(n104) );
  AOI22_X1 U134 ( .A1(N421), .A2(n18), .B1(addr_w_9[2]), .B2(n14), .ZN(n226)
         );
  INV_X1 U135 ( .A(n272), .ZN(n67) );
  AOI22_X1 U136 ( .A1(N222), .A2(n194), .B1(addr_w_0[1]), .B2(n14), .ZN(n272)
         );
  INV_X1 U137 ( .A(n252), .ZN(n83) );
  AOI22_X1 U138 ( .A1(N310), .A2(n17), .B1(addr_w_4[1]), .B2(n15), .ZN(n252)
         );
  INV_X1 U139 ( .A(n270), .ZN(n69) );
  AOI22_X1 U140 ( .A1(N224), .A2(n194), .B1(addr_w_0[3]), .B2(n14), .ZN(n270)
         );
  XOR2_X1 U141 ( .A(addr_w_0[3]), .B(\add_2341_S2/carry[3] ), .Z(N224) );
  INV_X1 U142 ( .A(n258), .ZN(n78) );
  AOI22_X1 U143 ( .A1(N287), .A2(n17), .B1(addr_w_3[0]), .B2(n15), .ZN(n258)
         );
  INV_X1 U144 ( .A(n208), .ZN(n118) );
  AOI22_X1 U145 ( .A1(N507), .A2(n17), .B1(addr_w_13[0]), .B2(n15), .ZN(n208)
         );
  INV_X1 U146 ( .A(n216), .ZN(n112) );
  AOI22_X1 U147 ( .A1(N465), .A2(n17), .B1(addr_w_11[2]), .B2(n16), .ZN(n216)
         );
  INV_X1 U148 ( .A(n197), .ZN(n127) );
  AOI22_X1 U149 ( .A1(N552), .A2(n17), .B1(addr_w_15[1]), .B2(n14), .ZN(n197)
         );
  INV_X1 U150 ( .A(n242), .ZN(n91) );
  AOI22_X1 U151 ( .A1(N354), .A2(n18), .B1(addr_w_6[1]), .B2(n16), .ZN(n242)
         );
  INV_X1 U152 ( .A(n232), .ZN(n99) );
  AOI22_X1 U153 ( .A1(N398), .A2(n18), .B1(addr_w_8[1]), .B2(n16), .ZN(n232)
         );
  INV_X1 U154 ( .A(n220), .ZN(n109) );
  AOI22_X1 U155 ( .A1(N444), .A2(n18), .B1(addr_w_10[3]), .B2(n15), .ZN(n220)
         );
  XOR2_X1 U156 ( .A(addr_w_10[3]), .B(\add_2421_S2/carry[3] ), .Z(N444) );
  INV_X1 U157 ( .A(n237), .ZN(n95) );
  AOI22_X1 U158 ( .A1(N376), .A2(n18), .B1(addr_w_7[1]), .B2(n16), .ZN(n237)
         );
  INV_X1 U159 ( .A(n248), .ZN(n86) );
  AOI22_X1 U160 ( .A1(N331), .A2(n17), .B1(addr_w_5[0]), .B2(n15), .ZN(n248)
         );
  INV_X1 U161 ( .A(n263), .ZN(n74) );
  AOI22_X1 U162 ( .A1(N265), .A2(n194), .B1(addr_w_2[0]), .B2(n14), .ZN(n263)
         );
  INV_X1 U163 ( .A(n267), .ZN(n71) );
  AOI22_X1 U164 ( .A1(N244), .A2(n194), .B1(addr_w_1[1]), .B2(n14), .ZN(n267)
         );
  INV_X1 U165 ( .A(n227), .ZN(n103) );
  AOI22_X1 U166 ( .A1(N420), .A2(n194), .B1(addr_w_9[1]), .B2(n195), .ZN(n227)
         );
  INV_X1 U167 ( .A(n207), .ZN(n119) );
  AOI22_X1 U168 ( .A1(N508), .A2(n18), .B1(addr_w_13[1]), .B2(n14), .ZN(n207)
         );
  INV_X1 U169 ( .A(n260), .ZN(n77) );
  AOI22_X1 U170 ( .A1(N268), .A2(n17), .B1(addr_w_2[3]), .B2(n14), .ZN(n260)
         );
  XOR2_X1 U171 ( .A(addr_w_2[3]), .B(\add_2357_S2/carry[3] ), .Z(N268) );
  INV_X1 U172 ( .A(n246), .ZN(n88) );
  AOI22_X1 U173 ( .A1(N333), .A2(n17), .B1(addr_w_5[2]), .B2(n15), .ZN(n246)
         );
  INV_X1 U174 ( .A(n231), .ZN(n100) );
  AOI22_X1 U175 ( .A1(N399), .A2(n18), .B1(addr_w_8[2]), .B2(n16), .ZN(n231)
         );
  INV_X1 U176 ( .A(n230), .ZN(n101) );
  AOI22_X1 U177 ( .A1(N400), .A2(n17), .B1(addr_w_8[3]), .B2(n16), .ZN(n230)
         );
  XOR2_X1 U178 ( .A(addr_w_8[3]), .B(\add_2405_S2/carry[3] ), .Z(N400) );
  INV_X1 U179 ( .A(n221), .ZN(n108) );
  AOI22_X1 U180 ( .A1(N443), .A2(n194), .B1(addr_w_10[2]), .B2(n195), .ZN(n221) );
  INV_X1 U181 ( .A(n225), .ZN(n105) );
  AOI22_X1 U182 ( .A1(N422), .A2(n194), .B1(addr_w_9[3]), .B2(n195), .ZN(n225)
         );
  XOR2_X1 U183 ( .A(addr_w_9[3]), .B(\add_2413_S2/carry[3] ), .Z(N422) );
  INV_X1 U184 ( .A(n205), .ZN(n121) );
  AOI22_X1 U185 ( .A1(N510), .A2(n18), .B1(addr_w_13[3]), .B2(n16), .ZN(n205)
         );
  XOR2_X1 U186 ( .A(addr_w_13[3]), .B(\add_2445_S2/carry[3] ), .Z(N510) );
  INV_X1 U187 ( .A(n262), .ZN(n75) );
  AOI22_X1 U188 ( .A1(N266), .A2(n194), .B1(addr_w_2[1]), .B2(n14), .ZN(n262)
         );
  INV_X1 U189 ( .A(n210), .ZN(n117) );
  AOI22_X1 U190 ( .A1(N488), .A2(n17), .B1(addr_w_12[3]), .B2(n16), .ZN(n210)
         );
  XOR2_X1 U191 ( .A(addr_w_12[3]), .B(\add_2437_S2/carry[3] ), .Z(N488) );
  INV_X1 U192 ( .A(n211), .ZN(n116) );
  AOI22_X1 U193 ( .A1(N487), .A2(n17), .B1(addr_w_12[2]), .B2(n15), .ZN(n211)
         );
  INV_X1 U194 ( .A(n265), .ZN(n73) );
  AOI22_X1 U195 ( .A1(N246), .A2(n194), .B1(addr_w_1[3]), .B2(n14), .ZN(n265)
         );
  XOR2_X1 U196 ( .A(addr_w_1[3]), .B(\add_2349_S2/carry[3] ), .Z(N246) );
  INV_X1 U197 ( .A(n284), .ZN(n65) );
  AOI22_X1 U198 ( .A1(n285), .A2(addr_x[1]), .B1(n28), .B2(n283), .ZN(n284) );
  INV_X1 U199 ( .A(n202), .ZN(n123) );
  AOI22_X1 U200 ( .A1(N530), .A2(n18), .B1(addr_w_14[1]), .B2(n14), .ZN(n202)
         );
  INV_X1 U201 ( .A(n257), .ZN(n79) );
  AOI22_X1 U202 ( .A1(N288), .A2(n17), .B1(addr_w_3[1]), .B2(n15), .ZN(n257)
         );
  INV_X1 U203 ( .A(reset), .ZN(n62) );
  OAI21_X1 U204 ( .B1(n176), .B2(n295), .A(n296), .ZN(n343) );
  INV_X1 U205 ( .A(n155), .ZN(n21) );
  NAND2_X1 U206 ( .A1(n289), .A2(n21), .ZN(n19) );
  NAND2_X1 U207 ( .A1(n288), .A2(n19), .ZN(n338) );
  OAI21_X1 U208 ( .B1(n281), .B2(n156), .A(n282), .ZN(n336) );
  NAND3_X1 U209 ( .A1(n152), .A2(n151), .A3(n153), .ZN(n54) );
  INV_X1 U210 ( .A(s_valid), .ZN(n26) );
  NAND2_X1 U211 ( .A1(n13), .A2(n153), .ZN(n35) );
  INV_X1 U212 ( .A(n156), .ZN(n20) );
  NAND2_X1 U213 ( .A1(n21), .A2(n20), .ZN(n27) );
  NAND2_X1 U214 ( .A1(n132), .A2(sel[0]), .ZN(n38) );
  INV_X1 U215 ( .A(n40), .ZN(n22) );
  NAND4_X1 U216 ( .A1(n177), .A2(m_valid), .A3(m_ready), .A4(n22), .ZN(n23) );
  NAND2_X1 U217 ( .A1(n13), .A2(state[0]), .ZN(n130) );
  INV_X1 U218 ( .A(n130), .ZN(n61) );
  NAND2_X1 U219 ( .A1(n23), .A2(n61), .ZN(n45) );
  INV_X1 U220 ( .A(n45), .ZN(n24) );
  AOI21_X1 U221 ( .B1(n12), .B2(n27), .A(n24), .ZN(n25) );
  OAI211_X1 U222 ( .C1(n54), .C2(n26), .A(n35), .B(n25), .ZN(n47) );
  INV_X1 U223 ( .A(n47), .ZN(n33) );
  INV_X1 U224 ( .A(n27), .ZN(n42) );
  INV_X1 U225 ( .A(addr_x[3]), .ZN(n30) );
  NOR3_X1 U226 ( .A1(n30), .A2(n29), .A3(n28), .ZN(n31) );
  OAI21_X1 U227 ( .B1(n42), .B2(n31), .A(n11), .ZN(n32) );
  NAND2_X1 U228 ( .A1(n33), .A2(n32), .ZN(n52) );
  INV_X1 U229 ( .A(n52), .ZN(n34) );
  NOR2_X1 U230 ( .A1(reset), .A2(n34), .ZN(N11) );
  OR3_X1 U231 ( .A1(state[0]), .A2(n152), .A3(state[2]), .ZN(n57) );
  NAND2_X1 U232 ( .A1(n57), .A2(n35), .ZN(n43) );
  INV_X1 U233 ( .A(n43), .ZN(n36) );
  NAND3_X1 U234 ( .A1(m_ready), .A2(m_valid), .A3(n9), .ZN(n50) );
  NAND2_X1 U235 ( .A1(n9), .A2(n50), .ZN(n49) );
  OAI22_X1 U236 ( .A1(n186), .A2(n49), .B1(sel[0]), .B2(n50), .ZN(n344) );
  OAI22_X1 U237 ( .A1(n37), .A2(n50), .B1(n185), .B2(n49), .ZN(n341) );
  XOR2_X1 U238 ( .A(n38), .B(sel[2]), .Z(n39) );
  OAI22_X1 U239 ( .A1(n50), .A2(n39), .B1(n184), .B2(n49), .ZN(n340) );
  XOR2_X1 U240 ( .A(n40), .B(sel[4]), .Z(n41) );
  OAI221_X1 U241 ( .B1(n50), .B2(n41), .C1(n177), .C2(n49), .A(n62), .ZN(n342)
         );
  NAND3_X1 U242 ( .A1(state[0]), .A2(state[2]), .A3(n152), .ZN(n46) );
  NOR3_X1 U243 ( .A1(n7), .A2(n11), .A3(n43), .ZN(n44) );
  NAND3_X1 U244 ( .A1(n45), .A2(n46), .A3(n44), .ZN(n191) );
  INV_X1 U245 ( .A(n46), .ZN(n131) );
  INV_X1 U246 ( .A(n1), .ZN(n60) );
  XOR2_X1 U247 ( .A(n48), .B(sel[3]), .Z(n51) );
  OAI22_X1 U248 ( .A1(n51), .A2(n50), .B1(n183), .B2(n49), .ZN(n339) );
  INV_X1 U249 ( .A(n191), .ZN(n53) );
  INV_X1 U250 ( .A(n57), .ZN(n306) );
  INV_X1 U251 ( .A(\r444/GE_LT_GT_LE ), .ZN(n59) );
  INV_X1 U252 ( .A(n291), .ZN(n58) );
  OAI21_X1 U253 ( .B1(n8), .B2(wr_en_x), .A(n62), .ZN(n287) );
  INV_X1 U254 ( .A(n287), .ZN(n64) );
  AND4_X1 U255 ( .A1(sel[3]), .A2(sel[2]), .A3(n132), .A4(sel[0]), .ZN(n63) );
  NOR2_X1 U256 ( .A1(n63), .A2(sel[4]), .ZN(\r444/GE_LT_GT_LE ) );
endmodule


module layer3_16_12_16_16 ( clk, reset, s_valid, m_ready, data_in, m_valid, 
        s_ready, data_out );
  input [15:0] data_in;
  output [15:0] data_out;
  input clk, reset, s_valid, m_ready;
  output m_valid, s_ready;
  wire   wr_en_x, \addr_b_0[0] , \addr_b_1[0] , \addr_b_2[0] , \addr_b_3[0] ,
         \addr_b_4[0] , \addr_b_5[0] , \addr_b_6[0] , \addr_b_7[0] ,
         \addr_b_8[0] , \addr_b_9[0] , \addr_b_10[0] , \addr_b_11[0] ,
         \addr_b_12[0] , \addr_b_13[0] , \addr_b_14[0] , \addr_b_15[0] ,
         clear_acc, wr_en_y, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276;
  wire   [15:0] data_out_x;
  wire   [3:0] addr_x;
  wire   [3:0] addr_w_0;
  wire   [15:0] data_out_w_0;
  wire   [15:0] data_out_b_0;
  wire   [3:0] addr_w_1;
  wire   [15:0] data_out_w_1;
  wire   [15:0] data_out_b_1;
  wire   [3:0] addr_w_2;
  wire   [15:0] data_out_w_2;
  wire   [15:0] data_out_b_2;
  wire   [3:0] addr_w_3;
  wire   [15:0] data_out_w_3;
  wire   [15:0] data_out_b_3;
  wire   [3:0] addr_w_4;
  wire   [15:0] data_out_w_4;
  wire   [15:0] data_out_b_4;
  wire   [3:0] addr_w_5;
  wire   [15:0] data_out_w_5;
  wire   [15:0] data_out_b_5;
  wire   [3:0] addr_w_6;
  wire   [15:0] data_out_w_6;
  wire   [15:0] data_out_b_6;
  wire   [3:0] addr_w_7;
  wire   [15:0] data_out_w_7;
  wire   [15:0] data_out_b_7;
  wire   [3:0] addr_w_8;
  wire   [15:0] data_out_w_8;
  wire   [15:0] data_out_b_8;
  wire   [3:0] addr_w_9;
  wire   [15:0] data_out_w_9;
  wire   [15:0] data_out_b_9;
  wire   [3:0] addr_w_10;
  wire   [15:0] data_out_w_10;
  wire   [15:0] data_out_b_10;
  wire   [3:0] addr_w_11;
  wire   [15:0] data_out_w_11;
  wire   [15:0] data_out_b_11;
  wire   [3:0] addr_w_12;
  wire   [15:0] data_out_w_12;
  wire   [15:0] data_out_b_12;
  wire   [3:0] addr_w_13;
  wire   [15:0] data_out_w_13;
  wire   [15:0] data_out_b_13;
  wire   [3:0] addr_w_14;
  wire   [15:0] data_out_w_14;
  wire   [15:0] data_out_b_14;
  wire   [3:0] addr_w_15;
  wire   [15:0] data_out_w_15;
  wire   [15:0] data_out_b_15;
  wire   [15:0] data_out_0;
  wire   [4:0] sel;
  wire   [15:0] data_out_1;
  wire   [15:0] data_out_2;
  wire   [15:0] data_out_3;
  wire   [15:0] data_out_4;
  wire   [15:0] data_out_5;
  wire   [15:0] data_out_6;
  wire   [15:0] data_out_7;
  wire   [15:0] data_out_8;
  wire   [15:0] data_out_9;
  wire   [15:0] data_out_10;
  wire   [15:0] data_out_11;
  wire   [15:0] data_out_12;
  wire   [15:0] data_out_13;
  wire   [15:0] data_out_14;
  wire   [15:0] data_out_15;
  wire   SYNOPSYS_UNCONNECTED__0;

  memory_WIDTH16_SIZE12_LOGSIZE4 mem_x ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_x), .addr(addr_x), .wr_en(wr_en_x) );
  layer3_16_12_16_16_W_rom_0 mem_w_0 ( .clk(clk), .addr(addr_w_0), .z(
        data_out_w_0) );
  layer3_16_12_16_16_B_rom_0 mem_b_0 ( .clk(clk), .addr(\addr_b_0[0] ) );
  layer3_16_12_16_16_W_rom_1 mem_w_1 ( .clk(clk), .addr(addr_w_1), .z(
        data_out_w_1) );
  layer3_16_12_16_16_B_rom_1 mem_b_1 ( .clk(clk), .addr(\addr_b_1[0] ) );
  layer3_16_12_16_16_W_rom_2 mem_w_2 ( .clk(clk), .addr(addr_w_2), .z(
        data_out_w_2) );
  layer3_16_12_16_16_B_rom_2 mem_b_2 ( .clk(clk), .addr(\addr_b_2[0] ) );
  layer3_16_12_16_16_W_rom_3 mem_w_3 ( .clk(clk), .addr(addr_w_3), .z(
        data_out_w_3) );
  layer3_16_12_16_16_B_rom_3 mem_b_3 ( .clk(clk), .addr(\addr_b_3[0] ) );
  layer3_16_12_16_16_W_rom_4 mem_w_4 ( .clk(clk), .addr(addr_w_4), .z(
        data_out_w_4) );
  layer3_16_12_16_16_B_rom_4 mem_b_4 ( .clk(clk), .addr(\addr_b_4[0] ) );
  layer3_16_12_16_16_W_rom_5 mem_w_5 ( .clk(clk), .addr(addr_w_5), .z(
        data_out_w_5) );
  layer3_16_12_16_16_B_rom_5 mem_b_5 ( .clk(clk), .addr(\addr_b_5[0] ) );
  layer3_16_12_16_16_W_rom_6 mem_w_6 ( .clk(clk), .addr(addr_w_6), .z({
        data_out_w_6[15:5], SYNOPSYS_UNCONNECTED__0, data_out_w_6[3:0]}) );
  layer3_16_12_16_16_B_rom_6 mem_b_6 ( .clk(clk), .addr(\addr_b_6[0] ) );
  layer3_16_12_16_16_W_rom_7 mem_w_7 ( .clk(clk), .addr(addr_w_7), .z(
        data_out_w_7) );
  layer3_16_12_16_16_B_rom_7 mem_b_7 ( .clk(clk), .addr(\addr_b_7[0] ) );
  layer3_16_12_16_16_W_rom_8 mem_w_8 ( .clk(clk), .addr(addr_w_8), .z(
        data_out_w_8) );
  layer3_16_12_16_16_B_rom_8 mem_b_8 ( .clk(clk), .addr(\addr_b_8[0] ) );
  layer3_16_12_16_16_W_rom_9 mem_w_9 ( .clk(clk), .addr(addr_w_9), .z(
        data_out_w_9) );
  layer3_16_12_16_16_B_rom_9 mem_b_9 ( .clk(clk), .addr(\addr_b_9[0] ) );
  layer3_16_12_16_16_W_rom_10 mem_w_10 ( .clk(clk), .addr(addr_w_10), .z(
        data_out_w_10) );
  layer3_16_12_16_16_B_rom_10 mem_b_10 ( .clk(clk), .addr(\addr_b_10[0] ) );
  layer3_16_12_16_16_W_rom_11 mem_w_11 ( .clk(clk), .addr(addr_w_11), .z(
        data_out_w_11) );
  layer3_16_12_16_16_B_rom_11 mem_b_11 ( .clk(clk), .addr(\addr_b_11[0] ) );
  layer3_16_12_16_16_W_rom_12 mem_w_12 ( .clk(clk), .addr(addr_w_12), .z(
        data_out_w_12) );
  layer3_16_12_16_16_B_rom_12 mem_b_12 ( .clk(clk), .addr(\addr_b_12[0] ) );
  layer3_16_12_16_16_W_rom_13 mem_w_13 ( .clk(clk), .addr(addr_w_13), .z(
        data_out_w_13) );
  layer3_16_12_16_16_B_rom_13 mem_b_13 ( .clk(clk), .addr(\addr_b_13[0] ) );
  layer3_16_12_16_16_W_rom_14 mem_w_14 ( .clk(clk), .addr(addr_w_14), .z(
        data_out_w_14) );
  layer3_16_12_16_16_B_rom_14 mem_b_14 ( .clk(clk), .addr(\addr_b_14[0] ) );
  layer3_16_12_16_16_W_rom_15 mem_w_15 ( .clk(clk), .addr(addr_w_15), .z(
        data_out_w_15) );
  layer3_16_12_16_16_B_rom_15 mem_b_15 ( .clk(clk), .addr(\addr_b_15[0] ) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_0 d_0 ( .clk(clk), .clear_acc(
        n225), .data_out_x({n255, n5, n252, n251, n7, n246, n1, n243, n241, 
        n239, n236, n6, n232, n13, n229, n17}), .data_out(data_out_0), 
        .data_out_w(data_out_w_0), .data_out_b({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1}), 
        .wr_en_y(n224), .m_valid(m_valid), .m_ready(m_ready), .sel(sel) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_15 d_1 ( .clk(clk), .clear_acc(
        clear_acc), .data_out_x({n256, n4, n253, n250, n248, n246, n245, n242, 
        n3, n15, n9, n235, n11, n13, n221, n226}), .data_out(data_out_1), 
        .data_out_w(data_out_w_1), .data_out_b({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1}), 
        .wr_en_y(wr_en_y), .m_valid(m_valid), .m_ready(m_ready), .sel(sel) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_14 d_2 ( .clk(clk), .clear_acc(
        clear_acc), .data_out_x({n256, n4, n253, n250, n249, n12, n1, n243, n2, 
        n238, n236, n234, n232, n230, n222, n227}), .data_out(data_out_2), 
        .data_out_w(data_out_w_2), .data_out_b({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1}), 
        .wr_en_y(wr_en_y), .m_valid(m_valid), .m_ready(m_ready), .sel(sel) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_13 d_3 ( .clk(clk), .clear_acc(
        clear_acc), .data_out_x({n256, n5, n253, n250, n249, n247, n244, n16, 
        n2, n15, n236, n234, n11, n231, n221, n227}), .data_out(data_out_3), 
        .data_out_w(data_out_w_3), .data_out_b({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1}), 
        .wr_en_y(wr_en_y), .m_valid(m_valid), .m_ready(m_ready), .sel(sel) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_12 d_4 ( .clk(clk), .clear_acc(
        clear_acc), .data_out_x({n256, n4, n253, n250, n249, n12, n244, n243, 
        n3, n239, n9, n10, n233, n230, n229, n226}), .data_out(data_out_4), 
        .data_out_w(data_out_w_4), .data_out_b({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .wr_en_y(wr_en_y), .m_valid(m_valid), .m_ready(m_ready), .sel(sel) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_11 d_5 ( .clk(clk), .clear_acc(
        clear_acc), .data_out_x({n255, n5, n252, n250, n248, n246, n245, n242, 
        n2, n8, n236, n235, n233, n13, n228, n227}), .data_out(data_out_5), 
        .data_out_w(data_out_w_5), .data_out_b({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1}), 
        .wr_en_y(wr_en_y), .m_valid(m_valid), .m_ready(m_ready), .sel(sel) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_10 d_6 ( .clk(clk), .clear_acc(
        clear_acc), .data_out_x({n255, n4, n252, n250, n248, n246, n1, n242, 
        n240, n238, n236, n234, n232, n14, n228, n19}), .data_out(data_out_6), 
        .data_out_w({data_out_w_6[15:5], 1'b1, data_out_w_6[3:0]}), 
        .data_out_b({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1}), .wr_en_y(wr_en_y), 
        .m_valid(m_valid), .m_ready(m_ready), .sel(sel) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_9 d_7 ( .clk(clk), .clear_acc(
        clear_acc), .data_out_x({n255, n254, n252, n250, n7, n12, n245, n243, 
        n240, n239, n9, n10, n232, n14, n229, n18}), .data_out(data_out_7), 
        .data_out_w(data_out_w_7), .data_out_b({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0}), 
        .wr_en_y(wr_en_y), .m_valid(m_valid), .m_ready(m_ready), .sel(sel) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_8 d_8 ( .clk(clk), .clear_acc(
        clear_acc), .data_out_x({n255, n254, n252, n250, n248, n12, n245, n16, 
        n3, n15, n9, n235, n233, n14, n228, n18}), .data_out(data_out_8), 
        .data_out_w(data_out_w_8), .data_out_b({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0}), 
        .wr_en_y(wr_en_y), .m_valid(m_valid), .m_ready(m_ready), .sel(sel) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_7 d_9 ( .clk(clk), .clear_acc(
        clear_acc), .data_out_x({n255, n4, n252, n250, n248, n247, n1, n243, 
        n241, n8, n9, n6, n11, n231, n229, n17}), .data_out(data_out_9), 
        .data_out_w(data_out_w_9), .data_out_b({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), 
        .wr_en_y(wr_en_y), .m_valid(m_valid), .m_ready(m_ready), .sel(sel) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_6 d_10 ( .clk(clk), .clear_acc(
        clear_acc), .data_out_x({n255, n254, n252, n250, n7, n247, n1, n16, n2, 
        n15, n9, n10, n11, n231, n222, n19}), .data_out(data_out_10), 
        .data_out_w(data_out_w_10), .data_out_b({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0}), 
        .wr_en_y(n224), .m_valid(m_valid), .m_ready(m_ready), .sel(sel) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_5 d_11 ( .clk(clk), .clear_acc(
        clear_acc), .data_out_x({n255, n5, n252, n250, n248, n246, n1, n16, 
        n241, n8, n237, n10, n11, n14, n228, n18}), .data_out(data_out_11), 
        .data_out_w(data_out_w_11), .data_out_b({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1}), 
        .wr_en_y(n224), .m_valid(m_valid), .m_ready(m_ready), .sel(sel) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_4 d_12 ( .clk(clk), .clear_acc(
        clear_acc), .data_out_x({n255, n4, n252, n250, n7, n12, n1, n242, n3, 
        n15, n9, n6, n11, n230, n20, n17}), .data_out(data_out_12), 
        .data_out_w(data_out_w_12), .data_out_b({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1}), 
        .wr_en_y(n224), .m_valid(m_valid), .m_ready(m_ready), .sel(sel) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_3 d_13 ( .clk(clk), .clear_acc(
        n225), .data_out_x({n255, n4, n252, n251, n248, n247, n244, n242, n2, 
        n8, n237, n234, n233, n230, n222, n17}), .data_out(data_out_13), 
        .data_out_w(data_out_w_13), .data_out_b({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1}), 
        .wr_en_y(n224), .m_valid(m_valid), .m_ready(m_ready), .sel(sel) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_2 d_14 ( .clk(clk), .clear_acc(
        n225), .data_out_x({n255, n5, n252, n251, n7, n247, n245, n243, n240, 
        n8, n237, n6, n233, n231, n221, n19}), .data_out(data_out_14), 
        .data_out_w(data_out_w_14), .data_out_b({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0}), 
        .wr_en_y(n224), .m_valid(m_valid), .m_ready(m_ready), .sel(sel) );
  layer3_16_12_16_16_datapath_M16_N12_T16_P16_1 d_15 ( .clk(clk), .clear_acc(
        n225), .data_out_x({n255, n5, n252, n251, n7, n247, n244, n16, n3, 
        n239, n237, n6, n11, n13, n229, n226}), .data_out(data_out_15), 
        .data_out_w(data_out_w_15), .data_out_b({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0}), 
        .wr_en_y(n224), .m_valid(m_valid), .m_ready(m_ready), .sel(sel) );
  layer3_16_12_16_16_ctrlpath_M16_N12_T16_P16 c ( .clk(clk), .reset(reset), 
        .s_valid(s_valid), .s_ready(s_ready), .m_valid(m_valid), .m_ready(
        m_ready), .clear_acc(clear_acc), .wr_en_x(wr_en_x), .wr_en_y(wr_en_y), 
        .sel(sel), .addr_x(addr_x), .addr_w_0(addr_w_0), .addr_b_0(
        \addr_b_0[0] ), .addr_w_1(addr_w_1), .addr_b_1(\addr_b_1[0] ), 
        .addr_w_2(addr_w_2), .addr_b_2(\addr_b_2[0] ), .addr_w_3(addr_w_3), 
        .addr_b_3(\addr_b_3[0] ), .addr_w_4(addr_w_4), .addr_b_4(\addr_b_4[0] ), .addr_w_5(addr_w_5), .addr_b_5(\addr_b_5[0] ), .addr_w_6(addr_w_6), 
        .addr_b_6(\addr_b_6[0] ), .addr_w_7(addr_w_7), .addr_b_7(\addr_b_7[0] ), .addr_w_8(addr_w_8), .addr_b_8(\addr_b_8[0] ), .addr_w_9(addr_w_9), 
        .addr_b_9(\addr_b_9[0] ), .addr_w_10(addr_w_10), .addr_b_10(
        \addr_b_10[0] ), .addr_w_11(addr_w_11), .addr_b_11(\addr_b_11[0] ), 
        .addr_w_12(addr_w_12), .addr_b_12(\addr_b_12[0] ), .addr_w_13(
        addr_w_13), .addr_b_13(\addr_b_13[0] ), .addr_w_14(addr_w_14), 
        .addr_b_14(\addr_b_14[0] ), .addr_w_15(addr_w_15), .addr_b_15(
        \addr_b_15[0] ) );
  CLKBUF_X3 U1 ( .A(data_out_x[9]), .Z(n1) );
  CLKBUF_X2 U2 ( .A(data_out_x[9]), .Z(n244) );
  CLKBUF_X3 U3 ( .A(data_out_x[0]), .Z(n19) );
  CLKBUF_X3 U4 ( .A(data_out_x[5]), .Z(n236) );
  BUF_X2 U5 ( .A(data_out_x[7]), .Z(n2) );
  BUF_X2 U6 ( .A(data_out_x[7]), .Z(n3) );
  BUF_X1 U7 ( .A(data_out_x[7]), .Z(n241) );
  BUF_X1 U8 ( .A(data_out_x[1]), .Z(n222) );
  CLKBUF_X3 U9 ( .A(data_out_x[1]), .Z(n229) );
  BUF_X1 U10 ( .A(data_out_x[1]), .Z(n228) );
  CLKBUF_X3 U11 ( .A(data_out_x[10]), .Z(n246) );
  CLKBUF_X3 U12 ( .A(data_out_x[10]), .Z(n247) );
  CLKBUF_X3 U13 ( .A(data_out_x[4]), .Z(n234) );
  CLKBUF_X3 U14 ( .A(data_out_x[8]), .Z(n243) );
  BUF_X2 U15 ( .A(data_out_x[3]), .Z(n11) );
  CLKBUF_X3 U16 ( .A(data_out_x[2]), .Z(n231) );
  CLKBUF_X3 U17 ( .A(data_out_x[14]), .Z(n4) );
  CLKBUF_X3 U18 ( .A(data_out_x[14]), .Z(n5) );
  CLKBUF_X1 U19 ( .A(data_out_x[14]), .Z(n254) );
  CLKBUF_X3 U20 ( .A(data_out_x[4]), .Z(n6) );
  CLKBUF_X2 U21 ( .A(data_out_x[4]), .Z(n10) );
  CLKBUF_X3 U22 ( .A(data_out_x[11]), .Z(n7) );
  BUF_X2 U23 ( .A(data_out_x[6]), .Z(n238) );
  BUF_X2 U24 ( .A(n222), .Z(n20) );
  CLKBUF_X3 U25 ( .A(data_out_x[8]), .Z(n242) );
  CLKBUF_X3 U26 ( .A(data_out_x[6]), .Z(n8) );
  BUF_X2 U27 ( .A(data_out_x[5]), .Z(n9) );
  CLKBUF_X3 U28 ( .A(data_out_x[3]), .Z(n233) );
  CLKBUF_X3 U29 ( .A(data_out_x[0]), .Z(n227) );
  CLKBUF_X3 U30 ( .A(data_out_x[15]), .Z(n255) );
  CLKBUF_X3 U31 ( .A(data_out_x[2]), .Z(n13) );
  CLKBUF_X3 U32 ( .A(data_out_x[4]), .Z(n235) );
  CLKBUF_X3 U33 ( .A(data_out_x[2]), .Z(n230) );
  CLKBUF_X3 U34 ( .A(data_out_x[10]), .Z(n12) );
  CLKBUF_X3 U35 ( .A(data_out_x[2]), .Z(n14) );
  CLKBUF_X3 U36 ( .A(data_out_x[6]), .Z(n15) );
  CLKBUF_X3 U37 ( .A(data_out_x[8]), .Z(n16) );
  CLKBUF_X3 U38 ( .A(data_out_x[0]), .Z(n17) );
  CLKBUF_X3 U39 ( .A(data_out_x[0]), .Z(n18) );
  CLKBUF_X3 U40 ( .A(data_out_x[0]), .Z(n226) );
  BUF_X2 U41 ( .A(data_out_x[7]), .Z(n240) );
  CLKBUF_X3 U42 ( .A(data_out_x[6]), .Z(n239) );
  CLKBUF_X3 U43 ( .A(data_out_x[3]), .Z(n232) );
  BUF_X1 U44 ( .A(data_out_x[1]), .Z(n221) );
  NOR2_X1 U45 ( .A1(n276), .A2(n273), .ZN(n220) );
  AND2_X1 U46 ( .A1(n214), .A2(n220), .ZN(n46) );
  AND2_X1 U47 ( .A1(n213), .A2(n220), .ZN(n44) );
  AND2_X1 U48 ( .A1(n211), .A2(n212), .ZN(n30) );
  AND2_X1 U49 ( .A1(n211), .A2(n213), .ZN(n32) );
  AND2_X1 U50 ( .A1(n211), .A2(n210), .ZN(n28) );
  AND2_X1 U51 ( .A1(n211), .A2(n214), .ZN(n34) );
  AND2_X1 U52 ( .A1(n210), .A2(n220), .ZN(n40) );
  AND2_X1 U53 ( .A1(n212), .A2(n220), .ZN(n42) );
  AND2_X1 U54 ( .A1(n214), .A2(n219), .ZN(n47) );
  AND2_X1 U55 ( .A1(n219), .A2(n210), .ZN(n41) );
  AND2_X1 U56 ( .A1(n213), .A2(n219), .ZN(n45) );
  AND2_X1 U57 ( .A1(n209), .A2(n212), .ZN(n31) );
  AND2_X1 U58 ( .A1(n209), .A2(n213), .ZN(n33) );
  AND2_X1 U59 ( .A1(n209), .A2(n210), .ZN(n29) );
  AND2_X1 U60 ( .A1(n209), .A2(n214), .ZN(n35) );
  AND2_X1 U61 ( .A1(n212), .A2(n219), .ZN(n43) );
  BUF_X1 U62 ( .A(n274), .Z(n223) );
  NOR2_X1 U63 ( .A1(sel[2]), .A2(sel[1]), .ZN(n214) );
  NOR2_X1 U64 ( .A1(n275), .A2(sel[2]), .ZN(n213) );
  NOR2_X1 U65 ( .A1(n276), .A2(sel[0]), .ZN(n219) );
  NOR2_X1 U66 ( .A1(sel[3]), .A2(sel[0]), .ZN(n209) );
  NOR2_X1 U67 ( .A1(n273), .A2(sel[3]), .ZN(n211) );
  BUF_X4 U68 ( .A(data_out_x[12]), .Z(n250) );
  BUF_X2 U69 ( .A(data_out_x[12]), .Z(n251) );
  AOI22_X1 U70 ( .A1(data_out_15[0]), .A2(n40), .B1(data_out_14[0]), .B2(n41), 
        .ZN(n218) );
  AOI22_X1 U71 ( .A1(data_out_15[1]), .A2(n40), .B1(data_out_14[1]), .B2(n41), 
        .ZN(n135) );
  AOI22_X1 U72 ( .A1(data_out_15[2]), .A2(n40), .B1(data_out_14[2]), .B2(n41), 
        .ZN(n124) );
  AOI22_X1 U73 ( .A1(data_out_15[3]), .A2(n40), .B1(data_out_14[3]), .B2(n41), 
        .ZN(n113) );
  AOI22_X1 U74 ( .A1(data_out_15[4]), .A2(n40), .B1(data_out_14[4]), .B2(n41), 
        .ZN(n102) );
  AOI22_X1 U75 ( .A1(data_out_15[5]), .A2(n40), .B1(data_out_14[5]), .B2(n41), 
        .ZN(n91) );
  AOI22_X1 U76 ( .A1(data_out_15[6]), .A2(n40), .B1(data_out_14[6]), .B2(n41), 
        .ZN(n80) );
  AOI22_X1 U77 ( .A1(data_out_15[7]), .A2(n40), .B1(data_out_14[7]), .B2(n41), 
        .ZN(n69) );
  AOI22_X1 U78 ( .A1(data_out_15[8]), .A2(n40), .B1(data_out_14[8]), .B2(n41), 
        .ZN(n58) );
  AOI22_X1 U79 ( .A1(data_out_15[9]), .A2(n40), .B1(data_out_14[9]), .B2(n41), 
        .ZN(n39) );
  AOI22_X1 U80 ( .A1(data_out_15[10]), .A2(n40), .B1(data_out_14[10]), .B2(n41), .ZN(n201) );
  AOI22_X1 U81 ( .A1(data_out_15[11]), .A2(n40), .B1(data_out_14[11]), .B2(n41), .ZN(n190) );
  AOI22_X1 U82 ( .A1(data_out_15[12]), .A2(n40), .B1(data_out_14[12]), .B2(n41), .ZN(n179) );
  AOI22_X1 U83 ( .A1(data_out_15[13]), .A2(n40), .B1(data_out_14[13]), .B2(n41), .ZN(n168) );
  AOI22_X1 U84 ( .A1(data_out_15[14]), .A2(n40), .B1(data_out_14[14]), .B2(n41), .ZN(n157) );
  AOI22_X1 U85 ( .A1(data_out_15[15]), .A2(n40), .B1(data_out_14[15]), .B2(n41), .ZN(n146) );
  AOI22_X1 U86 ( .A1(data_out_5[0]), .A2(n30), .B1(data_out_4[0]), .B2(n31), 
        .ZN(n207) );
  AOI22_X1 U87 ( .A1(data_out_13[0]), .A2(n42), .B1(data_out_12[0]), .B2(n43), 
        .ZN(n217) );
  AOI22_X1 U88 ( .A1(data_out_5[1]), .A2(n30), .B1(data_out_4[1]), .B2(n31), 
        .ZN(n130) );
  AOI22_X1 U89 ( .A1(data_out_13[1]), .A2(n42), .B1(data_out_12[1]), .B2(n43), 
        .ZN(n134) );
  AOI22_X1 U90 ( .A1(data_out_5[2]), .A2(n30), .B1(data_out_4[2]), .B2(n31), 
        .ZN(n119) );
  AOI22_X1 U91 ( .A1(data_out_13[2]), .A2(n42), .B1(data_out_12[2]), .B2(n43), 
        .ZN(n123) );
  AOI22_X1 U92 ( .A1(data_out_5[3]), .A2(n30), .B1(data_out_4[3]), .B2(n31), 
        .ZN(n108) );
  AOI22_X1 U93 ( .A1(data_out_13[3]), .A2(n42), .B1(data_out_12[3]), .B2(n43), 
        .ZN(n112) );
  AOI22_X1 U94 ( .A1(data_out_5[4]), .A2(n30), .B1(data_out_4[4]), .B2(n31), 
        .ZN(n97) );
  AOI22_X1 U95 ( .A1(data_out_13[4]), .A2(n42), .B1(data_out_12[4]), .B2(n43), 
        .ZN(n101) );
  AOI22_X1 U96 ( .A1(data_out_5[5]), .A2(n30), .B1(data_out_4[5]), .B2(n31), 
        .ZN(n86) );
  AOI22_X1 U97 ( .A1(data_out_13[5]), .A2(n42), .B1(data_out_12[5]), .B2(n43), 
        .ZN(n90) );
  AOI22_X1 U98 ( .A1(data_out_5[6]), .A2(n30), .B1(data_out_4[6]), .B2(n31), 
        .ZN(n75) );
  AOI22_X1 U99 ( .A1(data_out_13[6]), .A2(n42), .B1(data_out_12[6]), .B2(n43), 
        .ZN(n79) );
  AOI22_X1 U100 ( .A1(data_out_5[7]), .A2(n30), .B1(data_out_4[7]), .B2(n31), 
        .ZN(n64) );
  AOI22_X1 U101 ( .A1(data_out_13[7]), .A2(n42), .B1(data_out_12[7]), .B2(n43), 
        .ZN(n68) );
  AOI22_X1 U102 ( .A1(data_out_5[8]), .A2(n30), .B1(data_out_4[8]), .B2(n31), 
        .ZN(n53) );
  AOI22_X1 U103 ( .A1(data_out_13[8]), .A2(n42), .B1(data_out_12[8]), .B2(n43), 
        .ZN(n57) );
  AOI22_X1 U104 ( .A1(data_out_5[9]), .A2(n30), .B1(data_out_4[9]), .B2(n31), 
        .ZN(n26) );
  AOI22_X1 U105 ( .A1(data_out_13[9]), .A2(n42), .B1(data_out_12[9]), .B2(n43), 
        .ZN(n38) );
  AOI22_X1 U106 ( .A1(data_out_5[10]), .A2(n30), .B1(data_out_4[10]), .B2(n31), 
        .ZN(n196) );
  AOI22_X1 U107 ( .A1(data_out_13[10]), .A2(n42), .B1(data_out_12[10]), .B2(
        n43), .ZN(n200) );
  AOI22_X1 U108 ( .A1(data_out_5[11]), .A2(n30), .B1(data_out_4[11]), .B2(n31), 
        .ZN(n185) );
  AOI22_X1 U109 ( .A1(data_out_13[11]), .A2(n42), .B1(data_out_12[11]), .B2(
        n43), .ZN(n189) );
  AOI22_X1 U110 ( .A1(data_out_5[12]), .A2(n30), .B1(data_out_4[12]), .B2(n31), 
        .ZN(n174) );
  AOI22_X1 U111 ( .A1(data_out_13[12]), .A2(n42), .B1(data_out_12[12]), .B2(
        n43), .ZN(n178) );
  AOI22_X1 U112 ( .A1(data_out_5[13]), .A2(n30), .B1(data_out_4[13]), .B2(n31), 
        .ZN(n163) );
  AOI22_X1 U113 ( .A1(data_out_13[13]), .A2(n42), .B1(data_out_12[13]), .B2(
        n43), .ZN(n167) );
  AOI22_X1 U114 ( .A1(data_out_5[14]), .A2(n30), .B1(data_out_4[14]), .B2(n31), 
        .ZN(n152) );
  AOI22_X1 U115 ( .A1(data_out_13[14]), .A2(n42), .B1(data_out_12[14]), .B2(
        n43), .ZN(n156) );
  AOI22_X1 U116 ( .A1(data_out_5[15]), .A2(n30), .B1(data_out_4[15]), .B2(n31), 
        .ZN(n141) );
  AOI22_X1 U117 ( .A1(data_out_13[15]), .A2(n42), .B1(data_out_12[15]), .B2(
        n43), .ZN(n145) );
  AOI22_X1 U118 ( .A1(data_out_11[0]), .A2(n44), .B1(data_out_10[0]), .B2(n45), 
        .ZN(n216) );
  AOI22_X1 U119 ( .A1(data_out_11[1]), .A2(n44), .B1(data_out_10[1]), .B2(n45), 
        .ZN(n133) );
  AOI22_X1 U120 ( .A1(data_out_11[2]), .A2(n44), .B1(data_out_10[2]), .B2(n45), 
        .ZN(n122) );
  AOI22_X1 U121 ( .A1(data_out_11[3]), .A2(n44), .B1(data_out_10[3]), .B2(n45), 
        .ZN(n111) );
  AOI22_X1 U122 ( .A1(data_out_11[4]), .A2(n44), .B1(data_out_10[4]), .B2(n45), 
        .ZN(n100) );
  AOI22_X1 U123 ( .A1(data_out_11[5]), .A2(n44), .B1(data_out_10[5]), .B2(n45), 
        .ZN(n89) );
  AOI22_X1 U124 ( .A1(data_out_11[6]), .A2(n44), .B1(data_out_10[6]), .B2(n45), 
        .ZN(n78) );
  AOI22_X1 U125 ( .A1(data_out_11[7]), .A2(n44), .B1(data_out_10[7]), .B2(n45), 
        .ZN(n67) );
  AOI22_X1 U126 ( .A1(data_out_11[8]), .A2(n44), .B1(data_out_10[8]), .B2(n45), 
        .ZN(n56) );
  AOI22_X1 U127 ( .A1(data_out_11[9]), .A2(n44), .B1(data_out_10[9]), .B2(n45), 
        .ZN(n37) );
  AOI22_X1 U128 ( .A1(data_out_11[10]), .A2(n44), .B1(data_out_10[10]), .B2(
        n45), .ZN(n199) );
  AOI22_X1 U129 ( .A1(data_out_11[11]), .A2(n44), .B1(data_out_10[11]), .B2(
        n45), .ZN(n188) );
  AOI22_X1 U130 ( .A1(data_out_11[12]), .A2(n44), .B1(data_out_10[12]), .B2(
        n45), .ZN(n177) );
  AOI22_X1 U131 ( .A1(data_out_11[13]), .A2(n44), .B1(data_out_10[13]), .B2(
        n45), .ZN(n166) );
  AOI22_X1 U132 ( .A1(data_out_11[14]), .A2(n44), .B1(data_out_10[14]), .B2(
        n45), .ZN(n155) );
  AOI22_X1 U133 ( .A1(data_out_11[15]), .A2(n44), .B1(data_out_10[15]), .B2(
        n45), .ZN(n144) );
  INV_X1 U134 ( .A(sel[4]), .ZN(n274) );
  AOI22_X1 U135 ( .A1(data_out_9[0]), .A2(n46), .B1(data_out_8[0]), .B2(n47), 
        .ZN(n215) );
  AOI22_X1 U136 ( .A1(data_out_9[1]), .A2(n46), .B1(data_out_8[1]), .B2(n47), 
        .ZN(n132) );
  AOI22_X1 U137 ( .A1(data_out_9[2]), .A2(n46), .B1(data_out_8[2]), .B2(n47), 
        .ZN(n121) );
  AOI22_X1 U138 ( .A1(data_out_9[3]), .A2(n46), .B1(data_out_8[3]), .B2(n47), 
        .ZN(n110) );
  AOI22_X1 U139 ( .A1(data_out_9[4]), .A2(n46), .B1(data_out_8[4]), .B2(n47), 
        .ZN(n99) );
  AOI22_X1 U140 ( .A1(data_out_9[5]), .A2(n46), .B1(data_out_8[5]), .B2(n47), 
        .ZN(n88) );
  AOI22_X1 U141 ( .A1(data_out_9[6]), .A2(n46), .B1(data_out_8[6]), .B2(n47), 
        .ZN(n77) );
  AOI22_X1 U142 ( .A1(data_out_9[7]), .A2(n46), .B1(data_out_8[7]), .B2(n47), 
        .ZN(n66) );
  AOI22_X1 U143 ( .A1(data_out_9[8]), .A2(n46), .B1(data_out_8[8]), .B2(n47), 
        .ZN(n55) );
  AOI22_X1 U144 ( .A1(data_out_9[9]), .A2(n46), .B1(data_out_8[9]), .B2(n47), 
        .ZN(n36) );
  AOI22_X1 U145 ( .A1(data_out_9[10]), .A2(n46), .B1(data_out_8[10]), .B2(n47), 
        .ZN(n198) );
  AOI22_X1 U146 ( .A1(data_out_9[11]), .A2(n46), .B1(data_out_8[11]), .B2(n47), 
        .ZN(n187) );
  AOI22_X1 U147 ( .A1(data_out_9[12]), .A2(n46), .B1(data_out_8[12]), .B2(n47), 
        .ZN(n176) );
  AOI22_X1 U148 ( .A1(data_out_9[13]), .A2(n46), .B1(data_out_8[13]), .B2(n47), 
        .ZN(n165) );
  AOI22_X1 U149 ( .A1(data_out_9[14]), .A2(n46), .B1(data_out_8[14]), .B2(n47), 
        .ZN(n154) );
  AOI22_X1 U150 ( .A1(data_out_9[15]), .A2(n46), .B1(data_out_8[15]), .B2(n47), 
        .ZN(n143) );
  AND2_X1 U151 ( .A1(sel[2]), .A2(sel[1]), .ZN(n210) );
  AND2_X1 U152 ( .A1(sel[2]), .A2(n275), .ZN(n212) );
  INV_X1 U153 ( .A(sel[3]), .ZN(n276) );
  INV_X1 U154 ( .A(sel[1]), .ZN(n275) );
  NAND4_X1 U155 ( .A1(n205), .A2(n206), .A3(n207), .A4(n208), .ZN(n204) );
  AOI22_X1 U156 ( .A1(data_out_1[0]), .A2(n34), .B1(data_out_0[0]), .B2(n35), 
        .ZN(n205) );
  AOI22_X1 U157 ( .A1(data_out_7[0]), .A2(n28), .B1(data_out_6[0]), .B2(n29), 
        .ZN(n208) );
  AOI22_X1 U158 ( .A1(data_out_3[0]), .A2(n32), .B1(data_out_2[0]), .B2(n33), 
        .ZN(n206) );
  NAND4_X1 U159 ( .A1(n128), .A2(n129), .A3(n130), .A4(n131), .ZN(n127) );
  AOI22_X1 U160 ( .A1(data_out_1[1]), .A2(n34), .B1(data_out_0[1]), .B2(n35), 
        .ZN(n128) );
  AOI22_X1 U161 ( .A1(data_out_7[1]), .A2(n28), .B1(data_out_6[1]), .B2(n29), 
        .ZN(n131) );
  AOI22_X1 U162 ( .A1(data_out_3[1]), .A2(n32), .B1(data_out_2[1]), .B2(n33), 
        .ZN(n129) );
  NAND4_X1 U163 ( .A1(n117), .A2(n118), .A3(n119), .A4(n120), .ZN(n116) );
  AOI22_X1 U164 ( .A1(data_out_1[2]), .A2(n34), .B1(data_out_0[2]), .B2(n35), 
        .ZN(n117) );
  AOI22_X1 U165 ( .A1(data_out_7[2]), .A2(n28), .B1(data_out_6[2]), .B2(n29), 
        .ZN(n120) );
  AOI22_X1 U166 ( .A1(data_out_3[2]), .A2(n32), .B1(data_out_2[2]), .B2(n33), 
        .ZN(n118) );
  NAND4_X1 U167 ( .A1(n106), .A2(n107), .A3(n108), .A4(n109), .ZN(n105) );
  AOI22_X1 U168 ( .A1(data_out_1[3]), .A2(n34), .B1(data_out_0[3]), .B2(n35), 
        .ZN(n106) );
  AOI22_X1 U169 ( .A1(data_out_7[3]), .A2(n28), .B1(data_out_6[3]), .B2(n29), 
        .ZN(n109) );
  AOI22_X1 U170 ( .A1(data_out_3[3]), .A2(n32), .B1(data_out_2[3]), .B2(n33), 
        .ZN(n107) );
  NAND4_X1 U171 ( .A1(n95), .A2(n96), .A3(n97), .A4(n98), .ZN(n94) );
  AOI22_X1 U172 ( .A1(data_out_1[4]), .A2(n34), .B1(data_out_0[4]), .B2(n35), 
        .ZN(n95) );
  AOI22_X1 U173 ( .A1(data_out_7[4]), .A2(n28), .B1(data_out_6[4]), .B2(n29), 
        .ZN(n98) );
  AOI22_X1 U174 ( .A1(data_out_3[4]), .A2(n32), .B1(data_out_2[4]), .B2(n33), 
        .ZN(n96) );
  NAND4_X1 U175 ( .A1(n84), .A2(n85), .A3(n86), .A4(n87), .ZN(n83) );
  AOI22_X1 U176 ( .A1(data_out_1[5]), .A2(n34), .B1(data_out_0[5]), .B2(n35), 
        .ZN(n84) );
  AOI22_X1 U177 ( .A1(data_out_7[5]), .A2(n28), .B1(data_out_6[5]), .B2(n29), 
        .ZN(n87) );
  AOI22_X1 U178 ( .A1(data_out_3[5]), .A2(n32), .B1(data_out_2[5]), .B2(n33), 
        .ZN(n85) );
  NAND4_X1 U179 ( .A1(n73), .A2(n74), .A3(n75), .A4(n76), .ZN(n72) );
  AOI22_X1 U180 ( .A1(data_out_1[6]), .A2(n34), .B1(data_out_0[6]), .B2(n35), 
        .ZN(n73) );
  AOI22_X1 U181 ( .A1(data_out_7[6]), .A2(n28), .B1(data_out_6[6]), .B2(n29), 
        .ZN(n76) );
  AOI22_X1 U182 ( .A1(data_out_3[6]), .A2(n32), .B1(data_out_2[6]), .B2(n33), 
        .ZN(n74) );
  NAND4_X1 U183 ( .A1(n62), .A2(n63), .A3(n64), .A4(n65), .ZN(n61) );
  AOI22_X1 U184 ( .A1(data_out_1[7]), .A2(n34), .B1(data_out_0[7]), .B2(n35), 
        .ZN(n62) );
  AOI22_X1 U185 ( .A1(data_out_7[7]), .A2(n28), .B1(data_out_6[7]), .B2(n29), 
        .ZN(n65) );
  AOI22_X1 U186 ( .A1(data_out_3[7]), .A2(n32), .B1(data_out_2[7]), .B2(n33), 
        .ZN(n63) );
  NAND4_X1 U187 ( .A1(n51), .A2(n52), .A3(n53), .A4(n54), .ZN(n50) );
  AOI22_X1 U188 ( .A1(data_out_1[8]), .A2(n34), .B1(data_out_0[8]), .B2(n35), 
        .ZN(n51) );
  AOI22_X1 U189 ( .A1(data_out_7[8]), .A2(n28), .B1(data_out_6[8]), .B2(n29), 
        .ZN(n54) );
  AOI22_X1 U190 ( .A1(data_out_3[8]), .A2(n32), .B1(data_out_2[8]), .B2(n33), 
        .ZN(n52) );
  NAND4_X1 U191 ( .A1(n24), .A2(n25), .A3(n26), .A4(n27), .ZN(n23) );
  AOI22_X1 U192 ( .A1(data_out_1[9]), .A2(n34), .B1(data_out_0[9]), .B2(n35), 
        .ZN(n24) );
  AOI22_X1 U193 ( .A1(data_out_7[9]), .A2(n28), .B1(data_out_6[9]), .B2(n29), 
        .ZN(n27) );
  AOI22_X1 U194 ( .A1(data_out_3[9]), .A2(n32), .B1(data_out_2[9]), .B2(n33), 
        .ZN(n25) );
  NAND4_X1 U195 ( .A1(n194), .A2(n195), .A3(n196), .A4(n197), .ZN(n193) );
  AOI22_X1 U196 ( .A1(data_out_1[10]), .A2(n34), .B1(data_out_0[10]), .B2(n35), 
        .ZN(n194) );
  AOI22_X1 U197 ( .A1(data_out_7[10]), .A2(n28), .B1(data_out_6[10]), .B2(n29), 
        .ZN(n197) );
  AOI22_X1 U198 ( .A1(data_out_3[10]), .A2(n32), .B1(data_out_2[10]), .B2(n33), 
        .ZN(n195) );
  NAND4_X1 U199 ( .A1(n183), .A2(n184), .A3(n185), .A4(n186), .ZN(n182) );
  AOI22_X1 U200 ( .A1(data_out_1[11]), .A2(n34), .B1(data_out_0[11]), .B2(n35), 
        .ZN(n183) );
  AOI22_X1 U201 ( .A1(data_out_7[11]), .A2(n28), .B1(data_out_6[11]), .B2(n29), 
        .ZN(n186) );
  AOI22_X1 U202 ( .A1(data_out_3[11]), .A2(n32), .B1(data_out_2[11]), .B2(n33), 
        .ZN(n184) );
  NAND4_X1 U203 ( .A1(n172), .A2(n173), .A3(n174), .A4(n175), .ZN(n171) );
  AOI22_X1 U204 ( .A1(data_out_1[12]), .A2(n34), .B1(data_out_0[12]), .B2(n35), 
        .ZN(n172) );
  AOI22_X1 U205 ( .A1(data_out_7[12]), .A2(n28), .B1(data_out_6[12]), .B2(n29), 
        .ZN(n175) );
  AOI22_X1 U206 ( .A1(data_out_3[12]), .A2(n32), .B1(data_out_2[12]), .B2(n33), 
        .ZN(n173) );
  NAND4_X1 U207 ( .A1(n161), .A2(n162), .A3(n163), .A4(n164), .ZN(n160) );
  AOI22_X1 U208 ( .A1(data_out_1[13]), .A2(n34), .B1(data_out_0[13]), .B2(n35), 
        .ZN(n161) );
  AOI22_X1 U209 ( .A1(data_out_7[13]), .A2(n28), .B1(data_out_6[13]), .B2(n29), 
        .ZN(n164) );
  AOI22_X1 U210 ( .A1(data_out_3[13]), .A2(n32), .B1(data_out_2[13]), .B2(n33), 
        .ZN(n162) );
  NAND4_X1 U211 ( .A1(n150), .A2(n151), .A3(n152), .A4(n153), .ZN(n149) );
  AOI22_X1 U212 ( .A1(data_out_1[14]), .A2(n34), .B1(data_out_0[14]), .B2(n35), 
        .ZN(n150) );
  AOI22_X1 U213 ( .A1(data_out_7[14]), .A2(n28), .B1(data_out_6[14]), .B2(n29), 
        .ZN(n153) );
  AOI22_X1 U214 ( .A1(data_out_3[14]), .A2(n32), .B1(data_out_2[14]), .B2(n33), 
        .ZN(n151) );
  NAND4_X1 U215 ( .A1(n139), .A2(n140), .A3(n141), .A4(n142), .ZN(n138) );
  AOI22_X1 U216 ( .A1(data_out_1[15]), .A2(n34), .B1(data_out_0[15]), .B2(n35), 
        .ZN(n139) );
  AOI22_X1 U217 ( .A1(data_out_7[15]), .A2(n28), .B1(data_out_6[15]), .B2(n29), 
        .ZN(n142) );
  AOI22_X1 U218 ( .A1(data_out_3[15]), .A2(n32), .B1(data_out_2[15]), .B2(n33), 
        .ZN(n140) );
  BUF_X1 U219 ( .A(clear_acc), .Z(n225) );
  INV_X1 U220 ( .A(sel[0]), .ZN(n273) );
  OAI21_X1 U221 ( .B1(n274), .B2(n271), .A(n125), .ZN(data_out[1]) );
  INV_X1 U222 ( .A(data_out_15[1]), .ZN(n271) );
  OAI21_X1 U223 ( .B1(n126), .B2(n127), .A(n223), .ZN(n125) );
  NAND4_X1 U224 ( .A1(n132), .A2(n133), .A3(n134), .A4(n135), .ZN(n126) );
  OAI21_X1 U225 ( .B1(n274), .B2(n262), .A(n191), .ZN(data_out[10]) );
  INV_X1 U226 ( .A(data_out_15[10]), .ZN(n262) );
  OAI21_X1 U227 ( .B1(n192), .B2(n193), .A(n274), .ZN(n191) );
  NAND4_X1 U228 ( .A1(n198), .A2(n199), .A3(n200), .A4(n201), .ZN(n192) );
  OAI21_X1 U229 ( .B1(n223), .B2(n261), .A(n180), .ZN(data_out[11]) );
  INV_X1 U230 ( .A(data_out_15[11]), .ZN(n261) );
  OAI21_X1 U231 ( .B1(n181), .B2(n182), .A(n274), .ZN(n180) );
  NAND4_X1 U232 ( .A1(n187), .A2(n188), .A3(n189), .A4(n190), .ZN(n181) );
  OAI21_X1 U233 ( .B1(n274), .B2(n260), .A(n169), .ZN(data_out[12]) );
  INV_X1 U234 ( .A(data_out_15[12]), .ZN(n260) );
  OAI21_X1 U235 ( .B1(n170), .B2(n171), .A(n274), .ZN(n169) );
  NAND4_X1 U236 ( .A1(n176), .A2(n177), .A3(n178), .A4(n179), .ZN(n170) );
  OAI21_X1 U237 ( .B1(n223), .B2(n259), .A(n158), .ZN(data_out[13]) );
  INV_X1 U238 ( .A(data_out_15[13]), .ZN(n259) );
  OAI21_X1 U239 ( .B1(n159), .B2(n160), .A(n274), .ZN(n158) );
  NAND4_X1 U240 ( .A1(n165), .A2(n166), .A3(n167), .A4(n168), .ZN(n159) );
  OAI21_X1 U241 ( .B1(n274), .B2(n258), .A(n147), .ZN(data_out[14]) );
  INV_X1 U242 ( .A(data_out_15[14]), .ZN(n258) );
  OAI21_X1 U243 ( .B1(n148), .B2(n149), .A(n274), .ZN(n147) );
  NAND4_X1 U244 ( .A1(n154), .A2(n155), .A3(n156), .A4(n157), .ZN(n148) );
  OAI21_X1 U245 ( .B1(n274), .B2(n257), .A(n136), .ZN(data_out[15]) );
  INV_X1 U246 ( .A(data_out_15[15]), .ZN(n257) );
  OAI21_X1 U247 ( .B1(n137), .B2(n138), .A(n274), .ZN(n136) );
  NAND4_X1 U248 ( .A1(n143), .A2(n144), .A3(n145), .A4(n146), .ZN(n137) );
  OAI21_X1 U249 ( .B1(n223), .B2(n272), .A(n202), .ZN(data_out[0]) );
  INV_X1 U250 ( .A(data_out_15[0]), .ZN(n272) );
  OAI21_X1 U251 ( .B1(n203), .B2(n204), .A(n274), .ZN(n202) );
  NAND4_X1 U252 ( .A1(n215), .A2(n216), .A3(n217), .A4(n218), .ZN(n203) );
  OAI21_X1 U253 ( .B1(n223), .B2(n270), .A(n114), .ZN(data_out[2]) );
  INV_X1 U254 ( .A(data_out_15[2]), .ZN(n270) );
  OAI21_X1 U255 ( .B1(n115), .B2(n116), .A(n223), .ZN(n114) );
  NAND4_X1 U256 ( .A1(n121), .A2(n122), .A3(n123), .A4(n124), .ZN(n115) );
  OAI21_X1 U257 ( .B1(n223), .B2(n269), .A(n103), .ZN(data_out[3]) );
  INV_X1 U258 ( .A(data_out_15[3]), .ZN(n269) );
  OAI21_X1 U259 ( .B1(n104), .B2(n105), .A(n223), .ZN(n103) );
  NAND4_X1 U260 ( .A1(n110), .A2(n111), .A3(n112), .A4(n113), .ZN(n104) );
  OAI21_X1 U261 ( .B1(n223), .B2(n268), .A(n92), .ZN(data_out[4]) );
  INV_X1 U262 ( .A(data_out_15[4]), .ZN(n268) );
  OAI21_X1 U263 ( .B1(n93), .B2(n94), .A(n223), .ZN(n92) );
  NAND4_X1 U264 ( .A1(n99), .A2(n100), .A3(n101), .A4(n102), .ZN(n93) );
  OAI21_X1 U265 ( .B1(n223), .B2(n267), .A(n81), .ZN(data_out[5]) );
  INV_X1 U266 ( .A(data_out_15[5]), .ZN(n267) );
  OAI21_X1 U267 ( .B1(n82), .B2(n83), .A(n223), .ZN(n81) );
  NAND4_X1 U268 ( .A1(n88), .A2(n89), .A3(n90), .A4(n91), .ZN(n82) );
  OAI21_X1 U269 ( .B1(n223), .B2(n266), .A(n70), .ZN(data_out[6]) );
  INV_X1 U270 ( .A(data_out_15[6]), .ZN(n266) );
  OAI21_X1 U271 ( .B1(n71), .B2(n72), .A(n223), .ZN(n70) );
  NAND4_X1 U272 ( .A1(n77), .A2(n78), .A3(n79), .A4(n80), .ZN(n71) );
  OAI21_X1 U273 ( .B1(n223), .B2(n265), .A(n59), .ZN(data_out[7]) );
  INV_X1 U274 ( .A(data_out_15[7]), .ZN(n265) );
  OAI21_X1 U275 ( .B1(n60), .B2(n61), .A(n274), .ZN(n59) );
  NAND4_X1 U276 ( .A1(n66), .A2(n67), .A3(n68), .A4(n69), .ZN(n60) );
  OAI21_X1 U277 ( .B1(n223), .B2(n264), .A(n48), .ZN(data_out[8]) );
  INV_X1 U278 ( .A(data_out_15[8]), .ZN(n264) );
  OAI21_X1 U279 ( .B1(n49), .B2(n50), .A(n274), .ZN(n48) );
  NAND4_X1 U280 ( .A1(n55), .A2(n56), .A3(n57), .A4(n58), .ZN(n49) );
  OAI21_X1 U281 ( .B1(n263), .B2(n274), .A(n21), .ZN(data_out[9]) );
  INV_X1 U282 ( .A(data_out_15[9]), .ZN(n263) );
  OAI21_X1 U283 ( .B1(n22), .B2(n23), .A(n274), .ZN(n21) );
  NAND4_X1 U284 ( .A1(n36), .A2(n37), .A3(n38), .A4(n39), .ZN(n22) );
  BUF_X1 U285 ( .A(data_out_x[11]), .Z(n249) );
  BUF_X1 U286 ( .A(data_out_x[13]), .Z(n253) );
  BUF_X1 U287 ( .A(data_out_x[15]), .Z(n256) );
  BUF_X2 U288 ( .A(data_out_x[5]), .Z(n237) );
  CLKBUF_X1 U289 ( .A(wr_en_y), .Z(n224) );
  CLKBUF_X3 U290 ( .A(data_out_x[9]), .Z(n245) );
  CLKBUF_X3 U291 ( .A(data_out_x[11]), .Z(n248) );
  CLKBUF_X3 U292 ( .A(data_out_x[13]), .Z(n252) );
endmodule


module network_4_8_12_16_36_16 ( clk, reset, s_valid, m_ready, data_in, 
        m_valid, s_ready, data_out );
  input [15:0] data_in;
  output [15:0] data_out;
  input clk, reset, s_valid, m_ready;
  output m_valid, s_ready;
  wire   ready_1, valid_1, ready_2, valid_2;
  wire   [15:0] data_1;
  wire   [15:0] data_2;

  layer1_8_4_8_16 layer1 ( .clk(clk), .reset(reset), .s_valid(s_valid), 
        .m_ready(ready_1), .data_in(data_in), .m_valid(valid_1), .s_ready(
        s_ready), .data_out(data_1) );
  layer2_12_8_12_16 layer2 ( .clk(clk), .reset(reset), .s_valid(valid_1), 
        .m_ready(ready_2), .data_in(data_1), .m_valid(valid_2), .s_ready(
        ready_1), .data_out(data_2) );
  layer3_16_12_16_16 layer3 ( .clk(clk), .reset(reset), .s_valid(valid_2), 
        .m_ready(m_ready), .data_in(data_2), .m_valid(m_valid), .s_ready(
        ready_2), .data_out(data_out) );
endmodule

