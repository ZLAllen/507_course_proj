
module memory_WIDTH32_SIZE16_LOGSIZE5 ( clk, data_in, data_out, addr, wr_en );
  input [31:0] data_in;
  output [31:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, \mem[15][31] , \mem[15][30] , \mem[15][29] ,
         \mem[15][28] , \mem[15][27] , \mem[15][26] , \mem[15][25] ,
         \mem[15][24] , \mem[15][23] , \mem[15][22] , \mem[15][21] ,
         \mem[15][20] , \mem[15][19] , \mem[15][18] , \mem[15][17] ,
         \mem[15][16] , \mem[15][15] , \mem[15][14] , \mem[15][13] ,
         \mem[15][12] , \mem[15][11] , \mem[15][10] , \mem[15][9] ,
         \mem[15][8] , \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] ,
         \mem[15][3] , \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][31] ,
         \mem[14][30] , \mem[14][29] , \mem[14][28] , \mem[14][27] ,
         \mem[14][26] , \mem[14][25] , \mem[14][24] , \mem[14][23] ,
         \mem[14][22] , \mem[14][21] , \mem[14][20] , \mem[14][19] ,
         \mem[14][18] , \mem[14][17] , \mem[14][16] , \mem[14][15] ,
         \mem[14][14] , \mem[14][13] , \mem[14][12] , \mem[14][11] ,
         \mem[14][10] , \mem[14][9] , \mem[14][8] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][31] , \mem[13][30] , \mem[13][29] ,
         \mem[13][28] , \mem[13][27] , \mem[13][26] , \mem[13][25] ,
         \mem[13][24] , \mem[13][23] , \mem[13][22] , \mem[13][21] ,
         \mem[13][20] , \mem[13][19] , \mem[13][18] , \mem[13][17] ,
         \mem[13][16] , \mem[13][15] , \mem[13][14] , \mem[13][13] ,
         \mem[13][12] , \mem[13][11] , \mem[13][10] , \mem[13][9] ,
         \mem[13][8] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][31] ,
         \mem[12][30] , \mem[12][29] , \mem[12][28] , \mem[12][27] ,
         \mem[12][26] , \mem[12][25] , \mem[12][24] , \mem[12][23] ,
         \mem[12][22] , \mem[12][21] , \mem[12][20] , \mem[12][19] ,
         \mem[12][18] , \mem[12][17] , \mem[12][16] , \mem[12][15] ,
         \mem[12][14] , \mem[12][13] , \mem[12][12] , \mem[12][11] ,
         \mem[12][10] , \mem[12][9] , \mem[12][8] , \mem[12][7] , \mem[12][6] ,
         \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] , \mem[12][1] ,
         \mem[12][0] , \mem[11][31] , \mem[11][30] , \mem[11][29] ,
         \mem[11][28] , \mem[11][27] , \mem[11][26] , \mem[11][25] ,
         \mem[11][24] , \mem[11][23] , \mem[11][22] , \mem[11][21] ,
         \mem[11][20] , \mem[11][19] , \mem[11][18] , \mem[11][17] ,
         \mem[11][16] , \mem[11][15] , \mem[11][14] , \mem[11][13] ,
         \mem[11][12] , \mem[11][11] , \mem[11][10] , \mem[11][9] ,
         \mem[11][8] , \mem[11][7] , \mem[11][6] , \mem[11][5] , \mem[11][4] ,
         \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] , \mem[10][31] ,
         \mem[10][30] , \mem[10][29] , \mem[10][28] , \mem[10][27] ,
         \mem[10][26] , \mem[10][25] , \mem[10][24] , \mem[10][23] ,
         \mem[10][22] , \mem[10][21] , \mem[10][20] , \mem[10][19] ,
         \mem[10][18] , \mem[10][17] , \mem[10][16] , \mem[10][15] ,
         \mem[10][14] , \mem[10][13] , \mem[10][12] , \mem[10][11] ,
         \mem[10][10] , \mem[10][9] , \mem[10][8] , \mem[10][7] , \mem[10][6] ,
         \mem[10][5] , \mem[10][4] , \mem[10][3] , \mem[10][2] , \mem[10][1] ,
         \mem[10][0] , \mem[9][31] , \mem[9][30] , \mem[9][29] , \mem[9][28] ,
         \mem[9][27] , \mem[9][26] , \mem[9][25] , \mem[9][24] , \mem[9][23] ,
         \mem[9][22] , \mem[9][21] , \mem[9][20] , \mem[9][19] , \mem[9][18] ,
         \mem[9][17] , \mem[9][16] , \mem[9][15] , \mem[9][14] , \mem[9][13] ,
         \mem[9][12] , \mem[9][11] , \mem[9][10] , \mem[9][9] , \mem[9][8] ,
         \mem[9][7] , \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] ,
         \mem[9][2] , \mem[9][1] , \mem[9][0] , \mem[8][31] , \mem[8][30] ,
         \mem[8][29] , \mem[8][28] , \mem[8][27] , \mem[8][26] , \mem[8][25] ,
         \mem[8][24] , \mem[8][23] , \mem[8][22] , \mem[8][21] , \mem[8][20] ,
         \mem[8][19] , \mem[8][18] , \mem[8][17] , \mem[8][16] , \mem[8][15] ,
         \mem[8][14] , \mem[8][13] , \mem[8][12] , \mem[8][11] , \mem[8][10] ,
         \mem[8][9] , \mem[8][8] , \mem[8][7] , \mem[8][6] , \mem[8][5] ,
         \mem[8][4] , \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] ,
         \mem[7][31] , \mem[7][30] , \mem[7][29] , \mem[7][28] , \mem[7][27] ,
         \mem[7][26] , \mem[7][25] , \mem[7][24] , \mem[7][23] , \mem[7][22] ,
         \mem[7][21] , \mem[7][20] , \mem[7][19] , \mem[7][18] , \mem[7][17] ,
         \mem[7][16] , \mem[7][15] , \mem[7][14] , \mem[7][13] , \mem[7][12] ,
         \mem[7][11] , \mem[7][10] , \mem[7][9] , \mem[7][8] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][31] , \mem[6][30] , \mem[6][29] ,
         \mem[6][28] , \mem[6][27] , \mem[6][26] , \mem[6][25] , \mem[6][24] ,
         \mem[6][23] , \mem[6][22] , \mem[6][21] , \mem[6][20] , \mem[6][19] ,
         \mem[6][18] , \mem[6][17] , \mem[6][16] , \mem[6][15] , \mem[6][14] ,
         \mem[6][13] , \mem[6][12] , \mem[6][11] , \mem[6][10] , \mem[6][9] ,
         \mem[6][8] , \mem[6][7] , \mem[6][6] , \mem[6][5] , \mem[6][4] ,
         \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] , \mem[5][31] ,
         \mem[5][30] , \mem[5][29] , \mem[5][28] , \mem[5][27] , \mem[5][26] ,
         \mem[5][25] , \mem[5][24] , \mem[5][23] , \mem[5][22] , \mem[5][21] ,
         \mem[5][20] , \mem[5][19] , \mem[5][18] , \mem[5][17] , \mem[5][16] ,
         \mem[5][15] , \mem[5][14] , \mem[5][13] , \mem[5][12] , \mem[5][11] ,
         \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[4][31] , \mem[4][30] , \mem[4][29] , \mem[4][28] ,
         \mem[4][27] , \mem[4][26] , \mem[4][25] , \mem[4][24] , \mem[4][23] ,
         \mem[4][22] , \mem[4][21] , \mem[4][20] , \mem[4][19] , \mem[4][18] ,
         \mem[4][17] , \mem[4][16] , \mem[4][15] , \mem[4][14] , \mem[4][13] ,
         \mem[4][12] , \mem[4][11] , \mem[4][10] , \mem[4][9] , \mem[4][8] ,
         \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] ,
         \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[3][31] , \mem[3][30] ,
         \mem[3][29] , \mem[3][28] , \mem[3][27] , \mem[3][26] , \mem[3][25] ,
         \mem[3][24] , \mem[3][23] , \mem[3][22] , \mem[3][21] , \mem[3][20] ,
         \mem[3][19] , \mem[3][18] , \mem[3][17] , \mem[3][16] , \mem[3][15] ,
         \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] , \mem[3][10] ,
         \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] , \mem[3][5] ,
         \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] ,
         \mem[2][31] , \mem[2][30] , \mem[2][29] , \mem[2][28] , \mem[2][27] ,
         \mem[2][26] , \mem[2][25] , \mem[2][24] , \mem[2][23] , \mem[2][22] ,
         \mem[2][21] , \mem[2][20] , \mem[2][19] , \mem[2][18] , \mem[2][17] ,
         \mem[2][16] , \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] ,
         \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][31] , \mem[1][30] , \mem[1][29] ,
         \mem[1][28] , \mem[1][27] , \mem[1][26] , \mem[1][25] , \mem[1][24] ,
         \mem[1][23] , \mem[1][22] , \mem[1][21] , \mem[1][20] , \mem[1][19] ,
         \mem[1][18] , \mem[1][17] , \mem[1][16] , \mem[1][15] , \mem[1][14] ,
         \mem[1][13] , \mem[1][12] , \mem[1][11] , \mem[1][10] , \mem[1][9] ,
         \mem[1][8] , \mem[1][7] , \mem[1][6] , \mem[1][5] , \mem[1][4] ,
         \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] , \mem[0][31] ,
         \mem[0][30] , \mem[0][29] , \mem[0][28] , \mem[0][27] , \mem[0][26] ,
         \mem[0][25] , \mem[0][24] , \mem[0][23] , \mem[0][22] , \mem[0][21] ,
         \mem[0][20] , \mem[0][19] , \mem[0][18] , \mem[0][17] , \mem[0][16] ,
         \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , N14, N16, N17, N19, N21, N25, N29, N37, N39, N43, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];

  DFF_X1 \data_out_reg[31]  ( .D(N14), .CK(clk), .Q(data_out[31]) );
  DFF_X1 \data_out_reg[29]  ( .D(N16), .CK(clk), .QN(n1) );
  DFF_X1 \data_out_reg[28]  ( .D(N17), .CK(clk), .Q(data_out[28]) );
  DFF_X1 \data_out_reg[26]  ( .D(N19), .CK(clk), .Q(data_out[26]) );
  DFF_X1 \data_out_reg[24]  ( .D(N21), .CK(clk), .Q(data_out[24]) );
  DFF_X1 \data_out_reg[20]  ( .D(N25), .CK(clk), .Q(data_out[20]) );
  DFF_X1 \data_out_reg[16]  ( .D(N29), .CK(clk), .Q(data_out[16]) );
  DFF_X1 \data_out_reg[8]  ( .D(N37), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[6]  ( .D(N39), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[2]  ( .D(N43), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[15][31]  ( .D(n1087), .CK(clk), .Q(\mem[15][31] ) );
  DFF_X1 \mem_reg[15][30]  ( .D(n1086), .CK(clk), .Q(\mem[15][30] ) );
  DFF_X1 \mem_reg[15][29]  ( .D(n1085), .CK(clk), .Q(\mem[15][29] ) );
  DFF_X1 \mem_reg[15][28]  ( .D(n1084), .CK(clk), .Q(\mem[15][28] ) );
  DFF_X1 \mem_reg[15][27]  ( .D(n1083), .CK(clk), .Q(\mem[15][27] ) );
  DFF_X1 \mem_reg[15][26]  ( .D(n1082), .CK(clk), .Q(\mem[15][26] ) );
  DFF_X1 \mem_reg[15][25]  ( .D(n1081), .CK(clk), .Q(\mem[15][25] ) );
  DFF_X1 \mem_reg[15][24]  ( .D(n1080), .CK(clk), .Q(\mem[15][24] ) );
  DFF_X1 \mem_reg[15][23]  ( .D(n1079), .CK(clk), .Q(\mem[15][23] ) );
  DFF_X1 \mem_reg[15][22]  ( .D(n1078), .CK(clk), .Q(\mem[15][22] ) );
  DFF_X1 \mem_reg[15][21]  ( .D(n1077), .CK(clk), .Q(\mem[15][21] ) );
  DFF_X1 \mem_reg[15][20]  ( .D(n1076), .CK(clk), .Q(\mem[15][20] ) );
  DFF_X1 \mem_reg[15][19]  ( .D(n1075), .CK(clk), .Q(\mem[15][19] ) );
  DFF_X1 \mem_reg[15][18]  ( .D(n1074), .CK(clk), .Q(\mem[15][18] ) );
  DFF_X1 \mem_reg[15][17]  ( .D(n1073), .CK(clk), .Q(\mem[15][17] ) );
  DFF_X1 \mem_reg[15][16]  ( .D(n1072), .CK(clk), .Q(\mem[15][16] ) );
  DFF_X1 \mem_reg[15][15]  ( .D(n1071), .CK(clk), .Q(\mem[15][15] ) );
  DFF_X1 \mem_reg[15][14]  ( .D(n1070), .CK(clk), .Q(\mem[15][14] ) );
  DFF_X1 \mem_reg[15][13]  ( .D(n1069), .CK(clk), .Q(\mem[15][13] ) );
  DFF_X1 \mem_reg[15][12]  ( .D(n1068), .CK(clk), .Q(\mem[15][12] ) );
  DFF_X1 \mem_reg[15][11]  ( .D(n1067), .CK(clk), .Q(\mem[15][11] ) );
  DFF_X1 \mem_reg[15][10]  ( .D(n1066), .CK(clk), .Q(\mem[15][10] ) );
  DFF_X1 \mem_reg[15][9]  ( .D(n1065), .CK(clk), .Q(\mem[15][9] ) );
  DFF_X1 \mem_reg[15][8]  ( .D(n1064), .CK(clk), .Q(\mem[15][8] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n1063), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n1062), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n1061), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n1060), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n1059), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n1058), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n1057), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n1056), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][31]  ( .D(n1055), .CK(clk), .Q(\mem[14][31] ) );
  DFF_X1 \mem_reg[14][30]  ( .D(n1054), .CK(clk), .Q(\mem[14][30] ) );
  DFF_X1 \mem_reg[14][29]  ( .D(n1053), .CK(clk), .Q(\mem[14][29] ) );
  DFF_X1 \mem_reg[14][28]  ( .D(n1052), .CK(clk), .Q(\mem[14][28] ) );
  DFF_X1 \mem_reg[14][27]  ( .D(n1051), .CK(clk), .Q(\mem[14][27] ) );
  DFF_X1 \mem_reg[14][26]  ( .D(n1050), .CK(clk), .Q(\mem[14][26] ) );
  DFF_X1 \mem_reg[14][25]  ( .D(n1049), .CK(clk), .Q(\mem[14][25] ) );
  DFF_X1 \mem_reg[14][24]  ( .D(n1048), .CK(clk), .Q(\mem[14][24] ) );
  DFF_X1 \mem_reg[14][23]  ( .D(n1047), .CK(clk), .Q(\mem[14][23] ) );
  DFF_X1 \mem_reg[14][22]  ( .D(n1046), .CK(clk), .Q(\mem[14][22] ) );
  DFF_X1 \mem_reg[14][21]  ( .D(n1045), .CK(clk), .Q(\mem[14][21] ) );
  DFF_X1 \mem_reg[14][20]  ( .D(n1044), .CK(clk), .Q(\mem[14][20] ) );
  DFF_X1 \mem_reg[14][19]  ( .D(n1043), .CK(clk), .Q(\mem[14][19] ) );
  DFF_X1 \mem_reg[14][18]  ( .D(n1042), .CK(clk), .Q(\mem[14][18] ) );
  DFF_X1 \mem_reg[14][17]  ( .D(n1041), .CK(clk), .Q(\mem[14][17] ) );
  DFF_X1 \mem_reg[14][16]  ( .D(n1040), .CK(clk), .Q(\mem[14][16] ) );
  DFF_X1 \mem_reg[14][15]  ( .D(n1039), .CK(clk), .Q(\mem[14][15] ) );
  DFF_X1 \mem_reg[14][14]  ( .D(n1038), .CK(clk), .Q(\mem[14][14] ) );
  DFF_X1 \mem_reg[14][13]  ( .D(n1037), .CK(clk), .Q(\mem[14][13] ) );
  DFF_X1 \mem_reg[14][12]  ( .D(n1036), .CK(clk), .Q(\mem[14][12] ) );
  DFF_X1 \mem_reg[14][11]  ( .D(n1035), .CK(clk), .Q(\mem[14][11] ) );
  DFF_X1 \mem_reg[14][10]  ( .D(n1034), .CK(clk), .Q(\mem[14][10] ) );
  DFF_X1 \mem_reg[14][9]  ( .D(n1033), .CK(clk), .Q(\mem[14][9] ) );
  DFF_X1 \mem_reg[14][8]  ( .D(n1032), .CK(clk), .Q(\mem[14][8] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n1031), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n1030), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n1029), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n1028), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n1027), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n1026), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n1025), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n1024), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][31]  ( .D(n1023), .CK(clk), .Q(\mem[13][31] ) );
  DFF_X1 \mem_reg[13][30]  ( .D(n1022), .CK(clk), .Q(\mem[13][30] ) );
  DFF_X1 \mem_reg[13][29]  ( .D(n1021), .CK(clk), .Q(\mem[13][29] ) );
  DFF_X1 \mem_reg[13][28]  ( .D(n1020), .CK(clk), .Q(\mem[13][28] ) );
  DFF_X1 \mem_reg[13][27]  ( .D(n1019), .CK(clk), .Q(\mem[13][27] ) );
  DFF_X1 \mem_reg[13][26]  ( .D(n1018), .CK(clk), .Q(\mem[13][26] ) );
  DFF_X1 \mem_reg[13][25]  ( .D(n1017), .CK(clk), .Q(\mem[13][25] ) );
  DFF_X1 \mem_reg[13][24]  ( .D(n1016), .CK(clk), .Q(\mem[13][24] ) );
  DFF_X1 \mem_reg[13][23]  ( .D(n1015), .CK(clk), .Q(\mem[13][23] ) );
  DFF_X1 \mem_reg[13][22]  ( .D(n1014), .CK(clk), .Q(\mem[13][22] ) );
  DFF_X1 \mem_reg[13][21]  ( .D(n1013), .CK(clk), .Q(\mem[13][21] ) );
  DFF_X1 \mem_reg[13][20]  ( .D(n1012), .CK(clk), .Q(\mem[13][20] ) );
  DFF_X1 \mem_reg[13][19]  ( .D(n1011), .CK(clk), .Q(\mem[13][19] ) );
  DFF_X1 \mem_reg[13][18]  ( .D(n1010), .CK(clk), .Q(\mem[13][18] ) );
  DFF_X1 \mem_reg[13][17]  ( .D(n1009), .CK(clk), .Q(\mem[13][17] ) );
  DFF_X1 \mem_reg[13][16]  ( .D(n1008), .CK(clk), .Q(\mem[13][16] ) );
  DFF_X1 \mem_reg[13][15]  ( .D(n1007), .CK(clk), .Q(\mem[13][15] ) );
  DFF_X1 \mem_reg[13][14]  ( .D(n1006), .CK(clk), .Q(\mem[13][14] ) );
  DFF_X1 \mem_reg[13][13]  ( .D(n1005), .CK(clk), .Q(\mem[13][13] ) );
  DFF_X1 \mem_reg[13][12]  ( .D(n1004), .CK(clk), .Q(\mem[13][12] ) );
  DFF_X1 \mem_reg[13][11]  ( .D(n1003), .CK(clk), .Q(\mem[13][11] ) );
  DFF_X1 \mem_reg[13][10]  ( .D(n1002), .CK(clk), .Q(\mem[13][10] ) );
  DFF_X1 \mem_reg[13][9]  ( .D(n1001), .CK(clk), .Q(\mem[13][9] ) );
  DFF_X1 \mem_reg[13][8]  ( .D(n1000), .CK(clk), .Q(\mem[13][8] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n999), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n998), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n997), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n996), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n995), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n994), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n993), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n992), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][31]  ( .D(n991), .CK(clk), .Q(\mem[12][31] ) );
  DFF_X1 \mem_reg[12][30]  ( .D(n990), .CK(clk), .Q(\mem[12][30] ) );
  DFF_X1 \mem_reg[12][29]  ( .D(n989), .CK(clk), .Q(\mem[12][29] ) );
  DFF_X1 \mem_reg[12][28]  ( .D(n988), .CK(clk), .Q(\mem[12][28] ) );
  DFF_X1 \mem_reg[12][27]  ( .D(n987), .CK(clk), .Q(\mem[12][27] ) );
  DFF_X1 \mem_reg[12][26]  ( .D(n986), .CK(clk), .Q(\mem[12][26] ) );
  DFF_X1 \mem_reg[12][25]  ( .D(n985), .CK(clk), .Q(\mem[12][25] ) );
  DFF_X1 \mem_reg[12][24]  ( .D(n984), .CK(clk), .Q(\mem[12][24] ) );
  DFF_X1 \mem_reg[12][23]  ( .D(n983), .CK(clk), .Q(\mem[12][23] ) );
  DFF_X1 \mem_reg[12][22]  ( .D(n982), .CK(clk), .Q(\mem[12][22] ) );
  DFF_X1 \mem_reg[12][21]  ( .D(n981), .CK(clk), .Q(\mem[12][21] ) );
  DFF_X1 \mem_reg[12][20]  ( .D(n980), .CK(clk), .Q(\mem[12][20] ) );
  DFF_X1 \mem_reg[12][19]  ( .D(n979), .CK(clk), .Q(\mem[12][19] ) );
  DFF_X1 \mem_reg[12][18]  ( .D(n978), .CK(clk), .Q(\mem[12][18] ) );
  DFF_X1 \mem_reg[12][17]  ( .D(n977), .CK(clk), .Q(\mem[12][17] ) );
  DFF_X1 \mem_reg[12][16]  ( .D(n976), .CK(clk), .Q(\mem[12][16] ) );
  DFF_X1 \mem_reg[12][15]  ( .D(n975), .CK(clk), .Q(\mem[12][15] ) );
  DFF_X1 \mem_reg[12][14]  ( .D(n974), .CK(clk), .Q(\mem[12][14] ) );
  DFF_X1 \mem_reg[12][13]  ( .D(n973), .CK(clk), .Q(\mem[12][13] ) );
  DFF_X1 \mem_reg[12][12]  ( .D(n972), .CK(clk), .Q(\mem[12][12] ) );
  DFF_X1 \mem_reg[12][11]  ( .D(n971), .CK(clk), .Q(\mem[12][11] ) );
  DFF_X1 \mem_reg[12][10]  ( .D(n970), .CK(clk), .Q(\mem[12][10] ) );
  DFF_X1 \mem_reg[12][9]  ( .D(n969), .CK(clk), .Q(\mem[12][9] ) );
  DFF_X1 \mem_reg[12][8]  ( .D(n968), .CK(clk), .Q(\mem[12][8] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n967), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n966), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n965), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n964), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n963), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n962), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n961), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n960), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][31]  ( .D(n959), .CK(clk), .Q(\mem[11][31] ) );
  DFF_X1 \mem_reg[11][30]  ( .D(n958), .CK(clk), .Q(\mem[11][30] ) );
  DFF_X1 \mem_reg[11][29]  ( .D(n957), .CK(clk), .Q(\mem[11][29] ) );
  DFF_X1 \mem_reg[11][28]  ( .D(n956), .CK(clk), .Q(\mem[11][28] ) );
  DFF_X1 \mem_reg[11][27]  ( .D(n955), .CK(clk), .Q(\mem[11][27] ) );
  DFF_X1 \mem_reg[11][26]  ( .D(n954), .CK(clk), .Q(\mem[11][26] ) );
  DFF_X1 \mem_reg[11][25]  ( .D(n953), .CK(clk), .Q(\mem[11][25] ) );
  DFF_X1 \mem_reg[11][24]  ( .D(n952), .CK(clk), .Q(\mem[11][24] ) );
  DFF_X1 \mem_reg[11][23]  ( .D(n951), .CK(clk), .Q(\mem[11][23] ) );
  DFF_X1 \mem_reg[11][22]  ( .D(n950), .CK(clk), .Q(\mem[11][22] ) );
  DFF_X1 \mem_reg[11][21]  ( .D(n949), .CK(clk), .Q(\mem[11][21] ) );
  DFF_X1 \mem_reg[11][20]  ( .D(n948), .CK(clk), .Q(\mem[11][20] ) );
  DFF_X1 \mem_reg[11][19]  ( .D(n947), .CK(clk), .Q(\mem[11][19] ) );
  DFF_X1 \mem_reg[11][18]  ( .D(n946), .CK(clk), .Q(\mem[11][18] ) );
  DFF_X1 \mem_reg[11][17]  ( .D(n945), .CK(clk), .Q(\mem[11][17] ) );
  DFF_X1 \mem_reg[11][16]  ( .D(n944), .CK(clk), .Q(\mem[11][16] ) );
  DFF_X1 \mem_reg[11][15]  ( .D(n943), .CK(clk), .Q(\mem[11][15] ) );
  DFF_X1 \mem_reg[11][14]  ( .D(n942), .CK(clk), .Q(\mem[11][14] ) );
  DFF_X1 \mem_reg[11][13]  ( .D(n941), .CK(clk), .Q(\mem[11][13] ) );
  DFF_X1 \mem_reg[11][12]  ( .D(n940), .CK(clk), .Q(\mem[11][12] ) );
  DFF_X1 \mem_reg[11][11]  ( .D(n939), .CK(clk), .Q(\mem[11][11] ) );
  DFF_X1 \mem_reg[11][10]  ( .D(n938), .CK(clk), .Q(\mem[11][10] ) );
  DFF_X1 \mem_reg[11][9]  ( .D(n937), .CK(clk), .Q(\mem[11][9] ) );
  DFF_X1 \mem_reg[11][8]  ( .D(n936), .CK(clk), .Q(\mem[11][8] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n935), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n934), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n933), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n932), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n931), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n930), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n929), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n928), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][31]  ( .D(n927), .CK(clk), .Q(\mem[10][31] ) );
  DFF_X1 \mem_reg[10][30]  ( .D(n926), .CK(clk), .Q(\mem[10][30] ) );
  DFF_X1 \mem_reg[10][29]  ( .D(n925), .CK(clk), .Q(\mem[10][29] ) );
  DFF_X1 \mem_reg[10][28]  ( .D(n924), .CK(clk), .Q(\mem[10][28] ) );
  DFF_X1 \mem_reg[10][27]  ( .D(n923), .CK(clk), .Q(\mem[10][27] ) );
  DFF_X1 \mem_reg[10][26]  ( .D(n922), .CK(clk), .Q(\mem[10][26] ) );
  DFF_X1 \mem_reg[10][25]  ( .D(n921), .CK(clk), .Q(\mem[10][25] ) );
  DFF_X1 \mem_reg[10][24]  ( .D(n920), .CK(clk), .Q(\mem[10][24] ) );
  DFF_X1 \mem_reg[10][23]  ( .D(n919), .CK(clk), .Q(\mem[10][23] ) );
  DFF_X1 \mem_reg[10][22]  ( .D(n918), .CK(clk), .Q(\mem[10][22] ) );
  DFF_X1 \mem_reg[10][21]  ( .D(n917), .CK(clk), .Q(\mem[10][21] ) );
  DFF_X1 \mem_reg[10][20]  ( .D(n916), .CK(clk), .Q(\mem[10][20] ) );
  DFF_X1 \mem_reg[10][19]  ( .D(n915), .CK(clk), .Q(\mem[10][19] ) );
  DFF_X1 \mem_reg[10][18]  ( .D(n914), .CK(clk), .Q(\mem[10][18] ) );
  DFF_X1 \mem_reg[10][17]  ( .D(n913), .CK(clk), .Q(\mem[10][17] ) );
  DFF_X1 \mem_reg[10][16]  ( .D(n912), .CK(clk), .Q(\mem[10][16] ) );
  DFF_X1 \mem_reg[10][15]  ( .D(n911), .CK(clk), .Q(\mem[10][15] ) );
  DFF_X1 \mem_reg[10][14]  ( .D(n910), .CK(clk), .Q(\mem[10][14] ) );
  DFF_X1 \mem_reg[10][13]  ( .D(n909), .CK(clk), .Q(\mem[10][13] ) );
  DFF_X1 \mem_reg[10][12]  ( .D(n908), .CK(clk), .Q(\mem[10][12] ) );
  DFF_X1 \mem_reg[10][11]  ( .D(n907), .CK(clk), .Q(\mem[10][11] ) );
  DFF_X1 \mem_reg[10][10]  ( .D(n906), .CK(clk), .Q(\mem[10][10] ) );
  DFF_X1 \mem_reg[10][9]  ( .D(n905), .CK(clk), .Q(\mem[10][9] ) );
  DFF_X1 \mem_reg[10][8]  ( .D(n904), .CK(clk), .Q(\mem[10][8] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n903), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n902), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n901), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n900), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n899), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n898), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n897), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n896), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][31]  ( .D(n895), .CK(clk), .Q(\mem[9][31] ) );
  DFF_X1 \mem_reg[9][30]  ( .D(n894), .CK(clk), .Q(\mem[9][30] ) );
  DFF_X1 \mem_reg[9][29]  ( .D(n893), .CK(clk), .Q(\mem[9][29] ) );
  DFF_X1 \mem_reg[9][28]  ( .D(n892), .CK(clk), .Q(\mem[9][28] ) );
  DFF_X1 \mem_reg[9][27]  ( .D(n891), .CK(clk), .Q(\mem[9][27] ) );
  DFF_X1 \mem_reg[9][26]  ( .D(n890), .CK(clk), .Q(\mem[9][26] ) );
  DFF_X1 \mem_reg[9][25]  ( .D(n889), .CK(clk), .Q(\mem[9][25] ) );
  DFF_X1 \mem_reg[9][24]  ( .D(n888), .CK(clk), .Q(\mem[9][24] ) );
  DFF_X1 \mem_reg[9][23]  ( .D(n887), .CK(clk), .Q(\mem[9][23] ) );
  DFF_X1 \mem_reg[9][22]  ( .D(n886), .CK(clk), .Q(\mem[9][22] ) );
  DFF_X1 \mem_reg[9][21]  ( .D(n885), .CK(clk), .Q(\mem[9][21] ) );
  DFF_X1 \mem_reg[9][20]  ( .D(n884), .CK(clk), .Q(\mem[9][20] ) );
  DFF_X1 \mem_reg[9][19]  ( .D(n883), .CK(clk), .Q(\mem[9][19] ) );
  DFF_X1 \mem_reg[9][18]  ( .D(n882), .CK(clk), .Q(\mem[9][18] ) );
  DFF_X1 \mem_reg[9][17]  ( .D(n881), .CK(clk), .Q(\mem[9][17] ) );
  DFF_X1 \mem_reg[9][16]  ( .D(n880), .CK(clk), .Q(\mem[9][16] ) );
  DFF_X1 \mem_reg[9][15]  ( .D(n879), .CK(clk), .Q(\mem[9][15] ) );
  DFF_X1 \mem_reg[9][14]  ( .D(n878), .CK(clk), .Q(\mem[9][14] ) );
  DFF_X1 \mem_reg[9][13]  ( .D(n877), .CK(clk), .Q(\mem[9][13] ) );
  DFF_X1 \mem_reg[9][12]  ( .D(n876), .CK(clk), .Q(\mem[9][12] ) );
  DFF_X1 \mem_reg[9][11]  ( .D(n875), .CK(clk), .Q(\mem[9][11] ) );
  DFF_X1 \mem_reg[9][10]  ( .D(n874), .CK(clk), .Q(\mem[9][10] ) );
  DFF_X1 \mem_reg[9][9]  ( .D(n873), .CK(clk), .Q(\mem[9][9] ) );
  DFF_X1 \mem_reg[9][8]  ( .D(n872), .CK(clk), .Q(\mem[9][8] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n871), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n870), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n869), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n868), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n867), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n866), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n865), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n864), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][31]  ( .D(n863), .CK(clk), .Q(\mem[8][31] ) );
  DFF_X1 \mem_reg[8][30]  ( .D(n862), .CK(clk), .Q(\mem[8][30] ) );
  DFF_X1 \mem_reg[8][29]  ( .D(n861), .CK(clk), .Q(\mem[8][29] ) );
  DFF_X1 \mem_reg[8][28]  ( .D(n860), .CK(clk), .Q(\mem[8][28] ) );
  DFF_X1 \mem_reg[8][27]  ( .D(n859), .CK(clk), .Q(\mem[8][27] ) );
  DFF_X1 \mem_reg[8][26]  ( .D(n858), .CK(clk), .Q(\mem[8][26] ) );
  DFF_X1 \mem_reg[8][25]  ( .D(n857), .CK(clk), .Q(\mem[8][25] ) );
  DFF_X1 \mem_reg[8][24]  ( .D(n856), .CK(clk), .Q(\mem[8][24] ) );
  DFF_X1 \mem_reg[8][23]  ( .D(n855), .CK(clk), .Q(\mem[8][23] ) );
  DFF_X1 \mem_reg[8][22]  ( .D(n854), .CK(clk), .Q(\mem[8][22] ) );
  DFF_X1 \mem_reg[8][21]  ( .D(n853), .CK(clk), .Q(\mem[8][21] ) );
  DFF_X1 \mem_reg[8][20]  ( .D(n852), .CK(clk), .Q(\mem[8][20] ) );
  DFF_X1 \mem_reg[8][19]  ( .D(n851), .CK(clk), .Q(\mem[8][19] ) );
  DFF_X1 \mem_reg[8][18]  ( .D(n850), .CK(clk), .Q(\mem[8][18] ) );
  DFF_X1 \mem_reg[8][17]  ( .D(n849), .CK(clk), .Q(\mem[8][17] ) );
  DFF_X1 \mem_reg[8][16]  ( .D(n848), .CK(clk), .Q(\mem[8][16] ) );
  DFF_X1 \mem_reg[8][15]  ( .D(n847), .CK(clk), .Q(\mem[8][15] ) );
  DFF_X1 \mem_reg[8][14]  ( .D(n846), .CK(clk), .Q(\mem[8][14] ) );
  DFF_X1 \mem_reg[8][13]  ( .D(n845), .CK(clk), .Q(\mem[8][13] ) );
  DFF_X1 \mem_reg[8][12]  ( .D(n844), .CK(clk), .Q(\mem[8][12] ) );
  DFF_X1 \mem_reg[8][11]  ( .D(n843), .CK(clk), .Q(\mem[8][11] ) );
  DFF_X1 \mem_reg[8][10]  ( .D(n842), .CK(clk), .Q(\mem[8][10] ) );
  DFF_X1 \mem_reg[8][9]  ( .D(n841), .CK(clk), .Q(\mem[8][9] ) );
  DFF_X1 \mem_reg[8][8]  ( .D(n840), .CK(clk), .Q(\mem[8][8] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n839), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n838), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n837), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n836), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n835), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n834), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n833), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n832), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][31]  ( .D(n831), .CK(clk), .Q(\mem[7][31] ) );
  DFF_X1 \mem_reg[7][30]  ( .D(n830), .CK(clk), .Q(\mem[7][30] ) );
  DFF_X1 \mem_reg[7][29]  ( .D(n829), .CK(clk), .Q(\mem[7][29] ) );
  DFF_X1 \mem_reg[7][28]  ( .D(n828), .CK(clk), .Q(\mem[7][28] ) );
  DFF_X1 \mem_reg[7][27]  ( .D(n827), .CK(clk), .Q(\mem[7][27] ) );
  DFF_X1 \mem_reg[7][26]  ( .D(n826), .CK(clk), .Q(\mem[7][26] ) );
  DFF_X1 \mem_reg[7][25]  ( .D(n825), .CK(clk), .Q(\mem[7][25] ) );
  DFF_X1 \mem_reg[7][24]  ( .D(n824), .CK(clk), .Q(\mem[7][24] ) );
  DFF_X1 \mem_reg[7][23]  ( .D(n823), .CK(clk), .Q(\mem[7][23] ) );
  DFF_X1 \mem_reg[7][22]  ( .D(n822), .CK(clk), .Q(\mem[7][22] ) );
  DFF_X1 \mem_reg[7][21]  ( .D(n821), .CK(clk), .Q(\mem[7][21] ) );
  DFF_X1 \mem_reg[7][20]  ( .D(n820), .CK(clk), .Q(\mem[7][20] ) );
  DFF_X1 \mem_reg[7][19]  ( .D(n819), .CK(clk), .Q(\mem[7][19] ) );
  DFF_X1 \mem_reg[7][18]  ( .D(n818), .CK(clk), .Q(\mem[7][18] ) );
  DFF_X1 \mem_reg[7][17]  ( .D(n817), .CK(clk), .Q(\mem[7][17] ) );
  DFF_X1 \mem_reg[7][16]  ( .D(n816), .CK(clk), .Q(\mem[7][16] ) );
  DFF_X1 \mem_reg[7][15]  ( .D(n815), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n814), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n813), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n812), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n811), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n810), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n809), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n808), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n807), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n806), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n805), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n804), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n803), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n802), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n801), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n800), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][31]  ( .D(n799), .CK(clk), .Q(\mem[6][31] ) );
  DFF_X1 \mem_reg[6][30]  ( .D(n798), .CK(clk), .Q(\mem[6][30] ) );
  DFF_X1 \mem_reg[6][29]  ( .D(n797), .CK(clk), .Q(\mem[6][29] ) );
  DFF_X1 \mem_reg[6][28]  ( .D(n796), .CK(clk), .Q(\mem[6][28] ) );
  DFF_X1 \mem_reg[6][27]  ( .D(n795), .CK(clk), .Q(\mem[6][27] ) );
  DFF_X1 \mem_reg[6][26]  ( .D(n794), .CK(clk), .Q(\mem[6][26] ) );
  DFF_X1 \mem_reg[6][25]  ( .D(n793), .CK(clk), .Q(\mem[6][25] ) );
  DFF_X1 \mem_reg[6][24]  ( .D(n792), .CK(clk), .Q(\mem[6][24] ) );
  DFF_X1 \mem_reg[6][23]  ( .D(n791), .CK(clk), .Q(\mem[6][23] ) );
  DFF_X1 \mem_reg[6][22]  ( .D(n790), .CK(clk), .Q(\mem[6][22] ) );
  DFF_X1 \mem_reg[6][21]  ( .D(n789), .CK(clk), .Q(\mem[6][21] ) );
  DFF_X1 \mem_reg[6][20]  ( .D(n788), .CK(clk), .Q(\mem[6][20] ) );
  DFF_X1 \mem_reg[6][19]  ( .D(n787), .CK(clk), .Q(\mem[6][19] ) );
  DFF_X1 \mem_reg[6][18]  ( .D(n786), .CK(clk), .Q(\mem[6][18] ) );
  DFF_X1 \mem_reg[6][17]  ( .D(n785), .CK(clk), .Q(\mem[6][17] ) );
  DFF_X1 \mem_reg[6][16]  ( .D(n784), .CK(clk), .Q(\mem[6][16] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n781), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n774), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n773), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n772), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n771), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n770), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n769), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n768), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][31]  ( .D(n767), .CK(clk), .Q(\mem[5][31] ) );
  DFF_X1 \mem_reg[5][30]  ( .D(n766), .CK(clk), .Q(\mem[5][30] ) );
  DFF_X1 \mem_reg[5][29]  ( .D(n765), .CK(clk), .Q(\mem[5][29] ) );
  DFF_X1 \mem_reg[5][28]  ( .D(n764), .CK(clk), .Q(\mem[5][28] ) );
  DFF_X1 \mem_reg[5][27]  ( .D(n763), .CK(clk), .Q(\mem[5][27] ) );
  DFF_X1 \mem_reg[5][26]  ( .D(n762), .CK(clk), .Q(\mem[5][26] ) );
  DFF_X1 \mem_reg[5][25]  ( .D(n761), .CK(clk), .Q(\mem[5][25] ) );
  DFF_X1 \mem_reg[5][24]  ( .D(n760), .CK(clk), .Q(\mem[5][24] ) );
  DFF_X1 \mem_reg[5][23]  ( .D(n759), .CK(clk), .Q(\mem[5][23] ) );
  DFF_X1 \mem_reg[5][22]  ( .D(n758), .CK(clk), .Q(\mem[5][22] ) );
  DFF_X1 \mem_reg[5][21]  ( .D(n757), .CK(clk), .Q(\mem[5][21] ) );
  DFF_X1 \mem_reg[5][20]  ( .D(n756), .CK(clk), .Q(\mem[5][20] ) );
  DFF_X1 \mem_reg[5][19]  ( .D(n755), .CK(clk), .Q(\mem[5][19] ) );
  DFF_X1 \mem_reg[5][18]  ( .D(n754), .CK(clk), .Q(\mem[5][18] ) );
  DFF_X1 \mem_reg[5][17]  ( .D(n753), .CK(clk), .Q(\mem[5][17] ) );
  DFF_X1 \mem_reg[5][16]  ( .D(n752), .CK(clk), .Q(\mem[5][16] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n751), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n750), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n749), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n748), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n747), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n746), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n745), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n744), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n743), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n742), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n741), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n740), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n739), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n738), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n737), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n736), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][31]  ( .D(n735), .CK(clk), .Q(\mem[4][31] ) );
  DFF_X1 \mem_reg[4][30]  ( .D(n734), .CK(clk), .Q(\mem[4][30] ) );
  DFF_X1 \mem_reg[4][29]  ( .D(n733), .CK(clk), .Q(\mem[4][29] ) );
  DFF_X1 \mem_reg[4][28]  ( .D(n732), .CK(clk), .Q(\mem[4][28] ) );
  DFF_X1 \mem_reg[4][27]  ( .D(n731), .CK(clk), .Q(\mem[4][27] ) );
  DFF_X1 \mem_reg[4][26]  ( .D(n730), .CK(clk), .Q(\mem[4][26] ) );
  DFF_X1 \mem_reg[4][25]  ( .D(n729), .CK(clk), .Q(\mem[4][25] ) );
  DFF_X1 \mem_reg[4][24]  ( .D(n728), .CK(clk), .Q(\mem[4][24] ) );
  DFF_X1 \mem_reg[4][23]  ( .D(n727), .CK(clk), .Q(\mem[4][23] ) );
  DFF_X1 \mem_reg[4][22]  ( .D(n726), .CK(clk), .Q(\mem[4][22] ) );
  DFF_X1 \mem_reg[4][21]  ( .D(n725), .CK(clk), .Q(\mem[4][21] ) );
  DFF_X1 \mem_reg[4][20]  ( .D(n724), .CK(clk), .Q(\mem[4][20] ) );
  DFF_X1 \mem_reg[4][19]  ( .D(n723), .CK(clk), .Q(\mem[4][19] ) );
  DFF_X1 \mem_reg[4][18]  ( .D(n722), .CK(clk), .Q(\mem[4][18] ) );
  DFF_X1 \mem_reg[4][17]  ( .D(n721), .CK(clk), .Q(\mem[4][17] ) );
  DFF_X1 \mem_reg[4][16]  ( .D(n720), .CK(clk), .Q(\mem[4][16] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n717), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n710), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n709), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n708), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n707), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n706), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n705), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n704), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][31]  ( .D(n703), .CK(clk), .Q(\mem[3][31] ) );
  DFF_X1 \mem_reg[3][30]  ( .D(n702), .CK(clk), .Q(\mem[3][30] ) );
  DFF_X1 \mem_reg[3][29]  ( .D(n701), .CK(clk), .Q(\mem[3][29] ) );
  DFF_X1 \mem_reg[3][28]  ( .D(n700), .CK(clk), .Q(\mem[3][28] ) );
  DFF_X1 \mem_reg[3][27]  ( .D(n699), .CK(clk), .Q(\mem[3][27] ) );
  DFF_X1 \mem_reg[3][26]  ( .D(n698), .CK(clk), .Q(\mem[3][26] ) );
  DFF_X1 \mem_reg[3][25]  ( .D(n697), .CK(clk), .Q(\mem[3][25] ) );
  DFF_X1 \mem_reg[3][24]  ( .D(n696), .CK(clk), .Q(\mem[3][24] ) );
  DFF_X1 \mem_reg[3][23]  ( .D(n695), .CK(clk), .Q(\mem[3][23] ) );
  DFF_X1 \mem_reg[3][22]  ( .D(n694), .CK(clk), .Q(\mem[3][22] ) );
  DFF_X1 \mem_reg[3][21]  ( .D(n693), .CK(clk), .Q(\mem[3][21] ) );
  DFF_X1 \mem_reg[3][20]  ( .D(n692), .CK(clk), .Q(\mem[3][20] ) );
  DFF_X1 \mem_reg[3][19]  ( .D(n691), .CK(clk), .Q(\mem[3][19] ) );
  DFF_X1 \mem_reg[3][18]  ( .D(n690), .CK(clk), .Q(\mem[3][18] ) );
  DFF_X1 \mem_reg[3][17]  ( .D(n689), .CK(clk), .Q(\mem[3][17] ) );
  DFF_X1 \mem_reg[3][16]  ( .D(n688), .CK(clk), .Q(\mem[3][16] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n687), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n686), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n685), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n684), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n683), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n682), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n681), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n680), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n679), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n678), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n677), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n676), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n675), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n674), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n673), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n672), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][31]  ( .D(n671), .CK(clk), .Q(\mem[2][31] ) );
  DFF_X1 \mem_reg[2][30]  ( .D(n670), .CK(clk), .Q(\mem[2][30] ) );
  DFF_X1 \mem_reg[2][29]  ( .D(n669), .CK(clk), .Q(\mem[2][29] ) );
  DFF_X1 \mem_reg[2][28]  ( .D(n668), .CK(clk), .Q(\mem[2][28] ) );
  DFF_X1 \mem_reg[2][27]  ( .D(n667), .CK(clk), .Q(\mem[2][27] ) );
  DFF_X1 \mem_reg[2][26]  ( .D(n666), .CK(clk), .Q(\mem[2][26] ) );
  DFF_X1 \mem_reg[2][25]  ( .D(n665), .CK(clk), .Q(\mem[2][25] ) );
  DFF_X1 \mem_reg[2][24]  ( .D(n664), .CK(clk), .Q(\mem[2][24] ) );
  DFF_X1 \mem_reg[2][23]  ( .D(n663), .CK(clk), .Q(\mem[2][23] ) );
  DFF_X1 \mem_reg[2][22]  ( .D(n662), .CK(clk), .Q(\mem[2][22] ) );
  DFF_X1 \mem_reg[2][21]  ( .D(n661), .CK(clk), .Q(\mem[2][21] ) );
  DFF_X1 \mem_reg[2][20]  ( .D(n660), .CK(clk), .Q(\mem[2][20] ) );
  DFF_X1 \mem_reg[2][19]  ( .D(n659), .CK(clk), .Q(\mem[2][19] ) );
  DFF_X1 \mem_reg[2][18]  ( .D(n658), .CK(clk), .Q(\mem[2][18] ) );
  DFF_X1 \mem_reg[2][17]  ( .D(n657), .CK(clk), .Q(\mem[2][17] ) );
  DFF_X1 \mem_reg[2][16]  ( .D(n656), .CK(clk), .Q(\mem[2][16] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n653), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n646), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n645), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n644), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n643), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n642), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n641), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n640), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[0][28]  ( .D(n604), .CK(clk), .Q(\mem[0][28] ) );
  DFF_X1 \mem_reg[0][27]  ( .D(n603), .CK(clk), .Q(\mem[0][27] ) );
  DFF_X1 \mem_reg[0][26]  ( .D(n602), .CK(clk), .Q(\mem[0][26] ) );
  DFF_X1 \mem_reg[0][25]  ( .D(n601), .CK(clk), .Q(\mem[0][25] ) );
  DFF_X1 \mem_reg[0][24]  ( .D(n600), .CK(clk), .Q(\mem[0][24] ) );
  DFF_X1 \mem_reg[0][23]  ( .D(n599), .CK(clk), .Q(\mem[0][23] ) );
  DFF_X1 \mem_reg[0][22]  ( .D(n598), .CK(clk), .Q(\mem[0][22] ) );
  DFF_X1 \mem_reg[0][21]  ( .D(n597), .CK(clk), .Q(\mem[0][21] ) );
  DFF_X1 \mem_reg[0][20]  ( .D(n596), .CK(clk), .Q(\mem[0][20] ) );
  DFF_X1 \mem_reg[0][19]  ( .D(n595), .CK(clk), .Q(\mem[0][19] ) );
  DFF_X1 \mem_reg[0][18]  ( .D(n594), .CK(clk), .Q(\mem[0][18] ) );
  DFF_X1 \mem_reg[0][17]  ( .D(n593), .CK(clk), .Q(\mem[0][17] ) );
  DFF_X1 \mem_reg[0][16]  ( .D(n592), .CK(clk), .Q(\mem[0][16] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n591), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n590), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n589), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n588), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n587), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n586), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n585), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n584), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n583), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n582), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n581), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n580), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n579), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n578), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n577), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n576), .CK(clk), .Q(\mem[0][0] ) );
  SDFF_X1 \data_out_reg[11]  ( .D(n1215), .SI(n1222), .SE(n1593), .CK(clk), 
        .Q(data_out[11]) );
  SDFF_X1 \data_out_reg[9]  ( .D(n1187), .SI(n1194), .SE(n1593), .CK(clk), .Q(
        data_out[9]) );
  SDFF_X1 \data_out_reg[10]  ( .D(n1201), .SI(n1208), .SE(n1593), .CK(clk), 
        .Q(data_out[10]) );
  SDFF_X1 \data_out_reg[17]  ( .D(n1299), .SI(n1306), .SE(n1593), .CK(clk), 
        .Q(data_out[17]) );
  SDFF_X1 \data_out_reg[1]  ( .D(n24), .SI(n31), .SE(n1593), .CK(clk), .Q(
        data_out[1]) );
  SDFF_X1 \data_out_reg[23]  ( .D(n1383), .SI(n1390), .SE(n1593), .CK(clk), 
        .Q(data_out[23]) );
  SDFF_X1 \data_out_reg[13]  ( .D(n1243), .SI(n1250), .SE(n1593), .CK(clk), 
        .Q(data_out[13]) );
  SDFF_X1 \data_out_reg[0]  ( .D(n10), .SI(n17), .SE(n1593), .CK(clk), .Q(
        data_out[0]) );
  SDFF_X1 \data_out_reg[15]  ( .D(n1271), .SI(n1278), .SE(n1593), .CK(clk), 
        .Q(data_out[15]) );
  SDFF_X1 \data_out_reg[18]  ( .D(n1313), .SI(n1320), .SE(n1593), .CK(clk), 
        .Q(data_out[18]) );
  SDFF_X1 \data_out_reg[3]  ( .D(n1103), .SI(n1110), .SE(n1593), .CK(clk), .Q(
        data_out[3]) );
  SDFF_X1 \data_out_reg[14]  ( .D(n1257), .SI(n1264), .SE(n1593), .CK(clk), 
        .Q(data_out[14]) );
  SDFF_X1 \data_out_reg[25]  ( .D(n1411), .SI(n1418), .SE(n1593), .CK(clk), 
        .Q(data_out[25]) );
  SDFF_X1 \data_out_reg[21]  ( .D(n1355), .SI(n1362), .SE(n1593), .CK(clk), 
        .Q(data_out[21]) );
  SDFF_X1 \data_out_reg[7]  ( .D(n1159), .SI(n1166), .SE(n1593), .CK(clk), .Q(
        data_out[7]) );
  SDFF_X1 \data_out_reg[5]  ( .D(n1131), .SI(n1138), .SE(n1593), .CK(clk), .Q(
        data_out[5]) );
  SDFF_X1 \data_out_reg[12]  ( .D(n1229), .SI(n1236), .SE(n1593), .CK(clk), 
        .Q(data_out[12]) );
  SDFF_X1 \data_out_reg[22]  ( .D(n1369), .SI(n1376), .SE(n1593), .CK(clk), 
        .Q(data_out[22]) );
  SDFF_X1 \data_out_reg[4]  ( .D(n1117), .SI(n1124), .SE(n1593), .CK(clk), .Q(
        data_out[4]) );
  DFF_X1 \mem_reg[1][15]  ( .D(n623), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n622), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n620), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n619), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n618), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n617), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n616), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n615), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][31]  ( .D(n639), .CK(clk), .Q(\mem[1][31] ) );
  DFF_X1 \mem_reg[1][30]  ( .D(n638), .CK(clk), .Q(\mem[1][30] ) );
  DFF_X1 \mem_reg[1][29]  ( .D(n637), .CK(clk), .Q(\mem[1][29] ) );
  DFF_X1 \mem_reg[1][28]  ( .D(n636), .CK(clk), .Q(\mem[1][28] ) );
  DFF_X1 \mem_reg[1][27]  ( .D(n635), .CK(clk), .Q(\mem[1][27] ) );
  DFF_X1 \mem_reg[1][26]  ( .D(n634), .CK(clk), .Q(\mem[1][26] ) );
  DFF_X1 \mem_reg[1][25]  ( .D(n633), .CK(clk), .Q(\mem[1][25] ) );
  DFF_X1 \mem_reg[1][24]  ( .D(n632), .CK(clk), .Q(\mem[1][24] ) );
  DFF_X1 \mem_reg[1][23]  ( .D(n631), .CK(clk), .Q(\mem[1][23] ) );
  DFF_X1 \mem_reg[1][22]  ( .D(n630), .CK(clk), .Q(\mem[1][22] ) );
  DFF_X1 \mem_reg[1][21]  ( .D(n629), .CK(clk), .Q(\mem[1][21] ) );
  DFF_X1 \mem_reg[1][20]  ( .D(n628), .CK(clk), .Q(\mem[1][20] ) );
  DFF_X1 \mem_reg[1][19]  ( .D(n627), .CK(clk), .Q(\mem[1][19] ) );
  DFF_X1 \mem_reg[1][18]  ( .D(n626), .CK(clk), .Q(\mem[1][18] ) );
  DFF_X1 \mem_reg[1][17]  ( .D(n625), .CK(clk), .Q(\mem[1][17] ) );
  DFF_X1 \mem_reg[1][16]  ( .D(n624), .CK(clk), .Q(\mem[1][16] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n621), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n614), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n613), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n612), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n611), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n610), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n609), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n608), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n783), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n782), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n780), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n779), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n778), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n777), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n776), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n775), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n719), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n718), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n716), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n715), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n714), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n713), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n712), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n711), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n655), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n654), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n652), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n651), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n650), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n649), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n648), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n647), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[0][31]  ( .D(n607), .CK(clk), .Q(\mem[0][31] ) );
  DFF_X1 \mem_reg[0][30]  ( .D(n606), .CK(clk), .Q(\mem[0][30] ) );
  DFF_X1 \mem_reg[0][29]  ( .D(n605), .CK(clk), .Q(\mem[0][29] ) );
  SDFF_X1 \data_out_reg[30]  ( .D(n1488), .SI(n1481), .SE(N13), .CK(clk), .Q(
        data_out[30]) );
  SDFF_X1 \data_out_reg[19]  ( .D(n1334), .SI(n1327), .SE(N13), .CK(clk), .Q(
        data_out[19]) );
  SDFF_X2 \data_out_reg[27]  ( .D(n1439), .SI(n1446), .SE(n1593), .CK(clk), 
        .Q(data_out[27]) );
  INV_X2 U3 ( .A(n1), .ZN(data_out[29]) );
  BUF_X1 U4 ( .A(N10), .Z(n1511) );
  BUF_X1 U5 ( .A(n1510), .Z(n1507) );
  BUF_X1 U6 ( .A(n1510), .Z(n1506) );
  NAND2_X1 U7 ( .A1(n105), .A2(n70), .ZN(n72) );
  NAND2_X1 U8 ( .A1(n70), .A2(n71), .ZN(n37) );
  NAND2_X1 U9 ( .A1(n139), .A2(n71), .ZN(n106) );
  NAND2_X1 U10 ( .A1(n139), .A2(n105), .ZN(n140) );
  NAND2_X1 U11 ( .A1(n206), .A2(n71), .ZN(n173) );
  NAND2_X1 U12 ( .A1(n206), .A2(n105), .ZN(n207) );
  NAND2_X1 U13 ( .A1(n273), .A2(n71), .ZN(n240) );
  NAND2_X1 U14 ( .A1(n273), .A2(n105), .ZN(n275) );
  NAND2_X1 U15 ( .A1(n342), .A2(n70), .ZN(n309) );
  NAND2_X1 U16 ( .A1(n376), .A2(n70), .ZN(n343) );
  NAND2_X1 U17 ( .A1(n342), .A2(n139), .ZN(n377) );
  NAND2_X1 U18 ( .A1(n376), .A2(n139), .ZN(n410) );
  NAND2_X1 U19 ( .A1(n342), .A2(n206), .ZN(n443) );
  NAND2_X1 U20 ( .A1(n376), .A2(n206), .ZN(n476) );
  NAND2_X1 U21 ( .A1(n342), .A2(n273), .ZN(n509) );
  NAND2_X1 U22 ( .A1(n376), .A2(n273), .ZN(n543) );
  BUF_X1 U23 ( .A(n1525), .Z(n1515) );
  BUF_X1 U24 ( .A(n1525), .Z(n1516) );
  BUF_X1 U25 ( .A(n1525), .Z(n1517) );
  BUF_X1 U26 ( .A(n1526), .Z(n1521) );
  BUF_X1 U27 ( .A(n1526), .Z(n1522) );
  BUF_X1 U28 ( .A(n1526), .Z(n1523) );
  BUF_X1 U29 ( .A(n1525), .Z(n1514) );
  BUF_X1 U30 ( .A(n1526), .Z(n1518) );
  BUF_X1 U31 ( .A(n1526), .Z(n1519) );
  BUF_X1 U32 ( .A(n1526), .Z(n1520) );
  BUF_X1 U33 ( .A(N10), .Z(n1512) );
  BUF_X1 U34 ( .A(N10), .Z(n1513) );
  BUF_X1 U35 ( .A(n1524), .Z(n1525) );
  BUF_X1 U36 ( .A(n1524), .Z(n1526) );
  BUF_X1 U37 ( .A(N10), .Z(n1524) );
  BUF_X1 U38 ( .A(n1510), .Z(n1508) );
  BUF_X1 U39 ( .A(N11), .Z(n1509) );
  BUF_X1 U40 ( .A(n72), .Z(n1584) );
  BUF_X1 U41 ( .A(n72), .Z(n1583) );
  BUF_X1 U42 ( .A(n309), .Z(n1556) );
  BUF_X1 U43 ( .A(n309), .Z(n1555) );
  BUF_X1 U44 ( .A(n343), .Z(n1552) );
  BUF_X1 U45 ( .A(n343), .Z(n1551) );
  BUF_X1 U46 ( .A(n377), .Z(n1548) );
  BUF_X1 U47 ( .A(n377), .Z(n1547) );
  BUF_X1 U48 ( .A(n410), .Z(n1544) );
  BUF_X1 U49 ( .A(n410), .Z(n1543) );
  BUF_X1 U50 ( .A(n37), .Z(n1588) );
  BUF_X1 U51 ( .A(n37), .Z(n1587) );
  BUF_X1 U52 ( .A(n140), .Z(n1576) );
  BUF_X1 U53 ( .A(n140), .Z(n1575) );
  BUF_X1 U54 ( .A(n173), .Z(n1572) );
  BUF_X1 U55 ( .A(n173), .Z(n1571) );
  BUF_X1 U56 ( .A(n240), .Z(n1564) );
  BUF_X1 U57 ( .A(n240), .Z(n1563) );
  BUF_X1 U58 ( .A(n275), .Z(n1560) );
  BUF_X1 U59 ( .A(n275), .Z(n1559) );
  BUF_X1 U60 ( .A(n443), .Z(n1540) );
  BUF_X1 U61 ( .A(n443), .Z(n1539) );
  BUF_X1 U62 ( .A(n476), .Z(n1536) );
  BUF_X1 U63 ( .A(n476), .Z(n1535) );
  BUF_X1 U64 ( .A(n509), .Z(n1532) );
  BUF_X1 U65 ( .A(n509), .Z(n1531) );
  BUF_X1 U66 ( .A(n37), .Z(n1589) );
  BUF_X1 U67 ( .A(n37), .Z(n1590) );
  BUF_X1 U68 ( .A(n309), .Z(n1557) );
  BUF_X1 U69 ( .A(n343), .Z(n1553) );
  BUF_X1 U70 ( .A(n377), .Z(n1549) );
  BUF_X1 U71 ( .A(n106), .Z(n1579) );
  BUF_X1 U72 ( .A(n140), .Z(n1577) );
  BUF_X1 U73 ( .A(n173), .Z(n1573) );
  BUF_X1 U74 ( .A(n207), .Z(n1567) );
  BUF_X1 U75 ( .A(n240), .Z(n1565) );
  BUF_X1 U76 ( .A(n275), .Z(n1561) );
  BUF_X1 U77 ( .A(n476), .Z(n1537) );
  BUF_X1 U78 ( .A(n509), .Z(n1533) );
  BUF_X1 U79 ( .A(n543), .Z(n1527) );
  BUF_X1 U80 ( .A(n72), .Z(n1585) );
  BUF_X1 U81 ( .A(n309), .Z(n1558) );
  BUF_X1 U82 ( .A(n343), .Z(n1554) );
  BUF_X1 U83 ( .A(n377), .Z(n1550) );
  BUF_X1 U84 ( .A(n410), .Z(n1545) );
  BUF_X1 U85 ( .A(n106), .Z(n1580) );
  BUF_X1 U86 ( .A(n106), .Z(n1581) );
  BUF_X1 U87 ( .A(n140), .Z(n1578) );
  BUF_X1 U88 ( .A(n173), .Z(n1574) );
  BUF_X1 U89 ( .A(n207), .Z(n1568) );
  BUF_X1 U90 ( .A(n207), .Z(n1569) );
  BUF_X1 U91 ( .A(n240), .Z(n1566) );
  BUF_X1 U92 ( .A(n275), .Z(n1562) );
  BUF_X1 U93 ( .A(n443), .Z(n1541) );
  BUF_X1 U94 ( .A(n476), .Z(n1538) );
  BUF_X1 U95 ( .A(n509), .Z(n1534) );
  BUF_X1 U96 ( .A(n543), .Z(n1528) );
  BUF_X1 U97 ( .A(n543), .Z(n1529) );
  AND2_X1 U98 ( .A1(n274), .A2(n1591), .ZN(n71) );
  AND2_X1 U99 ( .A1(N10), .A2(n274), .ZN(n105) );
  AND2_X1 U100 ( .A1(n542), .A2(N10), .ZN(n376) );
  AND2_X1 U101 ( .A1(n542), .A2(n1591), .ZN(n342) );
  BUF_X1 U102 ( .A(N11), .Z(n1510) );
  NOR2_X1 U103 ( .A1(n308), .A2(N13), .ZN(n274) );
  NOR2_X1 U104 ( .A1(n1593), .A2(n308), .ZN(n542) );
  NOR2_X1 U105 ( .A1(N11), .A2(N12), .ZN(n70) );
  NOR2_X1 U106 ( .A1(n1592), .A2(N12), .ZN(n139) );
  INV_X1 U107 ( .A(data_in[0]), .ZN(n1626) );
  INV_X1 U108 ( .A(data_in[1]), .ZN(n1625) );
  INV_X1 U109 ( .A(data_in[2]), .ZN(n1624) );
  INV_X1 U110 ( .A(data_in[3]), .ZN(n1623) );
  INV_X1 U111 ( .A(data_in[4]), .ZN(n1622) );
  INV_X1 U112 ( .A(data_in[5]), .ZN(n1621) );
  INV_X1 U113 ( .A(data_in[6]), .ZN(n1620) );
  INV_X1 U114 ( .A(data_in[7]), .ZN(n1619) );
  INV_X1 U115 ( .A(data_in[8]), .ZN(n1618) );
  INV_X1 U116 ( .A(data_in[9]), .ZN(n1617) );
  INV_X1 U117 ( .A(data_in[10]), .ZN(n1616) );
  INV_X1 U118 ( .A(data_in[11]), .ZN(n1615) );
  INV_X1 U119 ( .A(data_in[12]), .ZN(n1614) );
  INV_X1 U120 ( .A(data_in[13]), .ZN(n1613) );
  INV_X1 U121 ( .A(data_in[14]), .ZN(n1612) );
  INV_X1 U122 ( .A(data_in[15]), .ZN(n1611) );
  INV_X1 U123 ( .A(data_in[16]), .ZN(n1610) );
  INV_X1 U124 ( .A(data_in[17]), .ZN(n1609) );
  INV_X1 U125 ( .A(data_in[18]), .ZN(n1608) );
  INV_X1 U126 ( .A(data_in[19]), .ZN(n1607) );
  INV_X1 U127 ( .A(data_in[20]), .ZN(n1606) );
  INV_X1 U128 ( .A(data_in[21]), .ZN(n1605) );
  INV_X1 U129 ( .A(data_in[22]), .ZN(n1604) );
  INV_X1 U130 ( .A(data_in[23]), .ZN(n1603) );
  INV_X1 U131 ( .A(data_in[24]), .ZN(n1602) );
  INV_X1 U132 ( .A(data_in[25]), .ZN(n1601) );
  INV_X1 U133 ( .A(data_in[26]), .ZN(n1600) );
  INV_X1 U134 ( .A(data_in[27]), .ZN(n1599) );
  INV_X1 U135 ( .A(data_in[28]), .ZN(n1598) );
  INV_X1 U136 ( .A(data_in[29]), .ZN(n1597) );
  INV_X1 U137 ( .A(data_in[30]), .ZN(n1596) );
  INV_X1 U138 ( .A(data_in[31]), .ZN(n1595) );
  BUF_X1 U139 ( .A(N12), .Z(n1504) );
  BUF_X1 U140 ( .A(N12), .Z(n1505) );
  AND2_X1 U141 ( .A1(N12), .A2(n1592), .ZN(n206) );
  AND2_X1 U142 ( .A1(N12), .A2(N11), .ZN(n273) );
  OAI21_X1 U143 ( .B1(n1599), .B2(n1582), .A(n134), .ZN(n667) );
  NAND2_X1 U144 ( .A1(\mem[2][27] ), .A2(n1582), .ZN(n134) );
  OAI21_X1 U145 ( .B1(n1598), .B2(n1582), .A(n135), .ZN(n668) );
  NAND2_X1 U146 ( .A1(\mem[2][28] ), .A2(n1582), .ZN(n135) );
  OAI21_X1 U147 ( .B1(n1597), .B2(n1582), .A(n136), .ZN(n669) );
  NAND2_X1 U148 ( .A1(\mem[2][29] ), .A2(n1582), .ZN(n136) );
  OAI21_X1 U149 ( .B1(n1596), .B2(n1582), .A(n137), .ZN(n670) );
  NAND2_X1 U150 ( .A1(\mem[2][30] ), .A2(n1582), .ZN(n137) );
  OAI21_X1 U151 ( .B1(n1599), .B2(n1578), .A(n168), .ZN(n699) );
  NAND2_X1 U152 ( .A1(\mem[3][27] ), .A2(n1575), .ZN(n168) );
  OAI21_X1 U153 ( .B1(n1598), .B2(n140), .A(n169), .ZN(n700) );
  NAND2_X1 U154 ( .A1(\mem[3][28] ), .A2(n1575), .ZN(n169) );
  OAI21_X1 U155 ( .B1(n1597), .B2(n1578), .A(n170), .ZN(n701) );
  NAND2_X1 U156 ( .A1(\mem[3][29] ), .A2(n1575), .ZN(n170) );
  OAI21_X1 U157 ( .B1(n1596), .B2(n140), .A(n171), .ZN(n702) );
  NAND2_X1 U158 ( .A1(\mem[3][30] ), .A2(n1575), .ZN(n171) );
  OAI21_X1 U159 ( .B1(n1599), .B2(n1586), .A(n100), .ZN(n635) );
  NAND2_X1 U160 ( .A1(\mem[1][27] ), .A2(n1583), .ZN(n100) );
  OAI21_X1 U161 ( .B1(n1598), .B2(n1586), .A(n101), .ZN(n636) );
  NAND2_X1 U162 ( .A1(\mem[1][28] ), .A2(n1583), .ZN(n101) );
  OAI21_X1 U163 ( .B1(n1597), .B2(n1586), .A(n102), .ZN(n637) );
  NAND2_X1 U164 ( .A1(\mem[1][29] ), .A2(n1583), .ZN(n102) );
  OAI21_X1 U165 ( .B1(n1596), .B2(n1586), .A(n103), .ZN(n638) );
  NAND2_X1 U166 ( .A1(\mem[1][30] ), .A2(n1583), .ZN(n103) );
  OAI21_X1 U167 ( .B1(n1599), .B2(n1558), .A(n337), .ZN(n859) );
  NAND2_X1 U168 ( .A1(\mem[8][27] ), .A2(n1555), .ZN(n337) );
  OAI21_X1 U169 ( .B1(n1598), .B2(n309), .A(n338), .ZN(n860) );
  NAND2_X1 U170 ( .A1(\mem[8][28] ), .A2(n1555), .ZN(n338) );
  OAI21_X1 U171 ( .B1(n1597), .B2(n1558), .A(n339), .ZN(n861) );
  NAND2_X1 U172 ( .A1(\mem[8][29] ), .A2(n1555), .ZN(n339) );
  OAI21_X1 U173 ( .B1(n1596), .B2(n309), .A(n340), .ZN(n862) );
  NAND2_X1 U174 ( .A1(\mem[8][30] ), .A2(n1555), .ZN(n340) );
  OAI21_X1 U175 ( .B1(n1599), .B2(n1554), .A(n371), .ZN(n891) );
  NAND2_X1 U176 ( .A1(\mem[9][27] ), .A2(n1551), .ZN(n371) );
  OAI21_X1 U177 ( .B1(n1598), .B2(n343), .A(n372), .ZN(n892) );
  NAND2_X1 U178 ( .A1(\mem[9][28] ), .A2(n1551), .ZN(n372) );
  OAI21_X1 U179 ( .B1(n1597), .B2(n1554), .A(n373), .ZN(n893) );
  NAND2_X1 U180 ( .A1(\mem[9][29] ), .A2(n1551), .ZN(n373) );
  OAI21_X1 U181 ( .B1(n1596), .B2(n343), .A(n374), .ZN(n894) );
  NAND2_X1 U182 ( .A1(\mem[9][30] ), .A2(n1551), .ZN(n374) );
  OAI21_X1 U183 ( .B1(n1599), .B2(n1550), .A(n405), .ZN(n923) );
  NAND2_X1 U184 ( .A1(\mem[10][27] ), .A2(n1547), .ZN(n405) );
  OAI21_X1 U185 ( .B1(n1598), .B2(n377), .A(n406), .ZN(n924) );
  NAND2_X1 U186 ( .A1(\mem[10][28] ), .A2(n1547), .ZN(n406) );
  OAI21_X1 U187 ( .B1(n1597), .B2(n1550), .A(n407), .ZN(n925) );
  NAND2_X1 U188 ( .A1(\mem[10][29] ), .A2(n1547), .ZN(n407) );
  OAI21_X1 U189 ( .B1(n1596), .B2(n377), .A(n408), .ZN(n926) );
  NAND2_X1 U190 ( .A1(\mem[10][30] ), .A2(n1547), .ZN(n408) );
  OAI21_X1 U191 ( .B1(n1599), .B2(n1546), .A(n438), .ZN(n955) );
  NAND2_X1 U192 ( .A1(\mem[11][27] ), .A2(n1543), .ZN(n438) );
  OAI21_X1 U193 ( .B1(n1598), .B2(n1546), .A(n439), .ZN(n956) );
  NAND2_X1 U194 ( .A1(\mem[11][28] ), .A2(n1543), .ZN(n439) );
  OAI21_X1 U195 ( .B1(n1597), .B2(n1546), .A(n440), .ZN(n957) );
  NAND2_X1 U196 ( .A1(\mem[11][29] ), .A2(n1543), .ZN(n440) );
  OAI21_X1 U197 ( .B1(n1596), .B2(n1546), .A(n441), .ZN(n958) );
  NAND2_X1 U198 ( .A1(\mem[11][30] ), .A2(n1543), .ZN(n441) );
  OAI21_X1 U199 ( .B1(n1599), .B2(n1574), .A(n201), .ZN(n731) );
  NAND2_X1 U200 ( .A1(\mem[4][27] ), .A2(n1571), .ZN(n201) );
  OAI21_X1 U201 ( .B1(n1598), .B2(n173), .A(n202), .ZN(n732) );
  NAND2_X1 U202 ( .A1(\mem[4][28] ), .A2(n1571), .ZN(n202) );
  OAI21_X1 U203 ( .B1(n1597), .B2(n1574), .A(n203), .ZN(n733) );
  NAND2_X1 U204 ( .A1(\mem[4][29] ), .A2(n1571), .ZN(n203) );
  OAI21_X1 U205 ( .B1(n1596), .B2(n173), .A(n204), .ZN(n734) );
  NAND2_X1 U206 ( .A1(\mem[4][30] ), .A2(n1571), .ZN(n204) );
  OAI21_X1 U207 ( .B1(n1599), .B2(n1570), .A(n235), .ZN(n763) );
  NAND2_X1 U208 ( .A1(\mem[5][27] ), .A2(n1570), .ZN(n235) );
  OAI21_X1 U209 ( .B1(n1598), .B2(n1570), .A(n236), .ZN(n764) );
  NAND2_X1 U210 ( .A1(\mem[5][28] ), .A2(n1570), .ZN(n236) );
  OAI21_X1 U211 ( .B1(n1597), .B2(n1570), .A(n237), .ZN(n765) );
  NAND2_X1 U212 ( .A1(\mem[5][29] ), .A2(n1570), .ZN(n237) );
  OAI21_X1 U213 ( .B1(n1596), .B2(n1570), .A(n238), .ZN(n766) );
  NAND2_X1 U214 ( .A1(\mem[5][30] ), .A2(n1570), .ZN(n238) );
  OAI21_X1 U215 ( .B1(n1599), .B2(n1566), .A(n268), .ZN(n795) );
  NAND2_X1 U216 ( .A1(\mem[6][27] ), .A2(n1563), .ZN(n268) );
  OAI21_X1 U217 ( .B1(n1598), .B2(n240), .A(n269), .ZN(n796) );
  NAND2_X1 U218 ( .A1(\mem[6][28] ), .A2(n1563), .ZN(n269) );
  OAI21_X1 U219 ( .B1(n1597), .B2(n1566), .A(n270), .ZN(n797) );
  NAND2_X1 U220 ( .A1(\mem[6][29] ), .A2(n1563), .ZN(n270) );
  OAI21_X1 U221 ( .B1(n1596), .B2(n240), .A(n271), .ZN(n798) );
  NAND2_X1 U222 ( .A1(\mem[6][30] ), .A2(n1563), .ZN(n271) );
  OAI21_X1 U223 ( .B1(n1599), .B2(n1562), .A(n303), .ZN(n827) );
  NAND2_X1 U224 ( .A1(\mem[7][27] ), .A2(n1559), .ZN(n303) );
  OAI21_X1 U225 ( .B1(n1598), .B2(n275), .A(n304), .ZN(n828) );
  NAND2_X1 U226 ( .A1(\mem[7][28] ), .A2(n1559), .ZN(n304) );
  OAI21_X1 U227 ( .B1(n1597), .B2(n1562), .A(n305), .ZN(n829) );
  NAND2_X1 U228 ( .A1(\mem[7][29] ), .A2(n1559), .ZN(n305) );
  OAI21_X1 U229 ( .B1(n1596), .B2(n275), .A(n306), .ZN(n830) );
  NAND2_X1 U230 ( .A1(\mem[7][30] ), .A2(n1559), .ZN(n306) );
  OAI21_X1 U231 ( .B1(n1599), .B2(n1542), .A(n471), .ZN(n987) );
  NAND2_X1 U232 ( .A1(\mem[12][27] ), .A2(n1539), .ZN(n471) );
  OAI21_X1 U233 ( .B1(n1598), .B2(n1542), .A(n472), .ZN(n988) );
  NAND2_X1 U234 ( .A1(\mem[12][28] ), .A2(n1539), .ZN(n472) );
  OAI21_X1 U235 ( .B1(n1597), .B2(n1542), .A(n473), .ZN(n989) );
  NAND2_X1 U236 ( .A1(\mem[12][29] ), .A2(n1539), .ZN(n473) );
  OAI21_X1 U237 ( .B1(n1596), .B2(n1542), .A(n474), .ZN(n990) );
  NAND2_X1 U238 ( .A1(\mem[12][30] ), .A2(n1539), .ZN(n474) );
  OAI21_X1 U239 ( .B1(n1599), .B2(n1538), .A(n504), .ZN(n1019) );
  NAND2_X1 U240 ( .A1(\mem[13][27] ), .A2(n1535), .ZN(n504) );
  OAI21_X1 U241 ( .B1(n1598), .B2(n476), .A(n505), .ZN(n1020) );
  NAND2_X1 U242 ( .A1(\mem[13][28] ), .A2(n1535), .ZN(n505) );
  OAI21_X1 U243 ( .B1(n1597), .B2(n1538), .A(n506), .ZN(n1021) );
  NAND2_X1 U244 ( .A1(\mem[13][29] ), .A2(n1535), .ZN(n506) );
  OAI21_X1 U245 ( .B1(n1596), .B2(n476), .A(n507), .ZN(n1022) );
  NAND2_X1 U246 ( .A1(\mem[13][30] ), .A2(n1535), .ZN(n507) );
  OAI21_X1 U247 ( .B1(n1599), .B2(n1534), .A(n537), .ZN(n1051) );
  NAND2_X1 U248 ( .A1(\mem[14][27] ), .A2(n1531), .ZN(n537) );
  OAI21_X1 U249 ( .B1(n1598), .B2(n509), .A(n538), .ZN(n1052) );
  NAND2_X1 U250 ( .A1(\mem[14][28] ), .A2(n1531), .ZN(n538) );
  OAI21_X1 U251 ( .B1(n1597), .B2(n1534), .A(n539), .ZN(n1053) );
  NAND2_X1 U252 ( .A1(\mem[14][29] ), .A2(n1531), .ZN(n539) );
  OAI21_X1 U253 ( .B1(n1596), .B2(n509), .A(n540), .ZN(n1054) );
  NAND2_X1 U254 ( .A1(\mem[14][30] ), .A2(n1531), .ZN(n540) );
  OAI21_X1 U255 ( .B1(n1599), .B2(n1530), .A(n571), .ZN(n1083) );
  NAND2_X1 U256 ( .A1(\mem[15][27] ), .A2(n1530), .ZN(n571) );
  OAI21_X1 U257 ( .B1(n1598), .B2(n1530), .A(n572), .ZN(n1084) );
  NAND2_X1 U258 ( .A1(\mem[15][28] ), .A2(n1530), .ZN(n572) );
  OAI21_X1 U259 ( .B1(n1597), .B2(n1530), .A(n573), .ZN(n1085) );
  NAND2_X1 U260 ( .A1(\mem[15][29] ), .A2(n1530), .ZN(n573) );
  OAI21_X1 U261 ( .B1(n1596), .B2(n1530), .A(n574), .ZN(n1086) );
  NAND2_X1 U262 ( .A1(\mem[15][30] ), .A2(n1530), .ZN(n574) );
  NAND2_X1 U263 ( .A1(wr_en), .A2(n1594), .ZN(n308) );
  INV_X1 U264 ( .A(addr[4]), .ZN(n1594) );
  OAI21_X1 U265 ( .B1(n1589), .B2(n1597), .A(n67), .ZN(n605) );
  NAND2_X1 U266 ( .A1(\mem[0][29] ), .A2(n1587), .ZN(n67) );
  OAI21_X1 U267 ( .B1(n1590), .B2(n1596), .A(n68), .ZN(n606) );
  NAND2_X1 U268 ( .A1(\mem[0][30] ), .A2(n1587), .ZN(n68) );
  OAI21_X1 U269 ( .B1(n1626), .B2(n1586), .A(n73), .ZN(n608) );
  NAND2_X1 U270 ( .A1(\mem[1][0] ), .A2(n1583), .ZN(n73) );
  OAI21_X1 U271 ( .B1(n1625), .B2(n72), .A(n74), .ZN(n609) );
  NAND2_X1 U272 ( .A1(\mem[1][1] ), .A2(n1583), .ZN(n74) );
  OAI21_X1 U273 ( .B1(n1624), .B2(n1586), .A(n75), .ZN(n610) );
  NAND2_X1 U274 ( .A1(\mem[1][2] ), .A2(n1583), .ZN(n75) );
  OAI21_X1 U275 ( .B1(n1623), .B2(n1585), .A(n76), .ZN(n611) );
  NAND2_X1 U276 ( .A1(\mem[1][3] ), .A2(n1583), .ZN(n76) );
  OAI21_X1 U277 ( .B1(n1622), .B2(n72), .A(n77), .ZN(n612) );
  NAND2_X1 U278 ( .A1(\mem[1][4] ), .A2(n1584), .ZN(n77) );
  OAI21_X1 U279 ( .B1(n1621), .B2(n1586), .A(n78), .ZN(n613) );
  NAND2_X1 U280 ( .A1(\mem[1][5] ), .A2(n1584), .ZN(n78) );
  OAI21_X1 U281 ( .B1(n1620), .B2(n1586), .A(n79), .ZN(n614) );
  NAND2_X1 U282 ( .A1(\mem[1][6] ), .A2(n1584), .ZN(n79) );
  OAI21_X1 U283 ( .B1(n1619), .B2(n1586), .A(n80), .ZN(n615) );
  NAND2_X1 U284 ( .A1(\mem[1][7] ), .A2(n1584), .ZN(n80) );
  OAI21_X1 U285 ( .B1(n1618), .B2(n1586), .A(n81), .ZN(n616) );
  NAND2_X1 U286 ( .A1(\mem[1][8] ), .A2(n1583), .ZN(n81) );
  OAI21_X1 U287 ( .B1(n1617), .B2(n1586), .A(n82), .ZN(n617) );
  NAND2_X1 U288 ( .A1(\mem[1][9] ), .A2(n72), .ZN(n82) );
  OAI21_X1 U289 ( .B1(n1616), .B2(n1586), .A(n83), .ZN(n618) );
  NAND2_X1 U290 ( .A1(\mem[1][10] ), .A2(n72), .ZN(n83) );
  OAI21_X1 U291 ( .B1(n1615), .B2(n1585), .A(n84), .ZN(n619) );
  NAND2_X1 U292 ( .A1(\mem[1][11] ), .A2(n72), .ZN(n84) );
  OAI21_X1 U293 ( .B1(n1614), .B2(n1586), .A(n85), .ZN(n620) );
  NAND2_X1 U294 ( .A1(\mem[1][12] ), .A2(n72), .ZN(n85) );
  OAI21_X1 U295 ( .B1(n1613), .B2(n1585), .A(n86), .ZN(n621) );
  NAND2_X1 U296 ( .A1(\mem[1][13] ), .A2(n1584), .ZN(n86) );
  OAI21_X1 U297 ( .B1(n1612), .B2(n1586), .A(n87), .ZN(n622) );
  NAND2_X1 U298 ( .A1(\mem[1][14] ), .A2(n72), .ZN(n87) );
  OAI21_X1 U299 ( .B1(n1611), .B2(n1585), .A(n88), .ZN(n623) );
  NAND2_X1 U300 ( .A1(\mem[1][15] ), .A2(n72), .ZN(n88) );
  OAI21_X1 U301 ( .B1(n1610), .B2(n1585), .A(n89), .ZN(n624) );
  NAND2_X1 U302 ( .A1(\mem[1][16] ), .A2(n1584), .ZN(n89) );
  OAI21_X1 U303 ( .B1(n1609), .B2(n1585), .A(n90), .ZN(n625) );
  NAND2_X1 U304 ( .A1(\mem[1][17] ), .A2(n1584), .ZN(n90) );
  OAI21_X1 U305 ( .B1(n1608), .B2(n1585), .A(n91), .ZN(n626) );
  NAND2_X1 U306 ( .A1(\mem[1][18] ), .A2(n1584), .ZN(n91) );
  OAI21_X1 U307 ( .B1(n1607), .B2(n1585), .A(n92), .ZN(n627) );
  NAND2_X1 U308 ( .A1(\mem[1][19] ), .A2(n1584), .ZN(n92) );
  OAI21_X1 U309 ( .B1(n1606), .B2(n1585), .A(n93), .ZN(n628) );
  NAND2_X1 U310 ( .A1(\mem[1][20] ), .A2(n1584), .ZN(n93) );
  OAI21_X1 U311 ( .B1(n1605), .B2(n1585), .A(n94), .ZN(n629) );
  NAND2_X1 U312 ( .A1(\mem[1][21] ), .A2(n1584), .ZN(n94) );
  OAI21_X1 U313 ( .B1(n1604), .B2(n1585), .A(n95), .ZN(n630) );
  NAND2_X1 U314 ( .A1(\mem[1][22] ), .A2(n1584), .ZN(n95) );
  OAI21_X1 U315 ( .B1(n1603), .B2(n1585), .A(n96), .ZN(n631) );
  NAND2_X1 U316 ( .A1(\mem[1][23] ), .A2(n1584), .ZN(n96) );
  OAI21_X1 U317 ( .B1(n1602), .B2(n1585), .A(n97), .ZN(n632) );
  NAND2_X1 U318 ( .A1(\mem[1][24] ), .A2(n1583), .ZN(n97) );
  OAI21_X1 U319 ( .B1(n1601), .B2(n1585), .A(n98), .ZN(n633) );
  NAND2_X1 U320 ( .A1(\mem[1][25] ), .A2(n1583), .ZN(n98) );
  OAI21_X1 U321 ( .B1(n1600), .B2(n1585), .A(n99), .ZN(n634) );
  NAND2_X1 U322 ( .A1(\mem[1][26] ), .A2(n1583), .ZN(n99) );
  OAI21_X1 U323 ( .B1(n1595), .B2(n72), .A(n104), .ZN(n639) );
  NAND2_X1 U324 ( .A1(\mem[1][31] ), .A2(n1583), .ZN(n104) );
  OAI21_X1 U325 ( .B1(n1626), .B2(n1580), .A(n107), .ZN(n640) );
  NAND2_X1 U326 ( .A1(\mem[2][0] ), .A2(n1582), .ZN(n107) );
  OAI21_X1 U327 ( .B1(n1625), .B2(n1579), .A(n108), .ZN(n641) );
  NAND2_X1 U328 ( .A1(\mem[2][1] ), .A2(n1582), .ZN(n108) );
  OAI21_X1 U329 ( .B1(n1624), .B2(n1580), .A(n109), .ZN(n642) );
  NAND2_X1 U330 ( .A1(\mem[2][2] ), .A2(n1582), .ZN(n109) );
  OAI21_X1 U331 ( .B1(n1623), .B2(n1579), .A(n110), .ZN(n643) );
  NAND2_X1 U332 ( .A1(\mem[2][3] ), .A2(n1580), .ZN(n110) );
  OAI21_X1 U333 ( .B1(n1622), .B2(n1579), .A(n111), .ZN(n644) );
  NAND2_X1 U334 ( .A1(\mem[2][4] ), .A2(n1579), .ZN(n111) );
  OAI21_X1 U335 ( .B1(n1621), .B2(n1580), .A(n112), .ZN(n645) );
  NAND2_X1 U336 ( .A1(\mem[2][5] ), .A2(n1580), .ZN(n112) );
  OAI21_X1 U337 ( .B1(n1620), .B2(n1580), .A(n113), .ZN(n646) );
  NAND2_X1 U338 ( .A1(\mem[2][6] ), .A2(n1581), .ZN(n113) );
  OAI21_X1 U339 ( .B1(n1619), .B2(n1580), .A(n114), .ZN(n647) );
  NAND2_X1 U340 ( .A1(\mem[2][7] ), .A2(n1579), .ZN(n114) );
  OAI21_X1 U341 ( .B1(n1618), .B2(n1580), .A(n115), .ZN(n648) );
  NAND2_X1 U342 ( .A1(\mem[2][8] ), .A2(n1579), .ZN(n115) );
  OAI21_X1 U343 ( .B1(n1617), .B2(n1580), .A(n116), .ZN(n649) );
  NAND2_X1 U344 ( .A1(\mem[2][9] ), .A2(n1579), .ZN(n116) );
  OAI21_X1 U345 ( .B1(n1616), .B2(n1580), .A(n117), .ZN(n650) );
  NAND2_X1 U346 ( .A1(\mem[2][10] ), .A2(n1579), .ZN(n117) );
  OAI21_X1 U347 ( .B1(n1615), .B2(n1580), .A(n118), .ZN(n651) );
  NAND2_X1 U348 ( .A1(\mem[2][11] ), .A2(n1579), .ZN(n118) );
  OAI21_X1 U349 ( .B1(n1614), .B2(n1580), .A(n119), .ZN(n652) );
  NAND2_X1 U350 ( .A1(\mem[2][12] ), .A2(n1579), .ZN(n119) );
  OAI21_X1 U351 ( .B1(n1613), .B2(n1580), .A(n120), .ZN(n653) );
  NAND2_X1 U352 ( .A1(\mem[2][13] ), .A2(n106), .ZN(n120) );
  OAI21_X1 U353 ( .B1(n1612), .B2(n1580), .A(n121), .ZN(n654) );
  NAND2_X1 U354 ( .A1(\mem[2][14] ), .A2(n1579), .ZN(n121) );
  OAI21_X1 U355 ( .B1(n1611), .B2(n1581), .A(n122), .ZN(n655) );
  NAND2_X1 U356 ( .A1(\mem[2][15] ), .A2(n1579), .ZN(n122) );
  OAI21_X1 U357 ( .B1(n1610), .B2(n1581), .A(n123), .ZN(n656) );
  NAND2_X1 U358 ( .A1(\mem[2][16] ), .A2(n106), .ZN(n123) );
  OAI21_X1 U359 ( .B1(n1609), .B2(n1581), .A(n124), .ZN(n657) );
  NAND2_X1 U360 ( .A1(\mem[2][17] ), .A2(n106), .ZN(n124) );
  OAI21_X1 U361 ( .B1(n1608), .B2(n1581), .A(n125), .ZN(n658) );
  NAND2_X1 U362 ( .A1(\mem[2][18] ), .A2(n106), .ZN(n125) );
  OAI21_X1 U363 ( .B1(n1607), .B2(n1581), .A(n126), .ZN(n659) );
  NAND2_X1 U364 ( .A1(\mem[2][19] ), .A2(n106), .ZN(n126) );
  OAI21_X1 U365 ( .B1(n1606), .B2(n1581), .A(n127), .ZN(n660) );
  NAND2_X1 U366 ( .A1(\mem[2][20] ), .A2(n106), .ZN(n127) );
  OAI21_X1 U367 ( .B1(n1605), .B2(n1581), .A(n128), .ZN(n661) );
  NAND2_X1 U368 ( .A1(\mem[2][21] ), .A2(n106), .ZN(n128) );
  OAI21_X1 U369 ( .B1(n1604), .B2(n1581), .A(n129), .ZN(n662) );
  NAND2_X1 U370 ( .A1(\mem[2][22] ), .A2(n106), .ZN(n129) );
  OAI21_X1 U371 ( .B1(n1603), .B2(n1581), .A(n130), .ZN(n663) );
  NAND2_X1 U372 ( .A1(\mem[2][23] ), .A2(n106), .ZN(n130) );
  OAI21_X1 U373 ( .B1(n1602), .B2(n1581), .A(n131), .ZN(n664) );
  NAND2_X1 U374 ( .A1(\mem[2][24] ), .A2(n1581), .ZN(n131) );
  OAI21_X1 U375 ( .B1(n1601), .B2(n1581), .A(n132), .ZN(n665) );
  NAND2_X1 U376 ( .A1(\mem[2][25] ), .A2(n106), .ZN(n132) );
  OAI21_X1 U377 ( .B1(n1600), .B2(n1581), .A(n133), .ZN(n666) );
  NAND2_X1 U378 ( .A1(\mem[2][26] ), .A2(n106), .ZN(n133) );
  OAI21_X1 U379 ( .B1(n1595), .B2(n1579), .A(n138), .ZN(n671) );
  NAND2_X1 U380 ( .A1(\mem[2][31] ), .A2(n106), .ZN(n138) );
  OAI21_X1 U381 ( .B1(n1626), .B2(n1578), .A(n141), .ZN(n672) );
  NAND2_X1 U382 ( .A1(\mem[3][0] ), .A2(n1575), .ZN(n141) );
  OAI21_X1 U383 ( .B1(n1625), .B2(n1577), .A(n142), .ZN(n673) );
  NAND2_X1 U384 ( .A1(\mem[3][1] ), .A2(n1575), .ZN(n142) );
  OAI21_X1 U385 ( .B1(n1624), .B2(n1578), .A(n143), .ZN(n674) );
  NAND2_X1 U386 ( .A1(\mem[3][2] ), .A2(n1575), .ZN(n143) );
  OAI21_X1 U387 ( .B1(n1623), .B2(n1577), .A(n144), .ZN(n675) );
  NAND2_X1 U388 ( .A1(\mem[3][3] ), .A2(n1575), .ZN(n144) );
  OAI21_X1 U389 ( .B1(n1622), .B2(n1577), .A(n145), .ZN(n676) );
  NAND2_X1 U390 ( .A1(\mem[3][4] ), .A2(n1576), .ZN(n145) );
  OAI21_X1 U391 ( .B1(n1621), .B2(n1578), .A(n146), .ZN(n677) );
  NAND2_X1 U392 ( .A1(\mem[3][5] ), .A2(n1576), .ZN(n146) );
  OAI21_X1 U393 ( .B1(n1620), .B2(n1578), .A(n147), .ZN(n678) );
  NAND2_X1 U394 ( .A1(\mem[3][6] ), .A2(n1576), .ZN(n147) );
  OAI21_X1 U395 ( .B1(n1619), .B2(n1578), .A(n148), .ZN(n679) );
  NAND2_X1 U396 ( .A1(\mem[3][7] ), .A2(n1577), .ZN(n148) );
  OAI21_X1 U397 ( .B1(n1618), .B2(n1578), .A(n149), .ZN(n680) );
  NAND2_X1 U398 ( .A1(\mem[3][8] ), .A2(n1577), .ZN(n149) );
  OAI21_X1 U399 ( .B1(n1617), .B2(n1578), .A(n150), .ZN(n681) );
  NAND2_X1 U400 ( .A1(\mem[3][9] ), .A2(n1577), .ZN(n150) );
  OAI21_X1 U401 ( .B1(n1616), .B2(n1578), .A(n151), .ZN(n682) );
  NAND2_X1 U402 ( .A1(\mem[3][10] ), .A2(n1577), .ZN(n151) );
  OAI21_X1 U403 ( .B1(n1615), .B2(n1578), .A(n152), .ZN(n683) );
  NAND2_X1 U404 ( .A1(\mem[3][11] ), .A2(n1577), .ZN(n152) );
  OAI21_X1 U405 ( .B1(n1614), .B2(n1578), .A(n153), .ZN(n684) );
  NAND2_X1 U406 ( .A1(\mem[3][12] ), .A2(n1577), .ZN(n153) );
  OAI21_X1 U407 ( .B1(n1613), .B2(n1578), .A(n154), .ZN(n685) );
  NAND2_X1 U408 ( .A1(\mem[3][13] ), .A2(n1576), .ZN(n154) );
  OAI21_X1 U409 ( .B1(n1612), .B2(n1578), .A(n155), .ZN(n686) );
  NAND2_X1 U410 ( .A1(\mem[3][14] ), .A2(n1577), .ZN(n155) );
  OAI21_X1 U411 ( .B1(n1611), .B2(n1578), .A(n156), .ZN(n687) );
  NAND2_X1 U412 ( .A1(\mem[3][15] ), .A2(n1577), .ZN(n156) );
  OAI21_X1 U413 ( .B1(n1610), .B2(n140), .A(n157), .ZN(n688) );
  NAND2_X1 U414 ( .A1(\mem[3][16] ), .A2(n1576), .ZN(n157) );
  OAI21_X1 U415 ( .B1(n1609), .B2(n140), .A(n158), .ZN(n689) );
  NAND2_X1 U416 ( .A1(\mem[3][17] ), .A2(n1576), .ZN(n158) );
  OAI21_X1 U417 ( .B1(n1608), .B2(n140), .A(n159), .ZN(n690) );
  NAND2_X1 U418 ( .A1(\mem[3][18] ), .A2(n1576), .ZN(n159) );
  OAI21_X1 U419 ( .B1(n1607), .B2(n140), .A(n160), .ZN(n691) );
  NAND2_X1 U420 ( .A1(\mem[3][19] ), .A2(n1576), .ZN(n160) );
  OAI21_X1 U421 ( .B1(n1606), .B2(n140), .A(n161), .ZN(n692) );
  NAND2_X1 U422 ( .A1(\mem[3][20] ), .A2(n1576), .ZN(n161) );
  OAI21_X1 U423 ( .B1(n1605), .B2(n140), .A(n162), .ZN(n693) );
  NAND2_X1 U424 ( .A1(\mem[3][21] ), .A2(n1576), .ZN(n162) );
  OAI21_X1 U425 ( .B1(n1604), .B2(n140), .A(n163), .ZN(n694) );
  NAND2_X1 U426 ( .A1(\mem[3][22] ), .A2(n1576), .ZN(n163) );
  OAI21_X1 U427 ( .B1(n1603), .B2(n140), .A(n164), .ZN(n695) );
  NAND2_X1 U428 ( .A1(\mem[3][23] ), .A2(n1576), .ZN(n164) );
  OAI21_X1 U429 ( .B1(n1602), .B2(n140), .A(n165), .ZN(n696) );
  NAND2_X1 U430 ( .A1(\mem[3][24] ), .A2(n1575), .ZN(n165) );
  OAI21_X1 U431 ( .B1(n1601), .B2(n140), .A(n166), .ZN(n697) );
  NAND2_X1 U432 ( .A1(\mem[3][25] ), .A2(n1575), .ZN(n166) );
  OAI21_X1 U433 ( .B1(n1600), .B2(n140), .A(n167), .ZN(n698) );
  NAND2_X1 U434 ( .A1(\mem[3][26] ), .A2(n1575), .ZN(n167) );
  OAI21_X1 U435 ( .B1(n1595), .B2(n1577), .A(n172), .ZN(n703) );
  NAND2_X1 U436 ( .A1(\mem[3][31] ), .A2(n1575), .ZN(n172) );
  OAI21_X1 U437 ( .B1(n1626), .B2(n1574), .A(n174), .ZN(n704) );
  NAND2_X1 U438 ( .A1(\mem[4][0] ), .A2(n1571), .ZN(n174) );
  OAI21_X1 U439 ( .B1(n1625), .B2(n1573), .A(n175), .ZN(n705) );
  NAND2_X1 U440 ( .A1(\mem[4][1] ), .A2(n1571), .ZN(n175) );
  OAI21_X1 U441 ( .B1(n1624), .B2(n1574), .A(n176), .ZN(n706) );
  NAND2_X1 U442 ( .A1(\mem[4][2] ), .A2(n1571), .ZN(n176) );
  OAI21_X1 U443 ( .B1(n1623), .B2(n1573), .A(n177), .ZN(n707) );
  NAND2_X1 U444 ( .A1(\mem[4][3] ), .A2(n1571), .ZN(n177) );
  OAI21_X1 U445 ( .B1(n1622), .B2(n1573), .A(n178), .ZN(n708) );
  NAND2_X1 U446 ( .A1(\mem[4][4] ), .A2(n1572), .ZN(n178) );
  OAI21_X1 U447 ( .B1(n1621), .B2(n1574), .A(n179), .ZN(n709) );
  NAND2_X1 U448 ( .A1(\mem[4][5] ), .A2(n1572), .ZN(n179) );
  OAI21_X1 U449 ( .B1(n1620), .B2(n1574), .A(n180), .ZN(n710) );
  NAND2_X1 U450 ( .A1(\mem[4][6] ), .A2(n1572), .ZN(n180) );
  OAI21_X1 U451 ( .B1(n1619), .B2(n1574), .A(n181), .ZN(n711) );
  NAND2_X1 U452 ( .A1(\mem[4][7] ), .A2(n1573), .ZN(n181) );
  OAI21_X1 U453 ( .B1(n1618), .B2(n1574), .A(n182), .ZN(n712) );
  NAND2_X1 U454 ( .A1(\mem[4][8] ), .A2(n1573), .ZN(n182) );
  OAI21_X1 U455 ( .B1(n1617), .B2(n1574), .A(n183), .ZN(n713) );
  NAND2_X1 U456 ( .A1(\mem[4][9] ), .A2(n1573), .ZN(n183) );
  OAI21_X1 U457 ( .B1(n1616), .B2(n1574), .A(n184), .ZN(n714) );
  NAND2_X1 U458 ( .A1(\mem[4][10] ), .A2(n1573), .ZN(n184) );
  OAI21_X1 U459 ( .B1(n1615), .B2(n1574), .A(n185), .ZN(n715) );
  NAND2_X1 U460 ( .A1(\mem[4][11] ), .A2(n1573), .ZN(n185) );
  OAI21_X1 U461 ( .B1(n1614), .B2(n1574), .A(n186), .ZN(n716) );
  NAND2_X1 U462 ( .A1(\mem[4][12] ), .A2(n1573), .ZN(n186) );
  OAI21_X1 U463 ( .B1(n1613), .B2(n1574), .A(n187), .ZN(n717) );
  NAND2_X1 U464 ( .A1(\mem[4][13] ), .A2(n1572), .ZN(n187) );
  OAI21_X1 U465 ( .B1(n1612), .B2(n1574), .A(n188), .ZN(n718) );
  NAND2_X1 U466 ( .A1(\mem[4][14] ), .A2(n1573), .ZN(n188) );
  OAI21_X1 U467 ( .B1(n1611), .B2(n1574), .A(n189), .ZN(n719) );
  NAND2_X1 U468 ( .A1(\mem[4][15] ), .A2(n1573), .ZN(n189) );
  OAI21_X1 U469 ( .B1(n1610), .B2(n173), .A(n190), .ZN(n720) );
  NAND2_X1 U470 ( .A1(\mem[4][16] ), .A2(n1572), .ZN(n190) );
  OAI21_X1 U471 ( .B1(n1609), .B2(n173), .A(n191), .ZN(n721) );
  NAND2_X1 U472 ( .A1(\mem[4][17] ), .A2(n1572), .ZN(n191) );
  OAI21_X1 U473 ( .B1(n1608), .B2(n173), .A(n192), .ZN(n722) );
  NAND2_X1 U474 ( .A1(\mem[4][18] ), .A2(n1572), .ZN(n192) );
  OAI21_X1 U475 ( .B1(n1607), .B2(n173), .A(n193), .ZN(n723) );
  NAND2_X1 U476 ( .A1(\mem[4][19] ), .A2(n1572), .ZN(n193) );
  OAI21_X1 U477 ( .B1(n1606), .B2(n173), .A(n194), .ZN(n724) );
  NAND2_X1 U478 ( .A1(\mem[4][20] ), .A2(n1572), .ZN(n194) );
  OAI21_X1 U479 ( .B1(n1605), .B2(n173), .A(n195), .ZN(n725) );
  NAND2_X1 U480 ( .A1(\mem[4][21] ), .A2(n1572), .ZN(n195) );
  OAI21_X1 U481 ( .B1(n1604), .B2(n173), .A(n196), .ZN(n726) );
  NAND2_X1 U482 ( .A1(\mem[4][22] ), .A2(n1572), .ZN(n196) );
  OAI21_X1 U483 ( .B1(n1603), .B2(n173), .A(n197), .ZN(n727) );
  NAND2_X1 U484 ( .A1(\mem[4][23] ), .A2(n1572), .ZN(n197) );
  OAI21_X1 U485 ( .B1(n1602), .B2(n173), .A(n198), .ZN(n728) );
  NAND2_X1 U486 ( .A1(\mem[4][24] ), .A2(n1571), .ZN(n198) );
  OAI21_X1 U487 ( .B1(n1601), .B2(n173), .A(n199), .ZN(n729) );
  NAND2_X1 U488 ( .A1(\mem[4][25] ), .A2(n1571), .ZN(n199) );
  OAI21_X1 U489 ( .B1(n1600), .B2(n173), .A(n200), .ZN(n730) );
  NAND2_X1 U490 ( .A1(\mem[4][26] ), .A2(n1571), .ZN(n200) );
  OAI21_X1 U491 ( .B1(n1595), .B2(n1573), .A(n205), .ZN(n735) );
  NAND2_X1 U492 ( .A1(\mem[4][31] ), .A2(n1571), .ZN(n205) );
  OAI21_X1 U493 ( .B1(n1626), .B2(n1568), .A(n208), .ZN(n736) );
  NAND2_X1 U494 ( .A1(\mem[5][0] ), .A2(n1570), .ZN(n208) );
  OAI21_X1 U495 ( .B1(n1625), .B2(n1567), .A(n209), .ZN(n737) );
  NAND2_X1 U496 ( .A1(\mem[5][1] ), .A2(n1570), .ZN(n209) );
  OAI21_X1 U497 ( .B1(n1624), .B2(n1568), .A(n210), .ZN(n738) );
  NAND2_X1 U498 ( .A1(\mem[5][2] ), .A2(n1570), .ZN(n210) );
  OAI21_X1 U499 ( .B1(n1623), .B2(n1567), .A(n211), .ZN(n739) );
  NAND2_X1 U500 ( .A1(\mem[5][3] ), .A2(n1568), .ZN(n211) );
  OAI21_X1 U501 ( .B1(n1622), .B2(n1567), .A(n212), .ZN(n740) );
  NAND2_X1 U502 ( .A1(\mem[5][4] ), .A2(n1567), .ZN(n212) );
  OAI21_X1 U503 ( .B1(n1621), .B2(n1568), .A(n213), .ZN(n741) );
  NAND2_X1 U504 ( .A1(\mem[5][5] ), .A2(n207), .ZN(n213) );
  OAI21_X1 U505 ( .B1(n1620), .B2(n1568), .A(n214), .ZN(n742) );
  NAND2_X1 U506 ( .A1(\mem[5][6] ), .A2(n207), .ZN(n214) );
  OAI21_X1 U507 ( .B1(n1619), .B2(n1568), .A(n215), .ZN(n743) );
  NAND2_X1 U508 ( .A1(\mem[5][7] ), .A2(n1567), .ZN(n215) );
  OAI21_X1 U509 ( .B1(n1618), .B2(n1568), .A(n216), .ZN(n744) );
  NAND2_X1 U510 ( .A1(\mem[5][8] ), .A2(n1567), .ZN(n216) );
  OAI21_X1 U511 ( .B1(n1617), .B2(n1568), .A(n217), .ZN(n745) );
  NAND2_X1 U512 ( .A1(\mem[5][9] ), .A2(n1567), .ZN(n217) );
  OAI21_X1 U513 ( .B1(n1616), .B2(n1568), .A(n218), .ZN(n746) );
  NAND2_X1 U514 ( .A1(\mem[5][10] ), .A2(n1567), .ZN(n218) );
  OAI21_X1 U515 ( .B1(n1615), .B2(n1568), .A(n219), .ZN(n747) );
  NAND2_X1 U516 ( .A1(\mem[5][11] ), .A2(n1567), .ZN(n219) );
  OAI21_X1 U517 ( .B1(n1614), .B2(n1568), .A(n220), .ZN(n748) );
  NAND2_X1 U518 ( .A1(\mem[5][12] ), .A2(n1567), .ZN(n220) );
  OAI21_X1 U519 ( .B1(n1613), .B2(n1568), .A(n221), .ZN(n749) );
  NAND2_X1 U520 ( .A1(\mem[5][13] ), .A2(n207), .ZN(n221) );
  OAI21_X1 U521 ( .B1(n1612), .B2(n1568), .A(n222), .ZN(n750) );
  NAND2_X1 U522 ( .A1(\mem[5][14] ), .A2(n1567), .ZN(n222) );
  OAI21_X1 U523 ( .B1(n1611), .B2(n1569), .A(n223), .ZN(n751) );
  NAND2_X1 U524 ( .A1(\mem[5][15] ), .A2(n1567), .ZN(n223) );
  OAI21_X1 U525 ( .B1(n1610), .B2(n1569), .A(n224), .ZN(n752) );
  NAND2_X1 U526 ( .A1(\mem[5][16] ), .A2(n207), .ZN(n224) );
  OAI21_X1 U527 ( .B1(n1609), .B2(n1569), .A(n225), .ZN(n753) );
  NAND2_X1 U528 ( .A1(\mem[5][17] ), .A2(n207), .ZN(n225) );
  OAI21_X1 U529 ( .B1(n1608), .B2(n1569), .A(n226), .ZN(n754) );
  NAND2_X1 U530 ( .A1(\mem[5][18] ), .A2(n207), .ZN(n226) );
  OAI21_X1 U531 ( .B1(n1607), .B2(n1569), .A(n227), .ZN(n755) );
  NAND2_X1 U532 ( .A1(\mem[5][19] ), .A2(n207), .ZN(n227) );
  OAI21_X1 U533 ( .B1(n1606), .B2(n1569), .A(n228), .ZN(n756) );
  NAND2_X1 U534 ( .A1(\mem[5][20] ), .A2(n207), .ZN(n228) );
  OAI21_X1 U535 ( .B1(n1605), .B2(n1569), .A(n229), .ZN(n757) );
  NAND2_X1 U536 ( .A1(\mem[5][21] ), .A2(n207), .ZN(n229) );
  OAI21_X1 U537 ( .B1(n1604), .B2(n1569), .A(n230), .ZN(n758) );
  NAND2_X1 U538 ( .A1(\mem[5][22] ), .A2(n207), .ZN(n230) );
  OAI21_X1 U539 ( .B1(n1603), .B2(n1569), .A(n231), .ZN(n759) );
  NAND2_X1 U540 ( .A1(\mem[5][23] ), .A2(n207), .ZN(n231) );
  OAI21_X1 U541 ( .B1(n1602), .B2(n1569), .A(n232), .ZN(n760) );
  NAND2_X1 U542 ( .A1(\mem[5][24] ), .A2(n1569), .ZN(n232) );
  OAI21_X1 U543 ( .B1(n1601), .B2(n1569), .A(n233), .ZN(n761) );
  NAND2_X1 U544 ( .A1(\mem[5][25] ), .A2(n207), .ZN(n233) );
  OAI21_X1 U545 ( .B1(n1600), .B2(n1569), .A(n234), .ZN(n762) );
  NAND2_X1 U546 ( .A1(\mem[5][26] ), .A2(n207), .ZN(n234) );
  OAI21_X1 U547 ( .B1(n1595), .B2(n1567), .A(n239), .ZN(n767) );
  NAND2_X1 U548 ( .A1(\mem[5][31] ), .A2(n207), .ZN(n239) );
  OAI21_X1 U549 ( .B1(n1626), .B2(n1566), .A(n241), .ZN(n768) );
  NAND2_X1 U550 ( .A1(\mem[6][0] ), .A2(n1563), .ZN(n241) );
  OAI21_X1 U551 ( .B1(n1625), .B2(n1565), .A(n242), .ZN(n769) );
  NAND2_X1 U552 ( .A1(\mem[6][1] ), .A2(n1563), .ZN(n242) );
  OAI21_X1 U553 ( .B1(n1624), .B2(n1566), .A(n243), .ZN(n770) );
  NAND2_X1 U554 ( .A1(\mem[6][2] ), .A2(n1563), .ZN(n243) );
  OAI21_X1 U555 ( .B1(n1623), .B2(n1565), .A(n244), .ZN(n771) );
  NAND2_X1 U556 ( .A1(\mem[6][3] ), .A2(n1563), .ZN(n244) );
  OAI21_X1 U557 ( .B1(n1622), .B2(n1565), .A(n245), .ZN(n772) );
  NAND2_X1 U558 ( .A1(\mem[6][4] ), .A2(n1564), .ZN(n245) );
  OAI21_X1 U559 ( .B1(n1621), .B2(n1566), .A(n246), .ZN(n773) );
  NAND2_X1 U560 ( .A1(\mem[6][5] ), .A2(n1564), .ZN(n246) );
  OAI21_X1 U561 ( .B1(n1620), .B2(n1566), .A(n247), .ZN(n774) );
  NAND2_X1 U562 ( .A1(\mem[6][6] ), .A2(n1564), .ZN(n247) );
  OAI21_X1 U563 ( .B1(n1619), .B2(n1566), .A(n248), .ZN(n775) );
  NAND2_X1 U564 ( .A1(\mem[6][7] ), .A2(n1565), .ZN(n248) );
  OAI21_X1 U565 ( .B1(n1618), .B2(n1566), .A(n249), .ZN(n776) );
  NAND2_X1 U566 ( .A1(\mem[6][8] ), .A2(n1565), .ZN(n249) );
  OAI21_X1 U567 ( .B1(n1617), .B2(n1566), .A(n250), .ZN(n777) );
  NAND2_X1 U568 ( .A1(\mem[6][9] ), .A2(n1565), .ZN(n250) );
  OAI21_X1 U569 ( .B1(n1616), .B2(n1566), .A(n251), .ZN(n778) );
  NAND2_X1 U570 ( .A1(\mem[6][10] ), .A2(n1565), .ZN(n251) );
  OAI21_X1 U571 ( .B1(n1615), .B2(n1566), .A(n252), .ZN(n779) );
  NAND2_X1 U572 ( .A1(\mem[6][11] ), .A2(n1565), .ZN(n252) );
  OAI21_X1 U573 ( .B1(n1614), .B2(n1566), .A(n253), .ZN(n780) );
  NAND2_X1 U574 ( .A1(\mem[6][12] ), .A2(n1565), .ZN(n253) );
  OAI21_X1 U575 ( .B1(n1613), .B2(n1566), .A(n254), .ZN(n781) );
  NAND2_X1 U576 ( .A1(\mem[6][13] ), .A2(n1564), .ZN(n254) );
  OAI21_X1 U577 ( .B1(n1612), .B2(n1566), .A(n255), .ZN(n782) );
  NAND2_X1 U578 ( .A1(\mem[6][14] ), .A2(n1565), .ZN(n255) );
  OAI21_X1 U579 ( .B1(n1611), .B2(n1566), .A(n256), .ZN(n783) );
  NAND2_X1 U580 ( .A1(\mem[6][15] ), .A2(n1565), .ZN(n256) );
  OAI21_X1 U581 ( .B1(n1610), .B2(n240), .A(n257), .ZN(n784) );
  NAND2_X1 U582 ( .A1(\mem[6][16] ), .A2(n1564), .ZN(n257) );
  OAI21_X1 U583 ( .B1(n1609), .B2(n240), .A(n258), .ZN(n785) );
  NAND2_X1 U584 ( .A1(\mem[6][17] ), .A2(n1564), .ZN(n258) );
  OAI21_X1 U585 ( .B1(n1608), .B2(n240), .A(n259), .ZN(n786) );
  NAND2_X1 U586 ( .A1(\mem[6][18] ), .A2(n1564), .ZN(n259) );
  OAI21_X1 U587 ( .B1(n1607), .B2(n240), .A(n260), .ZN(n787) );
  NAND2_X1 U588 ( .A1(\mem[6][19] ), .A2(n1564), .ZN(n260) );
  OAI21_X1 U589 ( .B1(n1606), .B2(n240), .A(n261), .ZN(n788) );
  NAND2_X1 U590 ( .A1(\mem[6][20] ), .A2(n1564), .ZN(n261) );
  OAI21_X1 U591 ( .B1(n1605), .B2(n240), .A(n262), .ZN(n789) );
  NAND2_X1 U592 ( .A1(\mem[6][21] ), .A2(n1564), .ZN(n262) );
  OAI21_X1 U593 ( .B1(n1604), .B2(n240), .A(n263), .ZN(n790) );
  NAND2_X1 U594 ( .A1(\mem[6][22] ), .A2(n1564), .ZN(n263) );
  OAI21_X1 U595 ( .B1(n1603), .B2(n240), .A(n264), .ZN(n791) );
  NAND2_X1 U596 ( .A1(\mem[6][23] ), .A2(n1564), .ZN(n264) );
  OAI21_X1 U597 ( .B1(n1602), .B2(n240), .A(n265), .ZN(n792) );
  NAND2_X1 U598 ( .A1(\mem[6][24] ), .A2(n1563), .ZN(n265) );
  OAI21_X1 U599 ( .B1(n1601), .B2(n240), .A(n266), .ZN(n793) );
  NAND2_X1 U600 ( .A1(\mem[6][25] ), .A2(n1563), .ZN(n266) );
  OAI21_X1 U601 ( .B1(n1600), .B2(n240), .A(n267), .ZN(n794) );
  NAND2_X1 U602 ( .A1(\mem[6][26] ), .A2(n1563), .ZN(n267) );
  OAI21_X1 U603 ( .B1(n1595), .B2(n1565), .A(n272), .ZN(n799) );
  NAND2_X1 U604 ( .A1(\mem[6][31] ), .A2(n1563), .ZN(n272) );
  OAI21_X1 U605 ( .B1(n1626), .B2(n1562), .A(n276), .ZN(n800) );
  NAND2_X1 U606 ( .A1(\mem[7][0] ), .A2(n1559), .ZN(n276) );
  OAI21_X1 U607 ( .B1(n1625), .B2(n1561), .A(n277), .ZN(n801) );
  NAND2_X1 U608 ( .A1(\mem[7][1] ), .A2(n1559), .ZN(n277) );
  OAI21_X1 U609 ( .B1(n1624), .B2(n1562), .A(n278), .ZN(n802) );
  NAND2_X1 U610 ( .A1(\mem[7][2] ), .A2(n1559), .ZN(n278) );
  OAI21_X1 U611 ( .B1(n1623), .B2(n1561), .A(n279), .ZN(n803) );
  NAND2_X1 U612 ( .A1(\mem[7][3] ), .A2(n1559), .ZN(n279) );
  OAI21_X1 U613 ( .B1(n1622), .B2(n1561), .A(n280), .ZN(n804) );
  NAND2_X1 U614 ( .A1(\mem[7][4] ), .A2(n1560), .ZN(n280) );
  OAI21_X1 U615 ( .B1(n1621), .B2(n1562), .A(n281), .ZN(n805) );
  NAND2_X1 U616 ( .A1(\mem[7][5] ), .A2(n1560), .ZN(n281) );
  OAI21_X1 U617 ( .B1(n1620), .B2(n1562), .A(n282), .ZN(n806) );
  NAND2_X1 U618 ( .A1(\mem[7][6] ), .A2(n1560), .ZN(n282) );
  OAI21_X1 U619 ( .B1(n1619), .B2(n1562), .A(n283), .ZN(n807) );
  NAND2_X1 U620 ( .A1(\mem[7][7] ), .A2(n1561), .ZN(n283) );
  OAI21_X1 U621 ( .B1(n1618), .B2(n1562), .A(n284), .ZN(n808) );
  NAND2_X1 U622 ( .A1(\mem[7][8] ), .A2(n1561), .ZN(n284) );
  OAI21_X1 U623 ( .B1(n1617), .B2(n1562), .A(n285), .ZN(n809) );
  NAND2_X1 U624 ( .A1(\mem[7][9] ), .A2(n1561), .ZN(n285) );
  OAI21_X1 U625 ( .B1(n1616), .B2(n1562), .A(n286), .ZN(n810) );
  NAND2_X1 U626 ( .A1(\mem[7][10] ), .A2(n1561), .ZN(n286) );
  OAI21_X1 U627 ( .B1(n1615), .B2(n1562), .A(n287), .ZN(n811) );
  NAND2_X1 U628 ( .A1(\mem[7][11] ), .A2(n1561), .ZN(n287) );
  OAI21_X1 U629 ( .B1(n1614), .B2(n1562), .A(n288), .ZN(n812) );
  NAND2_X1 U630 ( .A1(\mem[7][12] ), .A2(n1561), .ZN(n288) );
  OAI21_X1 U631 ( .B1(n1613), .B2(n1562), .A(n289), .ZN(n813) );
  NAND2_X1 U632 ( .A1(\mem[7][13] ), .A2(n1560), .ZN(n289) );
  OAI21_X1 U633 ( .B1(n1612), .B2(n1562), .A(n290), .ZN(n814) );
  NAND2_X1 U634 ( .A1(\mem[7][14] ), .A2(n1561), .ZN(n290) );
  OAI21_X1 U635 ( .B1(n1611), .B2(n1562), .A(n291), .ZN(n815) );
  NAND2_X1 U636 ( .A1(\mem[7][15] ), .A2(n1561), .ZN(n291) );
  OAI21_X1 U637 ( .B1(n1610), .B2(n275), .A(n292), .ZN(n816) );
  NAND2_X1 U638 ( .A1(\mem[7][16] ), .A2(n1560), .ZN(n292) );
  OAI21_X1 U639 ( .B1(n1609), .B2(n275), .A(n293), .ZN(n817) );
  NAND2_X1 U640 ( .A1(\mem[7][17] ), .A2(n1560), .ZN(n293) );
  OAI21_X1 U641 ( .B1(n1608), .B2(n275), .A(n294), .ZN(n818) );
  NAND2_X1 U642 ( .A1(\mem[7][18] ), .A2(n1560), .ZN(n294) );
  OAI21_X1 U643 ( .B1(n1607), .B2(n275), .A(n295), .ZN(n819) );
  NAND2_X1 U644 ( .A1(\mem[7][19] ), .A2(n1560), .ZN(n295) );
  OAI21_X1 U645 ( .B1(n1606), .B2(n275), .A(n296), .ZN(n820) );
  NAND2_X1 U646 ( .A1(\mem[7][20] ), .A2(n1560), .ZN(n296) );
  OAI21_X1 U647 ( .B1(n1605), .B2(n275), .A(n297), .ZN(n821) );
  NAND2_X1 U648 ( .A1(\mem[7][21] ), .A2(n1560), .ZN(n297) );
  OAI21_X1 U649 ( .B1(n1604), .B2(n275), .A(n298), .ZN(n822) );
  NAND2_X1 U650 ( .A1(\mem[7][22] ), .A2(n1560), .ZN(n298) );
  OAI21_X1 U651 ( .B1(n1603), .B2(n275), .A(n299), .ZN(n823) );
  NAND2_X1 U652 ( .A1(\mem[7][23] ), .A2(n1560), .ZN(n299) );
  OAI21_X1 U653 ( .B1(n1602), .B2(n275), .A(n300), .ZN(n824) );
  NAND2_X1 U654 ( .A1(\mem[7][24] ), .A2(n1559), .ZN(n300) );
  OAI21_X1 U655 ( .B1(n1601), .B2(n275), .A(n301), .ZN(n825) );
  NAND2_X1 U656 ( .A1(\mem[7][25] ), .A2(n1559), .ZN(n301) );
  OAI21_X1 U657 ( .B1(n1600), .B2(n275), .A(n302), .ZN(n826) );
  NAND2_X1 U658 ( .A1(\mem[7][26] ), .A2(n1559), .ZN(n302) );
  OAI21_X1 U659 ( .B1(n1595), .B2(n1561), .A(n307), .ZN(n831) );
  NAND2_X1 U660 ( .A1(\mem[7][31] ), .A2(n1559), .ZN(n307) );
  OAI21_X1 U661 ( .B1(n1626), .B2(n1558), .A(n310), .ZN(n832) );
  NAND2_X1 U662 ( .A1(\mem[8][0] ), .A2(n1555), .ZN(n310) );
  OAI21_X1 U663 ( .B1(n1625), .B2(n1557), .A(n311), .ZN(n833) );
  NAND2_X1 U664 ( .A1(\mem[8][1] ), .A2(n1555), .ZN(n311) );
  OAI21_X1 U665 ( .B1(n1624), .B2(n1558), .A(n312), .ZN(n834) );
  NAND2_X1 U666 ( .A1(\mem[8][2] ), .A2(n1555), .ZN(n312) );
  OAI21_X1 U667 ( .B1(n1623), .B2(n1557), .A(n313), .ZN(n835) );
  NAND2_X1 U668 ( .A1(\mem[8][3] ), .A2(n1555), .ZN(n313) );
  OAI21_X1 U669 ( .B1(n1622), .B2(n1557), .A(n314), .ZN(n836) );
  NAND2_X1 U670 ( .A1(\mem[8][4] ), .A2(n1556), .ZN(n314) );
  OAI21_X1 U671 ( .B1(n1621), .B2(n1558), .A(n315), .ZN(n837) );
  NAND2_X1 U672 ( .A1(\mem[8][5] ), .A2(n1556), .ZN(n315) );
  OAI21_X1 U673 ( .B1(n1620), .B2(n1558), .A(n316), .ZN(n838) );
  NAND2_X1 U674 ( .A1(\mem[8][6] ), .A2(n1556), .ZN(n316) );
  OAI21_X1 U675 ( .B1(n1619), .B2(n1558), .A(n317), .ZN(n839) );
  NAND2_X1 U676 ( .A1(\mem[8][7] ), .A2(n1557), .ZN(n317) );
  OAI21_X1 U677 ( .B1(n1618), .B2(n1558), .A(n318), .ZN(n840) );
  NAND2_X1 U678 ( .A1(\mem[8][8] ), .A2(n1557), .ZN(n318) );
  OAI21_X1 U679 ( .B1(n1617), .B2(n1558), .A(n319), .ZN(n841) );
  NAND2_X1 U680 ( .A1(\mem[8][9] ), .A2(n1557), .ZN(n319) );
  OAI21_X1 U681 ( .B1(n1616), .B2(n1558), .A(n320), .ZN(n842) );
  NAND2_X1 U682 ( .A1(\mem[8][10] ), .A2(n1557), .ZN(n320) );
  OAI21_X1 U683 ( .B1(n1615), .B2(n1558), .A(n321), .ZN(n843) );
  NAND2_X1 U684 ( .A1(\mem[8][11] ), .A2(n1557), .ZN(n321) );
  OAI21_X1 U685 ( .B1(n1614), .B2(n1558), .A(n322), .ZN(n844) );
  NAND2_X1 U686 ( .A1(\mem[8][12] ), .A2(n1557), .ZN(n322) );
  OAI21_X1 U687 ( .B1(n1613), .B2(n1558), .A(n323), .ZN(n845) );
  NAND2_X1 U688 ( .A1(\mem[8][13] ), .A2(n1556), .ZN(n323) );
  OAI21_X1 U689 ( .B1(n1612), .B2(n1558), .A(n324), .ZN(n846) );
  NAND2_X1 U690 ( .A1(\mem[8][14] ), .A2(n1557), .ZN(n324) );
  OAI21_X1 U691 ( .B1(n1611), .B2(n1558), .A(n325), .ZN(n847) );
  NAND2_X1 U692 ( .A1(\mem[8][15] ), .A2(n1557), .ZN(n325) );
  OAI21_X1 U693 ( .B1(n1610), .B2(n309), .A(n326), .ZN(n848) );
  NAND2_X1 U694 ( .A1(\mem[8][16] ), .A2(n1556), .ZN(n326) );
  OAI21_X1 U695 ( .B1(n1609), .B2(n309), .A(n327), .ZN(n849) );
  NAND2_X1 U696 ( .A1(\mem[8][17] ), .A2(n1556), .ZN(n327) );
  OAI21_X1 U697 ( .B1(n1608), .B2(n309), .A(n328), .ZN(n850) );
  NAND2_X1 U698 ( .A1(\mem[8][18] ), .A2(n1556), .ZN(n328) );
  OAI21_X1 U699 ( .B1(n1607), .B2(n309), .A(n329), .ZN(n851) );
  NAND2_X1 U700 ( .A1(\mem[8][19] ), .A2(n1556), .ZN(n329) );
  OAI21_X1 U701 ( .B1(n1606), .B2(n309), .A(n330), .ZN(n852) );
  NAND2_X1 U702 ( .A1(\mem[8][20] ), .A2(n1556), .ZN(n330) );
  OAI21_X1 U703 ( .B1(n1605), .B2(n309), .A(n331), .ZN(n853) );
  NAND2_X1 U704 ( .A1(\mem[8][21] ), .A2(n1556), .ZN(n331) );
  OAI21_X1 U705 ( .B1(n1604), .B2(n309), .A(n332), .ZN(n854) );
  NAND2_X1 U706 ( .A1(\mem[8][22] ), .A2(n1556), .ZN(n332) );
  OAI21_X1 U707 ( .B1(n1603), .B2(n309), .A(n333), .ZN(n855) );
  NAND2_X1 U708 ( .A1(\mem[8][23] ), .A2(n1556), .ZN(n333) );
  OAI21_X1 U709 ( .B1(n1602), .B2(n309), .A(n334), .ZN(n856) );
  NAND2_X1 U710 ( .A1(\mem[8][24] ), .A2(n1555), .ZN(n334) );
  OAI21_X1 U711 ( .B1(n1601), .B2(n309), .A(n335), .ZN(n857) );
  NAND2_X1 U712 ( .A1(\mem[8][25] ), .A2(n1555), .ZN(n335) );
  OAI21_X1 U713 ( .B1(n1600), .B2(n309), .A(n336), .ZN(n858) );
  NAND2_X1 U714 ( .A1(\mem[8][26] ), .A2(n1555), .ZN(n336) );
  OAI21_X1 U715 ( .B1(n1595), .B2(n1557), .A(n341), .ZN(n863) );
  NAND2_X1 U716 ( .A1(\mem[8][31] ), .A2(n1555), .ZN(n341) );
  OAI21_X1 U717 ( .B1(n1626), .B2(n1554), .A(n344), .ZN(n864) );
  NAND2_X1 U718 ( .A1(\mem[9][0] ), .A2(n1551), .ZN(n344) );
  OAI21_X1 U719 ( .B1(n1625), .B2(n1553), .A(n345), .ZN(n865) );
  NAND2_X1 U720 ( .A1(\mem[9][1] ), .A2(n1551), .ZN(n345) );
  OAI21_X1 U721 ( .B1(n1624), .B2(n1554), .A(n346), .ZN(n866) );
  NAND2_X1 U722 ( .A1(\mem[9][2] ), .A2(n1551), .ZN(n346) );
  OAI21_X1 U723 ( .B1(n1623), .B2(n1553), .A(n347), .ZN(n867) );
  NAND2_X1 U724 ( .A1(\mem[9][3] ), .A2(n1551), .ZN(n347) );
  OAI21_X1 U725 ( .B1(n1622), .B2(n1553), .A(n348), .ZN(n868) );
  NAND2_X1 U726 ( .A1(\mem[9][4] ), .A2(n1552), .ZN(n348) );
  OAI21_X1 U727 ( .B1(n1621), .B2(n1554), .A(n349), .ZN(n869) );
  NAND2_X1 U728 ( .A1(\mem[9][5] ), .A2(n1552), .ZN(n349) );
  OAI21_X1 U729 ( .B1(n1620), .B2(n1554), .A(n350), .ZN(n870) );
  NAND2_X1 U730 ( .A1(\mem[9][6] ), .A2(n1552), .ZN(n350) );
  OAI21_X1 U731 ( .B1(n1619), .B2(n1554), .A(n351), .ZN(n871) );
  NAND2_X1 U732 ( .A1(\mem[9][7] ), .A2(n1553), .ZN(n351) );
  OAI21_X1 U733 ( .B1(n1618), .B2(n1554), .A(n352), .ZN(n872) );
  NAND2_X1 U734 ( .A1(\mem[9][8] ), .A2(n1553), .ZN(n352) );
  OAI21_X1 U735 ( .B1(n1617), .B2(n1554), .A(n353), .ZN(n873) );
  NAND2_X1 U736 ( .A1(\mem[9][9] ), .A2(n1553), .ZN(n353) );
  OAI21_X1 U737 ( .B1(n1616), .B2(n1554), .A(n354), .ZN(n874) );
  NAND2_X1 U738 ( .A1(\mem[9][10] ), .A2(n1553), .ZN(n354) );
  OAI21_X1 U739 ( .B1(n1615), .B2(n1554), .A(n355), .ZN(n875) );
  NAND2_X1 U740 ( .A1(\mem[9][11] ), .A2(n1553), .ZN(n355) );
  OAI21_X1 U741 ( .B1(n1614), .B2(n1554), .A(n356), .ZN(n876) );
  NAND2_X1 U742 ( .A1(\mem[9][12] ), .A2(n1553), .ZN(n356) );
  OAI21_X1 U743 ( .B1(n1613), .B2(n1554), .A(n357), .ZN(n877) );
  NAND2_X1 U744 ( .A1(\mem[9][13] ), .A2(n1552), .ZN(n357) );
  OAI21_X1 U745 ( .B1(n1612), .B2(n1554), .A(n358), .ZN(n878) );
  NAND2_X1 U746 ( .A1(\mem[9][14] ), .A2(n1553), .ZN(n358) );
  OAI21_X1 U747 ( .B1(n1611), .B2(n1554), .A(n359), .ZN(n879) );
  NAND2_X1 U748 ( .A1(\mem[9][15] ), .A2(n1553), .ZN(n359) );
  OAI21_X1 U749 ( .B1(n1610), .B2(n343), .A(n360), .ZN(n880) );
  NAND2_X1 U750 ( .A1(\mem[9][16] ), .A2(n1552), .ZN(n360) );
  OAI21_X1 U751 ( .B1(n1609), .B2(n343), .A(n361), .ZN(n881) );
  NAND2_X1 U752 ( .A1(\mem[9][17] ), .A2(n1552), .ZN(n361) );
  OAI21_X1 U753 ( .B1(n1608), .B2(n343), .A(n362), .ZN(n882) );
  NAND2_X1 U754 ( .A1(\mem[9][18] ), .A2(n1552), .ZN(n362) );
  OAI21_X1 U755 ( .B1(n1607), .B2(n343), .A(n363), .ZN(n883) );
  NAND2_X1 U756 ( .A1(\mem[9][19] ), .A2(n1552), .ZN(n363) );
  OAI21_X1 U757 ( .B1(n1606), .B2(n343), .A(n364), .ZN(n884) );
  NAND2_X1 U758 ( .A1(\mem[9][20] ), .A2(n1552), .ZN(n364) );
  OAI21_X1 U759 ( .B1(n1605), .B2(n343), .A(n365), .ZN(n885) );
  NAND2_X1 U760 ( .A1(\mem[9][21] ), .A2(n1552), .ZN(n365) );
  OAI21_X1 U761 ( .B1(n1604), .B2(n343), .A(n366), .ZN(n886) );
  NAND2_X1 U762 ( .A1(\mem[9][22] ), .A2(n1552), .ZN(n366) );
  OAI21_X1 U763 ( .B1(n1603), .B2(n343), .A(n367), .ZN(n887) );
  NAND2_X1 U764 ( .A1(\mem[9][23] ), .A2(n1552), .ZN(n367) );
  OAI21_X1 U765 ( .B1(n1602), .B2(n343), .A(n368), .ZN(n888) );
  NAND2_X1 U766 ( .A1(\mem[9][24] ), .A2(n1551), .ZN(n368) );
  OAI21_X1 U767 ( .B1(n1601), .B2(n343), .A(n369), .ZN(n889) );
  NAND2_X1 U768 ( .A1(\mem[9][25] ), .A2(n1551), .ZN(n369) );
  OAI21_X1 U769 ( .B1(n1600), .B2(n343), .A(n370), .ZN(n890) );
  NAND2_X1 U770 ( .A1(\mem[9][26] ), .A2(n1551), .ZN(n370) );
  OAI21_X1 U771 ( .B1(n1595), .B2(n1553), .A(n375), .ZN(n895) );
  NAND2_X1 U772 ( .A1(\mem[9][31] ), .A2(n1551), .ZN(n375) );
  OAI21_X1 U773 ( .B1(n1626), .B2(n1550), .A(n378), .ZN(n896) );
  NAND2_X1 U774 ( .A1(\mem[10][0] ), .A2(n1547), .ZN(n378) );
  OAI21_X1 U775 ( .B1(n1625), .B2(n1549), .A(n379), .ZN(n897) );
  NAND2_X1 U776 ( .A1(\mem[10][1] ), .A2(n1547), .ZN(n379) );
  OAI21_X1 U777 ( .B1(n1624), .B2(n1550), .A(n380), .ZN(n898) );
  NAND2_X1 U778 ( .A1(\mem[10][2] ), .A2(n1547), .ZN(n380) );
  OAI21_X1 U779 ( .B1(n1623), .B2(n1549), .A(n381), .ZN(n899) );
  NAND2_X1 U780 ( .A1(\mem[10][3] ), .A2(n1547), .ZN(n381) );
  OAI21_X1 U781 ( .B1(n1622), .B2(n1549), .A(n382), .ZN(n900) );
  NAND2_X1 U782 ( .A1(\mem[10][4] ), .A2(n1548), .ZN(n382) );
  OAI21_X1 U783 ( .B1(n1621), .B2(n1550), .A(n383), .ZN(n901) );
  NAND2_X1 U784 ( .A1(\mem[10][5] ), .A2(n1548), .ZN(n383) );
  OAI21_X1 U785 ( .B1(n1620), .B2(n1550), .A(n384), .ZN(n902) );
  NAND2_X1 U786 ( .A1(\mem[10][6] ), .A2(n1548), .ZN(n384) );
  OAI21_X1 U787 ( .B1(n1619), .B2(n1550), .A(n385), .ZN(n903) );
  NAND2_X1 U788 ( .A1(\mem[10][7] ), .A2(n1549), .ZN(n385) );
  OAI21_X1 U789 ( .B1(n1618), .B2(n1550), .A(n386), .ZN(n904) );
  NAND2_X1 U790 ( .A1(\mem[10][8] ), .A2(n1549), .ZN(n386) );
  OAI21_X1 U791 ( .B1(n1617), .B2(n1550), .A(n387), .ZN(n905) );
  NAND2_X1 U792 ( .A1(\mem[10][9] ), .A2(n1549), .ZN(n387) );
  OAI21_X1 U793 ( .B1(n1616), .B2(n1550), .A(n388), .ZN(n906) );
  NAND2_X1 U794 ( .A1(\mem[10][10] ), .A2(n1549), .ZN(n388) );
  OAI21_X1 U795 ( .B1(n1615), .B2(n1550), .A(n389), .ZN(n907) );
  NAND2_X1 U796 ( .A1(\mem[10][11] ), .A2(n1549), .ZN(n389) );
  OAI21_X1 U797 ( .B1(n1614), .B2(n1550), .A(n390), .ZN(n908) );
  NAND2_X1 U798 ( .A1(\mem[10][12] ), .A2(n1549), .ZN(n390) );
  OAI21_X1 U799 ( .B1(n1613), .B2(n1550), .A(n391), .ZN(n909) );
  NAND2_X1 U800 ( .A1(\mem[10][13] ), .A2(n1548), .ZN(n391) );
  OAI21_X1 U801 ( .B1(n1612), .B2(n1550), .A(n392), .ZN(n910) );
  NAND2_X1 U802 ( .A1(\mem[10][14] ), .A2(n1549), .ZN(n392) );
  OAI21_X1 U803 ( .B1(n1611), .B2(n1550), .A(n393), .ZN(n911) );
  NAND2_X1 U804 ( .A1(\mem[10][15] ), .A2(n1549), .ZN(n393) );
  OAI21_X1 U805 ( .B1(n1610), .B2(n377), .A(n394), .ZN(n912) );
  NAND2_X1 U806 ( .A1(\mem[10][16] ), .A2(n1548), .ZN(n394) );
  OAI21_X1 U807 ( .B1(n1609), .B2(n377), .A(n395), .ZN(n913) );
  NAND2_X1 U808 ( .A1(\mem[10][17] ), .A2(n1548), .ZN(n395) );
  OAI21_X1 U809 ( .B1(n1608), .B2(n377), .A(n396), .ZN(n914) );
  NAND2_X1 U810 ( .A1(\mem[10][18] ), .A2(n1548), .ZN(n396) );
  OAI21_X1 U811 ( .B1(n1607), .B2(n377), .A(n397), .ZN(n915) );
  NAND2_X1 U812 ( .A1(\mem[10][19] ), .A2(n1548), .ZN(n397) );
  OAI21_X1 U813 ( .B1(n1606), .B2(n377), .A(n398), .ZN(n916) );
  NAND2_X1 U814 ( .A1(\mem[10][20] ), .A2(n1548), .ZN(n398) );
  OAI21_X1 U815 ( .B1(n1605), .B2(n377), .A(n399), .ZN(n917) );
  NAND2_X1 U816 ( .A1(\mem[10][21] ), .A2(n1548), .ZN(n399) );
  OAI21_X1 U817 ( .B1(n1604), .B2(n377), .A(n400), .ZN(n918) );
  NAND2_X1 U818 ( .A1(\mem[10][22] ), .A2(n1548), .ZN(n400) );
  OAI21_X1 U819 ( .B1(n1603), .B2(n377), .A(n401), .ZN(n919) );
  NAND2_X1 U820 ( .A1(\mem[10][23] ), .A2(n1548), .ZN(n401) );
  OAI21_X1 U821 ( .B1(n1602), .B2(n377), .A(n402), .ZN(n920) );
  NAND2_X1 U822 ( .A1(\mem[10][24] ), .A2(n1547), .ZN(n402) );
  OAI21_X1 U823 ( .B1(n1601), .B2(n377), .A(n403), .ZN(n921) );
  NAND2_X1 U824 ( .A1(\mem[10][25] ), .A2(n1547), .ZN(n403) );
  OAI21_X1 U825 ( .B1(n1600), .B2(n377), .A(n404), .ZN(n922) );
  NAND2_X1 U826 ( .A1(\mem[10][26] ), .A2(n1547), .ZN(n404) );
  OAI21_X1 U827 ( .B1(n1595), .B2(n1549), .A(n409), .ZN(n927) );
  NAND2_X1 U828 ( .A1(\mem[10][31] ), .A2(n1547), .ZN(n409) );
  OAI21_X1 U829 ( .B1(n1626), .B2(n1546), .A(n411), .ZN(n928) );
  NAND2_X1 U830 ( .A1(\mem[11][0] ), .A2(n1543), .ZN(n411) );
  OAI21_X1 U831 ( .B1(n1625), .B2(n410), .A(n412), .ZN(n929) );
  NAND2_X1 U832 ( .A1(\mem[11][1] ), .A2(n1543), .ZN(n412) );
  OAI21_X1 U833 ( .B1(n1624), .B2(n1546), .A(n413), .ZN(n930) );
  NAND2_X1 U834 ( .A1(\mem[11][2] ), .A2(n1543), .ZN(n413) );
  OAI21_X1 U835 ( .B1(n1623), .B2(n1545), .A(n414), .ZN(n931) );
  NAND2_X1 U836 ( .A1(\mem[11][3] ), .A2(n1543), .ZN(n414) );
  OAI21_X1 U837 ( .B1(n1622), .B2(n410), .A(n415), .ZN(n932) );
  NAND2_X1 U838 ( .A1(\mem[11][4] ), .A2(n1544), .ZN(n415) );
  OAI21_X1 U839 ( .B1(n1621), .B2(n1546), .A(n416), .ZN(n933) );
  NAND2_X1 U840 ( .A1(\mem[11][5] ), .A2(n1544), .ZN(n416) );
  OAI21_X1 U841 ( .B1(n1620), .B2(n1546), .A(n417), .ZN(n934) );
  NAND2_X1 U842 ( .A1(\mem[11][6] ), .A2(n1544), .ZN(n417) );
  OAI21_X1 U843 ( .B1(n1619), .B2(n1546), .A(n418), .ZN(n935) );
  NAND2_X1 U844 ( .A1(\mem[11][7] ), .A2(n1544), .ZN(n418) );
  OAI21_X1 U845 ( .B1(n1618), .B2(n1546), .A(n419), .ZN(n936) );
  NAND2_X1 U846 ( .A1(\mem[11][8] ), .A2(n1543), .ZN(n419) );
  OAI21_X1 U847 ( .B1(n1617), .B2(n1546), .A(n420), .ZN(n937) );
  NAND2_X1 U848 ( .A1(\mem[11][9] ), .A2(n410), .ZN(n420) );
  OAI21_X1 U849 ( .B1(n1616), .B2(n1546), .A(n421), .ZN(n938) );
  NAND2_X1 U850 ( .A1(\mem[11][10] ), .A2(n410), .ZN(n421) );
  OAI21_X1 U851 ( .B1(n1615), .B2(n1545), .A(n422), .ZN(n939) );
  NAND2_X1 U852 ( .A1(\mem[11][11] ), .A2(n410), .ZN(n422) );
  OAI21_X1 U853 ( .B1(n1614), .B2(n1546), .A(n423), .ZN(n940) );
  NAND2_X1 U854 ( .A1(\mem[11][12] ), .A2(n410), .ZN(n423) );
  OAI21_X1 U855 ( .B1(n1613), .B2(n1545), .A(n424), .ZN(n941) );
  NAND2_X1 U856 ( .A1(\mem[11][13] ), .A2(n1544), .ZN(n424) );
  OAI21_X1 U857 ( .B1(n1612), .B2(n1546), .A(n425), .ZN(n942) );
  NAND2_X1 U858 ( .A1(\mem[11][14] ), .A2(n410), .ZN(n425) );
  OAI21_X1 U859 ( .B1(n1611), .B2(n1545), .A(n426), .ZN(n943) );
  NAND2_X1 U860 ( .A1(\mem[11][15] ), .A2(n410), .ZN(n426) );
  OAI21_X1 U861 ( .B1(n1610), .B2(n1545), .A(n427), .ZN(n944) );
  NAND2_X1 U862 ( .A1(\mem[11][16] ), .A2(n1544), .ZN(n427) );
  OAI21_X1 U863 ( .B1(n1609), .B2(n1545), .A(n428), .ZN(n945) );
  NAND2_X1 U864 ( .A1(\mem[11][17] ), .A2(n1544), .ZN(n428) );
  OAI21_X1 U865 ( .B1(n1608), .B2(n1545), .A(n429), .ZN(n946) );
  NAND2_X1 U866 ( .A1(\mem[11][18] ), .A2(n1544), .ZN(n429) );
  OAI21_X1 U867 ( .B1(n1607), .B2(n1545), .A(n430), .ZN(n947) );
  NAND2_X1 U868 ( .A1(\mem[11][19] ), .A2(n1544), .ZN(n430) );
  OAI21_X1 U869 ( .B1(n1606), .B2(n1545), .A(n431), .ZN(n948) );
  NAND2_X1 U870 ( .A1(\mem[11][20] ), .A2(n1544), .ZN(n431) );
  OAI21_X1 U871 ( .B1(n1605), .B2(n1545), .A(n432), .ZN(n949) );
  NAND2_X1 U872 ( .A1(\mem[11][21] ), .A2(n1544), .ZN(n432) );
  OAI21_X1 U873 ( .B1(n1604), .B2(n1545), .A(n433), .ZN(n950) );
  NAND2_X1 U874 ( .A1(\mem[11][22] ), .A2(n1544), .ZN(n433) );
  OAI21_X1 U875 ( .B1(n1603), .B2(n1545), .A(n434), .ZN(n951) );
  NAND2_X1 U876 ( .A1(\mem[11][23] ), .A2(n1544), .ZN(n434) );
  OAI21_X1 U877 ( .B1(n1602), .B2(n1545), .A(n435), .ZN(n952) );
  NAND2_X1 U878 ( .A1(\mem[11][24] ), .A2(n1543), .ZN(n435) );
  OAI21_X1 U879 ( .B1(n1601), .B2(n1545), .A(n436), .ZN(n953) );
  NAND2_X1 U880 ( .A1(\mem[11][25] ), .A2(n1543), .ZN(n436) );
  OAI21_X1 U881 ( .B1(n1600), .B2(n1545), .A(n437), .ZN(n954) );
  NAND2_X1 U882 ( .A1(\mem[11][26] ), .A2(n1543), .ZN(n437) );
  OAI21_X1 U883 ( .B1(n1595), .B2(n410), .A(n442), .ZN(n959) );
  NAND2_X1 U884 ( .A1(\mem[11][31] ), .A2(n1543), .ZN(n442) );
  OAI21_X1 U885 ( .B1(n1626), .B2(n1542), .A(n444), .ZN(n960) );
  NAND2_X1 U886 ( .A1(\mem[12][0] ), .A2(n1539), .ZN(n444) );
  OAI21_X1 U887 ( .B1(n1625), .B2(n443), .A(n445), .ZN(n961) );
  NAND2_X1 U888 ( .A1(\mem[12][1] ), .A2(n1539), .ZN(n445) );
  OAI21_X1 U889 ( .B1(n1624), .B2(n1542), .A(n446), .ZN(n962) );
  NAND2_X1 U890 ( .A1(\mem[12][2] ), .A2(n1539), .ZN(n446) );
  OAI21_X1 U891 ( .B1(n1623), .B2(n1541), .A(n447), .ZN(n963) );
  NAND2_X1 U892 ( .A1(\mem[12][3] ), .A2(n1539), .ZN(n447) );
  OAI21_X1 U893 ( .B1(n1622), .B2(n443), .A(n448), .ZN(n964) );
  NAND2_X1 U894 ( .A1(\mem[12][4] ), .A2(n1540), .ZN(n448) );
  OAI21_X1 U895 ( .B1(n1621), .B2(n1542), .A(n449), .ZN(n965) );
  NAND2_X1 U896 ( .A1(\mem[12][5] ), .A2(n1540), .ZN(n449) );
  OAI21_X1 U897 ( .B1(n1620), .B2(n1542), .A(n450), .ZN(n966) );
  NAND2_X1 U898 ( .A1(\mem[12][6] ), .A2(n1540), .ZN(n450) );
  OAI21_X1 U899 ( .B1(n1619), .B2(n1542), .A(n451), .ZN(n967) );
  NAND2_X1 U900 ( .A1(\mem[12][7] ), .A2(n1540), .ZN(n451) );
  OAI21_X1 U901 ( .B1(n1618), .B2(n1542), .A(n452), .ZN(n968) );
  NAND2_X1 U902 ( .A1(\mem[12][8] ), .A2(n1539), .ZN(n452) );
  OAI21_X1 U903 ( .B1(n1617), .B2(n1542), .A(n453), .ZN(n969) );
  NAND2_X1 U904 ( .A1(\mem[12][9] ), .A2(n443), .ZN(n453) );
  OAI21_X1 U905 ( .B1(n1616), .B2(n1542), .A(n454), .ZN(n970) );
  NAND2_X1 U906 ( .A1(\mem[12][10] ), .A2(n443), .ZN(n454) );
  OAI21_X1 U907 ( .B1(n1615), .B2(n1541), .A(n455), .ZN(n971) );
  NAND2_X1 U908 ( .A1(\mem[12][11] ), .A2(n443), .ZN(n455) );
  OAI21_X1 U909 ( .B1(n1614), .B2(n1542), .A(n456), .ZN(n972) );
  NAND2_X1 U910 ( .A1(\mem[12][12] ), .A2(n443), .ZN(n456) );
  OAI21_X1 U911 ( .B1(n1613), .B2(n1541), .A(n457), .ZN(n973) );
  NAND2_X1 U912 ( .A1(\mem[12][13] ), .A2(n1540), .ZN(n457) );
  OAI21_X1 U913 ( .B1(n1612), .B2(n1542), .A(n458), .ZN(n974) );
  NAND2_X1 U914 ( .A1(\mem[12][14] ), .A2(n443), .ZN(n458) );
  OAI21_X1 U915 ( .B1(n1611), .B2(n1541), .A(n459), .ZN(n975) );
  NAND2_X1 U916 ( .A1(\mem[12][15] ), .A2(n443), .ZN(n459) );
  OAI21_X1 U917 ( .B1(n1610), .B2(n1541), .A(n460), .ZN(n976) );
  NAND2_X1 U918 ( .A1(\mem[12][16] ), .A2(n1540), .ZN(n460) );
  OAI21_X1 U919 ( .B1(n1609), .B2(n1541), .A(n461), .ZN(n977) );
  NAND2_X1 U920 ( .A1(\mem[12][17] ), .A2(n1540), .ZN(n461) );
  OAI21_X1 U921 ( .B1(n1608), .B2(n1541), .A(n462), .ZN(n978) );
  NAND2_X1 U922 ( .A1(\mem[12][18] ), .A2(n1540), .ZN(n462) );
  OAI21_X1 U923 ( .B1(n1607), .B2(n1541), .A(n463), .ZN(n979) );
  NAND2_X1 U924 ( .A1(\mem[12][19] ), .A2(n1540), .ZN(n463) );
  OAI21_X1 U925 ( .B1(n1606), .B2(n1541), .A(n464), .ZN(n980) );
  NAND2_X1 U926 ( .A1(\mem[12][20] ), .A2(n1540), .ZN(n464) );
  OAI21_X1 U927 ( .B1(n1605), .B2(n1541), .A(n465), .ZN(n981) );
  NAND2_X1 U928 ( .A1(\mem[12][21] ), .A2(n1540), .ZN(n465) );
  OAI21_X1 U929 ( .B1(n1604), .B2(n1541), .A(n466), .ZN(n982) );
  NAND2_X1 U930 ( .A1(\mem[12][22] ), .A2(n1540), .ZN(n466) );
  OAI21_X1 U931 ( .B1(n1603), .B2(n1541), .A(n467), .ZN(n983) );
  NAND2_X1 U932 ( .A1(\mem[12][23] ), .A2(n1540), .ZN(n467) );
  OAI21_X1 U933 ( .B1(n1602), .B2(n1541), .A(n468), .ZN(n984) );
  NAND2_X1 U934 ( .A1(\mem[12][24] ), .A2(n1539), .ZN(n468) );
  OAI21_X1 U935 ( .B1(n1601), .B2(n1541), .A(n469), .ZN(n985) );
  NAND2_X1 U936 ( .A1(\mem[12][25] ), .A2(n1539), .ZN(n469) );
  OAI21_X1 U937 ( .B1(n1600), .B2(n1541), .A(n470), .ZN(n986) );
  NAND2_X1 U938 ( .A1(\mem[12][26] ), .A2(n1539), .ZN(n470) );
  OAI21_X1 U939 ( .B1(n1595), .B2(n443), .A(n475), .ZN(n991) );
  NAND2_X1 U940 ( .A1(\mem[12][31] ), .A2(n1539), .ZN(n475) );
  OAI21_X1 U941 ( .B1(n1626), .B2(n1538), .A(n477), .ZN(n992) );
  NAND2_X1 U942 ( .A1(\mem[13][0] ), .A2(n1535), .ZN(n477) );
  OAI21_X1 U943 ( .B1(n1625), .B2(n1537), .A(n478), .ZN(n993) );
  NAND2_X1 U944 ( .A1(\mem[13][1] ), .A2(n1535), .ZN(n478) );
  OAI21_X1 U945 ( .B1(n1624), .B2(n1538), .A(n479), .ZN(n994) );
  NAND2_X1 U946 ( .A1(\mem[13][2] ), .A2(n1535), .ZN(n479) );
  OAI21_X1 U947 ( .B1(n1623), .B2(n1537), .A(n480), .ZN(n995) );
  NAND2_X1 U948 ( .A1(\mem[13][3] ), .A2(n1535), .ZN(n480) );
  OAI21_X1 U949 ( .B1(n1622), .B2(n1537), .A(n481), .ZN(n996) );
  NAND2_X1 U950 ( .A1(\mem[13][4] ), .A2(n1536), .ZN(n481) );
  OAI21_X1 U951 ( .B1(n1621), .B2(n1538), .A(n482), .ZN(n997) );
  NAND2_X1 U952 ( .A1(\mem[13][5] ), .A2(n1536), .ZN(n482) );
  OAI21_X1 U953 ( .B1(n1620), .B2(n1538), .A(n483), .ZN(n998) );
  NAND2_X1 U954 ( .A1(\mem[13][6] ), .A2(n1536), .ZN(n483) );
  OAI21_X1 U955 ( .B1(n1619), .B2(n1538), .A(n484), .ZN(n999) );
  NAND2_X1 U956 ( .A1(\mem[13][7] ), .A2(n1537), .ZN(n484) );
  OAI21_X1 U957 ( .B1(n1618), .B2(n1538), .A(n485), .ZN(n1000) );
  NAND2_X1 U958 ( .A1(\mem[13][8] ), .A2(n1537), .ZN(n485) );
  OAI21_X1 U959 ( .B1(n1617), .B2(n1538), .A(n486), .ZN(n1001) );
  NAND2_X1 U960 ( .A1(\mem[13][9] ), .A2(n1537), .ZN(n486) );
  OAI21_X1 U961 ( .B1(n1616), .B2(n1538), .A(n487), .ZN(n1002) );
  NAND2_X1 U962 ( .A1(\mem[13][10] ), .A2(n1537), .ZN(n487) );
  OAI21_X1 U963 ( .B1(n1615), .B2(n1538), .A(n488), .ZN(n1003) );
  NAND2_X1 U964 ( .A1(\mem[13][11] ), .A2(n1537), .ZN(n488) );
  OAI21_X1 U965 ( .B1(n1614), .B2(n1538), .A(n489), .ZN(n1004) );
  NAND2_X1 U966 ( .A1(\mem[13][12] ), .A2(n1537), .ZN(n489) );
  OAI21_X1 U967 ( .B1(n1613), .B2(n1538), .A(n490), .ZN(n1005) );
  NAND2_X1 U968 ( .A1(\mem[13][13] ), .A2(n1536), .ZN(n490) );
  OAI21_X1 U969 ( .B1(n1612), .B2(n1538), .A(n491), .ZN(n1006) );
  NAND2_X1 U970 ( .A1(\mem[13][14] ), .A2(n1537), .ZN(n491) );
  OAI21_X1 U971 ( .B1(n1611), .B2(n1538), .A(n492), .ZN(n1007) );
  NAND2_X1 U972 ( .A1(\mem[13][15] ), .A2(n1537), .ZN(n492) );
  OAI21_X1 U973 ( .B1(n1610), .B2(n476), .A(n493), .ZN(n1008) );
  NAND2_X1 U974 ( .A1(\mem[13][16] ), .A2(n1536), .ZN(n493) );
  OAI21_X1 U975 ( .B1(n1609), .B2(n476), .A(n494), .ZN(n1009) );
  NAND2_X1 U976 ( .A1(\mem[13][17] ), .A2(n1536), .ZN(n494) );
  OAI21_X1 U977 ( .B1(n1608), .B2(n476), .A(n495), .ZN(n1010) );
  NAND2_X1 U978 ( .A1(\mem[13][18] ), .A2(n1536), .ZN(n495) );
  OAI21_X1 U979 ( .B1(n1607), .B2(n476), .A(n496), .ZN(n1011) );
  NAND2_X1 U980 ( .A1(\mem[13][19] ), .A2(n1536), .ZN(n496) );
  OAI21_X1 U981 ( .B1(n1606), .B2(n476), .A(n497), .ZN(n1012) );
  NAND2_X1 U982 ( .A1(\mem[13][20] ), .A2(n1536), .ZN(n497) );
  OAI21_X1 U983 ( .B1(n1605), .B2(n476), .A(n498), .ZN(n1013) );
  NAND2_X1 U984 ( .A1(\mem[13][21] ), .A2(n1536), .ZN(n498) );
  OAI21_X1 U985 ( .B1(n1604), .B2(n476), .A(n499), .ZN(n1014) );
  NAND2_X1 U986 ( .A1(\mem[13][22] ), .A2(n1536), .ZN(n499) );
  OAI21_X1 U987 ( .B1(n1603), .B2(n476), .A(n500), .ZN(n1015) );
  NAND2_X1 U988 ( .A1(\mem[13][23] ), .A2(n1536), .ZN(n500) );
  OAI21_X1 U989 ( .B1(n1602), .B2(n476), .A(n501), .ZN(n1016) );
  NAND2_X1 U990 ( .A1(\mem[13][24] ), .A2(n1535), .ZN(n501) );
  OAI21_X1 U991 ( .B1(n1601), .B2(n476), .A(n502), .ZN(n1017) );
  NAND2_X1 U992 ( .A1(\mem[13][25] ), .A2(n1535), .ZN(n502) );
  OAI21_X1 U993 ( .B1(n1600), .B2(n476), .A(n503), .ZN(n1018) );
  NAND2_X1 U994 ( .A1(\mem[13][26] ), .A2(n1535), .ZN(n503) );
  OAI21_X1 U995 ( .B1(n1595), .B2(n1537), .A(n508), .ZN(n1023) );
  NAND2_X1 U996 ( .A1(\mem[13][31] ), .A2(n1535), .ZN(n508) );
  OAI21_X1 U997 ( .B1(n1626), .B2(n1534), .A(n510), .ZN(n1024) );
  NAND2_X1 U998 ( .A1(\mem[14][0] ), .A2(n1531), .ZN(n510) );
  OAI21_X1 U999 ( .B1(n1625), .B2(n1533), .A(n511), .ZN(n1025) );
  NAND2_X1 U1000 ( .A1(\mem[14][1] ), .A2(n1531), .ZN(n511) );
  OAI21_X1 U1001 ( .B1(n1624), .B2(n1534), .A(n512), .ZN(n1026) );
  NAND2_X1 U1002 ( .A1(\mem[14][2] ), .A2(n1531), .ZN(n512) );
  OAI21_X1 U1003 ( .B1(n1623), .B2(n1533), .A(n513), .ZN(n1027) );
  NAND2_X1 U1004 ( .A1(\mem[14][3] ), .A2(n1531), .ZN(n513) );
  OAI21_X1 U1005 ( .B1(n1622), .B2(n1533), .A(n514), .ZN(n1028) );
  NAND2_X1 U1006 ( .A1(\mem[14][4] ), .A2(n1532), .ZN(n514) );
  OAI21_X1 U1007 ( .B1(n1621), .B2(n1534), .A(n515), .ZN(n1029) );
  NAND2_X1 U1008 ( .A1(\mem[14][5] ), .A2(n1532), .ZN(n515) );
  OAI21_X1 U1009 ( .B1(n1620), .B2(n1534), .A(n516), .ZN(n1030) );
  NAND2_X1 U1010 ( .A1(\mem[14][6] ), .A2(n1532), .ZN(n516) );
  OAI21_X1 U1011 ( .B1(n1619), .B2(n1534), .A(n517), .ZN(n1031) );
  NAND2_X1 U1012 ( .A1(\mem[14][7] ), .A2(n1533), .ZN(n517) );
  OAI21_X1 U1013 ( .B1(n1618), .B2(n1534), .A(n518), .ZN(n1032) );
  NAND2_X1 U1014 ( .A1(\mem[14][8] ), .A2(n1533), .ZN(n518) );
  OAI21_X1 U1015 ( .B1(n1617), .B2(n1534), .A(n519), .ZN(n1033) );
  NAND2_X1 U1016 ( .A1(\mem[14][9] ), .A2(n1533), .ZN(n519) );
  OAI21_X1 U1017 ( .B1(n1616), .B2(n1534), .A(n520), .ZN(n1034) );
  NAND2_X1 U1018 ( .A1(\mem[14][10] ), .A2(n1533), .ZN(n520) );
  OAI21_X1 U1019 ( .B1(n1615), .B2(n1534), .A(n521), .ZN(n1035) );
  NAND2_X1 U1020 ( .A1(\mem[14][11] ), .A2(n1533), .ZN(n521) );
  OAI21_X1 U1021 ( .B1(n1614), .B2(n1534), .A(n522), .ZN(n1036) );
  NAND2_X1 U1022 ( .A1(\mem[14][12] ), .A2(n1533), .ZN(n522) );
  OAI21_X1 U1023 ( .B1(n1613), .B2(n1534), .A(n523), .ZN(n1037) );
  NAND2_X1 U1024 ( .A1(\mem[14][13] ), .A2(n1532), .ZN(n523) );
  OAI21_X1 U1025 ( .B1(n1612), .B2(n1534), .A(n524), .ZN(n1038) );
  NAND2_X1 U1026 ( .A1(\mem[14][14] ), .A2(n1533), .ZN(n524) );
  OAI21_X1 U1027 ( .B1(n1611), .B2(n1534), .A(n525), .ZN(n1039) );
  NAND2_X1 U1028 ( .A1(\mem[14][15] ), .A2(n1533), .ZN(n525) );
  OAI21_X1 U1029 ( .B1(n1610), .B2(n509), .A(n526), .ZN(n1040) );
  NAND2_X1 U1030 ( .A1(\mem[14][16] ), .A2(n1532), .ZN(n526) );
  OAI21_X1 U1031 ( .B1(n1609), .B2(n509), .A(n527), .ZN(n1041) );
  NAND2_X1 U1032 ( .A1(\mem[14][17] ), .A2(n1532), .ZN(n527) );
  OAI21_X1 U1033 ( .B1(n1608), .B2(n509), .A(n528), .ZN(n1042) );
  NAND2_X1 U1034 ( .A1(\mem[14][18] ), .A2(n1532), .ZN(n528) );
  OAI21_X1 U1035 ( .B1(n1607), .B2(n509), .A(n529), .ZN(n1043) );
  NAND2_X1 U1036 ( .A1(\mem[14][19] ), .A2(n1532), .ZN(n529) );
  OAI21_X1 U1037 ( .B1(n1606), .B2(n509), .A(n530), .ZN(n1044) );
  NAND2_X1 U1038 ( .A1(\mem[14][20] ), .A2(n1532), .ZN(n530) );
  OAI21_X1 U1039 ( .B1(n1605), .B2(n509), .A(n531), .ZN(n1045) );
  NAND2_X1 U1040 ( .A1(\mem[14][21] ), .A2(n1532), .ZN(n531) );
  OAI21_X1 U1041 ( .B1(n1604), .B2(n509), .A(n532), .ZN(n1046) );
  NAND2_X1 U1042 ( .A1(\mem[14][22] ), .A2(n1532), .ZN(n532) );
  OAI21_X1 U1043 ( .B1(n1603), .B2(n509), .A(n533), .ZN(n1047) );
  NAND2_X1 U1044 ( .A1(\mem[14][23] ), .A2(n1532), .ZN(n533) );
  OAI21_X1 U1045 ( .B1(n1602), .B2(n509), .A(n534), .ZN(n1048) );
  NAND2_X1 U1046 ( .A1(\mem[14][24] ), .A2(n1531), .ZN(n534) );
  OAI21_X1 U1047 ( .B1(n1601), .B2(n509), .A(n535), .ZN(n1049) );
  NAND2_X1 U1048 ( .A1(\mem[14][25] ), .A2(n1531), .ZN(n535) );
  OAI21_X1 U1049 ( .B1(n1600), .B2(n509), .A(n536), .ZN(n1050) );
  NAND2_X1 U1050 ( .A1(\mem[14][26] ), .A2(n1531), .ZN(n536) );
  OAI21_X1 U1051 ( .B1(n1595), .B2(n1533), .A(n541), .ZN(n1055) );
  NAND2_X1 U1052 ( .A1(\mem[14][31] ), .A2(n1531), .ZN(n541) );
  OAI21_X1 U1053 ( .B1(n1626), .B2(n1528), .A(n544), .ZN(n1056) );
  NAND2_X1 U1054 ( .A1(\mem[15][0] ), .A2(n1530), .ZN(n544) );
  OAI21_X1 U1055 ( .B1(n1625), .B2(n1527), .A(n545), .ZN(n1057) );
  NAND2_X1 U1056 ( .A1(\mem[15][1] ), .A2(n1530), .ZN(n545) );
  OAI21_X1 U1057 ( .B1(n1624), .B2(n1528), .A(n546), .ZN(n1058) );
  NAND2_X1 U1058 ( .A1(\mem[15][2] ), .A2(n1530), .ZN(n546) );
  OAI21_X1 U1059 ( .B1(n1623), .B2(n1527), .A(n547), .ZN(n1059) );
  NAND2_X1 U1060 ( .A1(\mem[15][3] ), .A2(n1528), .ZN(n547) );
  OAI21_X1 U1061 ( .B1(n1622), .B2(n1527), .A(n548), .ZN(n1060) );
  NAND2_X1 U1062 ( .A1(\mem[15][4] ), .A2(n1527), .ZN(n548) );
  OAI21_X1 U1063 ( .B1(n1621), .B2(n1528), .A(n549), .ZN(n1061) );
  NAND2_X1 U1064 ( .A1(\mem[15][5] ), .A2(n1528), .ZN(n549) );
  OAI21_X1 U1065 ( .B1(n1620), .B2(n1528), .A(n550), .ZN(n1062) );
  NAND2_X1 U1066 ( .A1(\mem[15][6] ), .A2(n1529), .ZN(n550) );
  OAI21_X1 U1067 ( .B1(n1619), .B2(n1528), .A(n551), .ZN(n1063) );
  NAND2_X1 U1068 ( .A1(\mem[15][7] ), .A2(n1527), .ZN(n551) );
  OAI21_X1 U1069 ( .B1(n1618), .B2(n1528), .A(n552), .ZN(n1064) );
  NAND2_X1 U1070 ( .A1(\mem[15][8] ), .A2(n1527), .ZN(n552) );
  OAI21_X1 U1071 ( .B1(n1617), .B2(n1528), .A(n553), .ZN(n1065) );
  NAND2_X1 U1072 ( .A1(\mem[15][9] ), .A2(n1527), .ZN(n553) );
  OAI21_X1 U1073 ( .B1(n1616), .B2(n1528), .A(n554), .ZN(n1066) );
  NAND2_X1 U1074 ( .A1(\mem[15][10] ), .A2(n1527), .ZN(n554) );
  OAI21_X1 U1075 ( .B1(n1615), .B2(n1528), .A(n555), .ZN(n1067) );
  NAND2_X1 U1076 ( .A1(\mem[15][11] ), .A2(n1527), .ZN(n555) );
  OAI21_X1 U1077 ( .B1(n1614), .B2(n1528), .A(n556), .ZN(n1068) );
  NAND2_X1 U1078 ( .A1(\mem[15][12] ), .A2(n1527), .ZN(n556) );
  OAI21_X1 U1079 ( .B1(n1613), .B2(n1528), .A(n557), .ZN(n1069) );
  NAND2_X1 U1080 ( .A1(\mem[15][13] ), .A2(n543), .ZN(n557) );
  OAI21_X1 U1081 ( .B1(n1612), .B2(n1528), .A(n558), .ZN(n1070) );
  NAND2_X1 U1082 ( .A1(\mem[15][14] ), .A2(n1527), .ZN(n558) );
  OAI21_X1 U1083 ( .B1(n1611), .B2(n1529), .A(n559), .ZN(n1071) );
  NAND2_X1 U1084 ( .A1(\mem[15][15] ), .A2(n1527), .ZN(n559) );
  OAI21_X1 U1085 ( .B1(n1610), .B2(n1529), .A(n560), .ZN(n1072) );
  NAND2_X1 U1086 ( .A1(\mem[15][16] ), .A2(n543), .ZN(n560) );
  OAI21_X1 U1087 ( .B1(n1609), .B2(n1529), .A(n561), .ZN(n1073) );
  NAND2_X1 U1088 ( .A1(\mem[15][17] ), .A2(n543), .ZN(n561) );
  OAI21_X1 U1089 ( .B1(n1608), .B2(n1529), .A(n562), .ZN(n1074) );
  NAND2_X1 U1090 ( .A1(\mem[15][18] ), .A2(n543), .ZN(n562) );
  OAI21_X1 U1091 ( .B1(n1607), .B2(n1529), .A(n563), .ZN(n1075) );
  NAND2_X1 U1092 ( .A1(\mem[15][19] ), .A2(n543), .ZN(n563) );
  OAI21_X1 U1093 ( .B1(n1606), .B2(n1529), .A(n564), .ZN(n1076) );
  NAND2_X1 U1094 ( .A1(\mem[15][20] ), .A2(n543), .ZN(n564) );
  OAI21_X1 U1095 ( .B1(n1605), .B2(n1529), .A(n565), .ZN(n1077) );
  NAND2_X1 U1096 ( .A1(\mem[15][21] ), .A2(n543), .ZN(n565) );
  OAI21_X1 U1097 ( .B1(n1604), .B2(n1529), .A(n566), .ZN(n1078) );
  NAND2_X1 U1098 ( .A1(\mem[15][22] ), .A2(n543), .ZN(n566) );
  OAI21_X1 U1099 ( .B1(n1603), .B2(n1529), .A(n567), .ZN(n1079) );
  NAND2_X1 U1100 ( .A1(\mem[15][23] ), .A2(n543), .ZN(n567) );
  OAI21_X1 U1101 ( .B1(n1602), .B2(n1529), .A(n568), .ZN(n1080) );
  NAND2_X1 U1102 ( .A1(\mem[15][24] ), .A2(n1529), .ZN(n568) );
  OAI21_X1 U1103 ( .B1(n1601), .B2(n1529), .A(n569), .ZN(n1081) );
  NAND2_X1 U1104 ( .A1(\mem[15][25] ), .A2(n543), .ZN(n569) );
  OAI21_X1 U1105 ( .B1(n1600), .B2(n1529), .A(n570), .ZN(n1082) );
  NAND2_X1 U1106 ( .A1(\mem[15][26] ), .A2(n543), .ZN(n570) );
  OAI21_X1 U1107 ( .B1(n1595), .B2(n1527), .A(n575), .ZN(n1087) );
  NAND2_X1 U1108 ( .A1(\mem[15][31] ), .A2(n543), .ZN(n575) );
  OAI21_X1 U1109 ( .B1(n1589), .B2(n1626), .A(n38), .ZN(n576) );
  NAND2_X1 U1110 ( .A1(\mem[0][0] ), .A2(n1587), .ZN(n38) );
  OAI21_X1 U1111 ( .B1(n1589), .B2(n1624), .A(n40), .ZN(n578) );
  NAND2_X1 U1112 ( .A1(\mem[0][2] ), .A2(n1587), .ZN(n40) );
  OAI21_X1 U1113 ( .B1(n1589), .B2(n1621), .A(n43), .ZN(n581) );
  NAND2_X1 U1114 ( .A1(\mem[0][5] ), .A2(n1588), .ZN(n43) );
  OAI21_X1 U1115 ( .B1(n1589), .B2(n1620), .A(n44), .ZN(n582) );
  NAND2_X1 U1116 ( .A1(\mem[0][6] ), .A2(n1588), .ZN(n44) );
  OAI21_X1 U1117 ( .B1(n1589), .B2(n1619), .A(n45), .ZN(n583) );
  NAND2_X1 U1118 ( .A1(\mem[0][7] ), .A2(n37), .ZN(n45) );
  OAI21_X1 U1119 ( .B1(n1589), .B2(n1618), .A(n46), .ZN(n584) );
  NAND2_X1 U1120 ( .A1(\mem[0][8] ), .A2(n37), .ZN(n46) );
  OAI21_X1 U1121 ( .B1(n1589), .B2(n1617), .A(n47), .ZN(n585) );
  NAND2_X1 U1122 ( .A1(\mem[0][9] ), .A2(n37), .ZN(n47) );
  OAI21_X1 U1123 ( .B1(n1589), .B2(n1616), .A(n48), .ZN(n586) );
  NAND2_X1 U1124 ( .A1(\mem[0][10] ), .A2(n37), .ZN(n48) );
  OAI21_X1 U1125 ( .B1(n1589), .B2(n1615), .A(n49), .ZN(n587) );
  NAND2_X1 U1126 ( .A1(\mem[0][11] ), .A2(n37), .ZN(n49) );
  OAI21_X1 U1127 ( .B1(n1589), .B2(n1614), .A(n50), .ZN(n588) );
  NAND2_X1 U1128 ( .A1(\mem[0][12] ), .A2(n37), .ZN(n50) );
  OAI21_X1 U1129 ( .B1(n1589), .B2(n1613), .A(n51), .ZN(n589) );
  NAND2_X1 U1130 ( .A1(\mem[0][13] ), .A2(n1588), .ZN(n51) );
  OAI21_X1 U1131 ( .B1(n1589), .B2(n1612), .A(n52), .ZN(n590) );
  NAND2_X1 U1132 ( .A1(\mem[0][14] ), .A2(n37), .ZN(n52) );
  OAI21_X1 U1133 ( .B1(n1589), .B2(n1611), .A(n53), .ZN(n591) );
  NAND2_X1 U1134 ( .A1(\mem[0][15] ), .A2(n37), .ZN(n53) );
  OAI21_X1 U1135 ( .B1(n1590), .B2(n1610), .A(n54), .ZN(n592) );
  NAND2_X1 U1136 ( .A1(\mem[0][16] ), .A2(n1588), .ZN(n54) );
  OAI21_X1 U1137 ( .B1(n1590), .B2(n1609), .A(n55), .ZN(n593) );
  NAND2_X1 U1138 ( .A1(\mem[0][17] ), .A2(n1588), .ZN(n55) );
  OAI21_X1 U1139 ( .B1(n1590), .B2(n1608), .A(n56), .ZN(n594) );
  NAND2_X1 U1140 ( .A1(\mem[0][18] ), .A2(n1588), .ZN(n56) );
  OAI21_X1 U1141 ( .B1(n1590), .B2(n1607), .A(n57), .ZN(n595) );
  NAND2_X1 U1142 ( .A1(\mem[0][19] ), .A2(n1588), .ZN(n57) );
  OAI21_X1 U1143 ( .B1(n1590), .B2(n1606), .A(n58), .ZN(n596) );
  NAND2_X1 U1144 ( .A1(\mem[0][20] ), .A2(n1588), .ZN(n58) );
  OAI21_X1 U1145 ( .B1(n1590), .B2(n1605), .A(n59), .ZN(n597) );
  NAND2_X1 U1146 ( .A1(\mem[0][21] ), .A2(n1588), .ZN(n59) );
  OAI21_X1 U1147 ( .B1(n1590), .B2(n1604), .A(n60), .ZN(n598) );
  NAND2_X1 U1148 ( .A1(\mem[0][22] ), .A2(n1588), .ZN(n60) );
  OAI21_X1 U1149 ( .B1(n1590), .B2(n1603), .A(n61), .ZN(n599) );
  NAND2_X1 U1150 ( .A1(\mem[0][23] ), .A2(n1588), .ZN(n61) );
  OAI21_X1 U1151 ( .B1(n1590), .B2(n1602), .A(n62), .ZN(n600) );
  NAND2_X1 U1152 ( .A1(\mem[0][24] ), .A2(n1587), .ZN(n62) );
  OAI21_X1 U1153 ( .B1(n1590), .B2(n1601), .A(n63), .ZN(n601) );
  NAND2_X1 U1154 ( .A1(\mem[0][25] ), .A2(n1587), .ZN(n63) );
  OAI21_X1 U1155 ( .B1(n1590), .B2(n1600), .A(n64), .ZN(n602) );
  NAND2_X1 U1156 ( .A1(\mem[0][26] ), .A2(n1587), .ZN(n64) );
  OAI21_X1 U1157 ( .B1(n1590), .B2(n1599), .A(n65), .ZN(n603) );
  NAND2_X1 U1158 ( .A1(\mem[0][27] ), .A2(n1587), .ZN(n65) );
  OAI21_X1 U1159 ( .B1(n1590), .B2(n1598), .A(n66), .ZN(n604) );
  NAND2_X1 U1160 ( .A1(\mem[0][28] ), .A2(n1587), .ZN(n66) );
  OAI21_X1 U1161 ( .B1(n1589), .B2(n1625), .A(n39), .ZN(n577) );
  NAND2_X1 U1162 ( .A1(\mem[0][1] ), .A2(n1587), .ZN(n39) );
  OAI21_X1 U1163 ( .B1(n1590), .B2(n1623), .A(n41), .ZN(n579) );
  NAND2_X1 U1164 ( .A1(\mem[0][3] ), .A2(n1587), .ZN(n41) );
  OAI21_X1 U1165 ( .B1(n37), .B2(n1622), .A(n42), .ZN(n580) );
  NAND2_X1 U1166 ( .A1(\mem[0][4] ), .A2(n1588), .ZN(n42) );
  OAI21_X1 U1167 ( .B1(n37), .B2(n1595), .A(n69), .ZN(n607) );
  NAND2_X1 U1168 ( .A1(\mem[0][31] ), .A2(n1587), .ZN(n69) );
  MUX2_X1 U1169 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n1511), .Z(n4) );
  MUX2_X1 U1170 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n1511), .Z(n5) );
  MUX2_X1 U1171 ( .A(n5), .B(n4), .S(n1506), .Z(n6) );
  MUX2_X1 U1172 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n1511), .Z(n7) );
  MUX2_X1 U1173 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n1511), .Z(n8) );
  MUX2_X1 U1174 ( .A(n8), .B(n7), .S(n1506), .Z(n9) );
  MUX2_X1 U1175 ( .A(n9), .B(n6), .S(n1503), .Z(n10) );
  MUX2_X1 U1176 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n1511), .Z(n11) );
  MUX2_X1 U1177 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n1511), .Z(n12) );
  MUX2_X1 U1178 ( .A(n12), .B(n11), .S(n1506), .Z(n13) );
  MUX2_X1 U1179 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n1511), .Z(n14) );
  MUX2_X1 U1180 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n1511), .Z(n15) );
  MUX2_X1 U1181 ( .A(n15), .B(n14), .S(n1506), .Z(n16) );
  MUX2_X1 U1182 ( .A(n16), .B(n13), .S(n1503), .Z(n17) );
  MUX2_X1 U1183 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n1513), .Z(n18) );
  MUX2_X1 U1184 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n1513), .Z(n19) );
  MUX2_X1 U1185 ( .A(n19), .B(n18), .S(n1506), .Z(n20) );
  MUX2_X1 U1186 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n1511), .Z(n21) );
  MUX2_X1 U1187 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n1511), .Z(n22) );
  MUX2_X1 U1188 ( .A(n22), .B(n21), .S(n1506), .Z(n23) );
  MUX2_X1 U1189 ( .A(n23), .B(n20), .S(n1503), .Z(n24) );
  MUX2_X1 U1190 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n1511), .Z(n25) );
  MUX2_X1 U1191 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n1511), .Z(n26) );
  MUX2_X1 U1192 ( .A(n26), .B(n25), .S(n1506), .Z(n27) );
  MUX2_X1 U1193 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n1511), .Z(n28) );
  MUX2_X1 U1194 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n1511), .Z(n29) );
  MUX2_X1 U1195 ( .A(n29), .B(n28), .S(n1506), .Z(n30) );
  MUX2_X1 U1196 ( .A(n30), .B(n27), .S(n1503), .Z(n31) );
  MUX2_X1 U1197 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n1512), .Z(n32) );
  MUX2_X1 U1198 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n1512), .Z(n33) );
  MUX2_X1 U1199 ( .A(n33), .B(n32), .S(n1506), .Z(n34) );
  MUX2_X1 U1200 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n1512), .Z(n35) );
  MUX2_X1 U1201 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n1512), .Z(n36) );
  MUX2_X1 U1202 ( .A(n36), .B(n35), .S(n1507), .Z(n1088) );
  MUX2_X1 U1203 ( .A(n1088), .B(n34), .S(n1504), .Z(n1089) );
  MUX2_X1 U1204 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n1512), .Z(n1090) );
  MUX2_X1 U1205 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n1512), .Z(n1091) );
  MUX2_X1 U1206 ( .A(n1091), .B(n1090), .S(n1506), .Z(n1092) );
  MUX2_X1 U1207 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n1512), .Z(n1093) );
  MUX2_X1 U1208 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n1512), .Z(n1094) );
  MUX2_X1 U1209 ( .A(n1094), .B(n1093), .S(n1508), .Z(n1095) );
  MUX2_X1 U1210 ( .A(n1095), .B(n1092), .S(n1505), .Z(n1096) );
  MUX2_X1 U1211 ( .A(n1096), .B(n1089), .S(N13), .Z(N43) );
  MUX2_X1 U1212 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n1512), .Z(n1097) );
  MUX2_X1 U1213 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n1512), .Z(n1098) );
  MUX2_X1 U1214 ( .A(n1098), .B(n1097), .S(n1507), .Z(n1099) );
  MUX2_X1 U1215 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n1512), .Z(n1100) );
  MUX2_X1 U1216 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n1512), .Z(n1101) );
  MUX2_X1 U1217 ( .A(n1101), .B(n1100), .S(n1507), .Z(n1102) );
  MUX2_X1 U1218 ( .A(n1102), .B(n1099), .S(n1503), .Z(n1103) );
  MUX2_X1 U1219 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n1513), .Z(n1104) );
  MUX2_X1 U1220 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n1513), .Z(n1105) );
  MUX2_X1 U1221 ( .A(n1105), .B(n1104), .S(n1506), .Z(n1106) );
  MUX2_X1 U1222 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n1513), .Z(n1107) );
  MUX2_X1 U1223 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n1513), .Z(n1108) );
  MUX2_X1 U1224 ( .A(n1108), .B(n1107), .S(n1508), .Z(n1109) );
  MUX2_X1 U1225 ( .A(n1109), .B(n1106), .S(n1505), .Z(n1110) );
  MUX2_X1 U1226 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n1513), .Z(n1111) );
  MUX2_X1 U1227 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n1513), .Z(n1112) );
  MUX2_X1 U1228 ( .A(n1112), .B(n1111), .S(n1508), .Z(n1113) );
  MUX2_X1 U1229 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n1513), .Z(n1114) );
  MUX2_X1 U1230 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n1513), .Z(n1115) );
  MUX2_X1 U1231 ( .A(n1115), .B(n1114), .S(n1508), .Z(n1116) );
  MUX2_X1 U1232 ( .A(n1116), .B(n1113), .S(n1505), .Z(n1117) );
  MUX2_X1 U1233 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n1513), .Z(n1118) );
  MUX2_X1 U1234 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n1513), .Z(n1119) );
  MUX2_X1 U1235 ( .A(n1119), .B(n1118), .S(n1507), .Z(n1120) );
  MUX2_X1 U1236 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n1513), .Z(n1121) );
  MUX2_X1 U1237 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n1513), .Z(n1122) );
  MUX2_X1 U1238 ( .A(n1122), .B(n1121), .S(n1506), .Z(n1123) );
  MUX2_X1 U1239 ( .A(n1123), .B(n1120), .S(n1504), .Z(n1124) );
  MUX2_X1 U1240 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n1513), .Z(n1125) );
  MUX2_X1 U1241 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n1515), .Z(n1126) );
  MUX2_X1 U1242 ( .A(n1126), .B(n1125), .S(n1510), .Z(n1127) );
  MUX2_X1 U1243 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n1524), .Z(n1128) );
  MUX2_X1 U1244 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n1514), .Z(n1129) );
  MUX2_X1 U1245 ( .A(n1129), .B(n1128), .S(n1510), .Z(n1130) );
  MUX2_X1 U1246 ( .A(n1130), .B(n1127), .S(n1504), .Z(n1131) );
  MUX2_X1 U1247 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n1513), .Z(n1132) );
  MUX2_X1 U1248 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(N10), .Z(n1133) );
  MUX2_X1 U1249 ( .A(n1133), .B(n1132), .S(n1510), .Z(n1134) );
  MUX2_X1 U1250 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(N10), .Z(n1135) );
  MUX2_X1 U1251 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n1511), .Z(n1136) );
  MUX2_X1 U1252 ( .A(n1136), .B(n1135), .S(n1510), .Z(n1137) );
  MUX2_X1 U1253 ( .A(n1137), .B(n1134), .S(n1503), .Z(n1138) );
  MUX2_X1 U1254 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n1512), .Z(n1139) );
  MUX2_X1 U1255 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n1524), .Z(n1140) );
  MUX2_X1 U1256 ( .A(n1140), .B(n1139), .S(n1507), .Z(n1141) );
  MUX2_X1 U1257 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n1526), .Z(n1142) );
  MUX2_X1 U1258 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(N10), .Z(n1143) );
  MUX2_X1 U1259 ( .A(n1143), .B(n1142), .S(n1510), .Z(n1144) );
  MUX2_X1 U1260 ( .A(n1144), .B(n1141), .S(n1503), .Z(n1145) );
  MUX2_X1 U1261 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n1526), .Z(n1146) );
  MUX2_X1 U1262 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n1511), .Z(n1147) );
  MUX2_X1 U1263 ( .A(n1147), .B(n1146), .S(n1510), .Z(n1148) );
  MUX2_X1 U1264 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n1525), .Z(n1149) );
  MUX2_X1 U1265 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(N10), .Z(n1150) );
  MUX2_X1 U1266 ( .A(n1150), .B(n1149), .S(n1506), .Z(n1151) );
  MUX2_X1 U1267 ( .A(n1151), .B(n1148), .S(n1503), .Z(n1152) );
  MUX2_X1 U1268 ( .A(n1152), .B(n1145), .S(N13), .Z(N39) );
  MUX2_X1 U1269 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n1526), .Z(n1153) );
  MUX2_X1 U1270 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n1514), .Z(n1154) );
  MUX2_X1 U1271 ( .A(n1154), .B(n1153), .S(n1510), .Z(n1155) );
  MUX2_X1 U1272 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n1515), .Z(n1156) );
  MUX2_X1 U1273 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(N10), .Z(n1157) );
  MUX2_X1 U1274 ( .A(n1157), .B(n1156), .S(n1510), .Z(n1158) );
  MUX2_X1 U1275 ( .A(n1158), .B(n1155), .S(n1503), .Z(n1159) );
  MUX2_X1 U1276 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n1513), .Z(n1160) );
  MUX2_X1 U1277 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n1517), .Z(n1161) );
  MUX2_X1 U1278 ( .A(n1161), .B(n1160), .S(n1510), .Z(n1162) );
  MUX2_X1 U1279 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n1526), .Z(n1163) );
  MUX2_X1 U1280 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n1517), .Z(n1164) );
  MUX2_X1 U1281 ( .A(n1164), .B(n1163), .S(n1510), .Z(n1165) );
  MUX2_X1 U1282 ( .A(n1165), .B(n1162), .S(n1505), .Z(n1166) );
  MUX2_X1 U1283 ( .A(\mem[14][8] ), .B(\mem[15][8] ), .S(n1512), .Z(n1167) );
  MUX2_X1 U1284 ( .A(\mem[12][8] ), .B(\mem[13][8] ), .S(n1524), .Z(n1168) );
  MUX2_X1 U1285 ( .A(n1168), .B(n1167), .S(n1507), .Z(n1169) );
  MUX2_X1 U1286 ( .A(\mem[10][8] ), .B(\mem[11][8] ), .S(n1524), .Z(n1170) );
  MUX2_X1 U1287 ( .A(\mem[8][8] ), .B(\mem[9][8] ), .S(N10), .Z(n1171) );
  MUX2_X1 U1288 ( .A(n1171), .B(n1170), .S(n1507), .Z(n1172) );
  MUX2_X1 U1289 ( .A(n1172), .B(n1169), .S(n1504), .Z(n1173) );
  MUX2_X1 U1290 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n1524), .Z(n1174) );
  MUX2_X1 U1291 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n1524), .Z(n1175) );
  MUX2_X1 U1292 ( .A(n1175), .B(n1174), .S(n1507), .Z(n1176) );
  MUX2_X1 U1293 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n1526), .Z(n1177) );
  MUX2_X1 U1294 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(N10), .Z(n1178) );
  MUX2_X1 U1295 ( .A(n1178), .B(n1177), .S(n1507), .Z(n1179) );
  MUX2_X1 U1296 ( .A(n1179), .B(n1176), .S(n1504), .Z(n1180) );
  MUX2_X1 U1297 ( .A(n1180), .B(n1173), .S(N13), .Z(N37) );
  MUX2_X1 U1298 ( .A(\mem[14][9] ), .B(\mem[15][9] ), .S(n1517), .Z(n1181) );
  MUX2_X1 U1299 ( .A(\mem[12][9] ), .B(\mem[13][9] ), .S(n1515), .Z(n1182) );
  MUX2_X1 U1300 ( .A(n1182), .B(n1181), .S(n1507), .Z(n1183) );
  MUX2_X1 U1301 ( .A(\mem[10][9] ), .B(\mem[11][9] ), .S(n1524), .Z(n1184) );
  MUX2_X1 U1302 ( .A(\mem[8][9] ), .B(\mem[9][9] ), .S(n1514), .Z(n1185) );
  MUX2_X1 U1303 ( .A(n1185), .B(n1184), .S(n1507), .Z(n1186) );
  MUX2_X1 U1304 ( .A(n1186), .B(n1183), .S(n1503), .Z(n1187) );
  MUX2_X1 U1305 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n1524), .Z(n1188) );
  MUX2_X1 U1306 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n1524), .Z(n1189) );
  MUX2_X1 U1307 ( .A(n1189), .B(n1188), .S(n1507), .Z(n1190) );
  MUX2_X1 U1308 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n1516), .Z(n1191) );
  MUX2_X1 U1309 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n1524), .Z(n1192) );
  MUX2_X1 U1310 ( .A(n1192), .B(n1191), .S(n1507), .Z(n1193) );
  MUX2_X1 U1311 ( .A(n1193), .B(n1190), .S(n1505), .Z(n1194) );
  MUX2_X1 U1312 ( .A(\mem[14][10] ), .B(\mem[15][10] ), .S(N10), .Z(n1195) );
  MUX2_X1 U1313 ( .A(\mem[12][10] ), .B(\mem[13][10] ), .S(N10), .Z(n1196) );
  MUX2_X1 U1314 ( .A(n1196), .B(n1195), .S(n1507), .Z(n1197) );
  MUX2_X1 U1315 ( .A(\mem[10][10] ), .B(\mem[11][10] ), .S(N10), .Z(n1198) );
  MUX2_X1 U1316 ( .A(\mem[8][10] ), .B(\mem[9][10] ), .S(N10), .Z(n1199) );
  MUX2_X1 U1317 ( .A(n1199), .B(n1198), .S(n1507), .Z(n1200) );
  MUX2_X1 U1318 ( .A(n1200), .B(n1197), .S(n1505), .Z(n1201) );
  MUX2_X1 U1319 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n1513), .Z(n1202) );
  MUX2_X1 U1320 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n1525), .Z(n1203) );
  MUX2_X1 U1321 ( .A(n1203), .B(n1202), .S(n1507), .Z(n1204) );
  MUX2_X1 U1322 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n1525), .Z(n1205) );
  MUX2_X1 U1323 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(N10), .Z(n1206) );
  MUX2_X1 U1324 ( .A(n1206), .B(n1205), .S(n1507), .Z(n1207) );
  MUX2_X1 U1325 ( .A(n1207), .B(n1204), .S(n1503), .Z(n1208) );
  MUX2_X1 U1326 ( .A(\mem[14][11] ), .B(\mem[15][11] ), .S(n1514), .Z(n1209)
         );
  MUX2_X1 U1327 ( .A(\mem[12][11] ), .B(\mem[13][11] ), .S(n1525), .Z(n1210)
         );
  MUX2_X1 U1328 ( .A(n1210), .B(n1209), .S(n1506), .Z(n1211) );
  MUX2_X1 U1329 ( .A(\mem[10][11] ), .B(\mem[11][11] ), .S(n1524), .Z(n1212)
         );
  MUX2_X1 U1330 ( .A(\mem[8][11] ), .B(\mem[9][11] ), .S(N10), .Z(n1213) );
  MUX2_X1 U1331 ( .A(n1213), .B(n1212), .S(n1510), .Z(n1214) );
  MUX2_X1 U1332 ( .A(n1214), .B(n1211), .S(n1504), .Z(n1215) );
  MUX2_X1 U1333 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n1513), .Z(n1216) );
  MUX2_X1 U1334 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n1526), .Z(n1217) );
  MUX2_X1 U1335 ( .A(n1217), .B(n1216), .S(n1509), .Z(n1218) );
  MUX2_X1 U1336 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n1515), .Z(n1219) );
  MUX2_X1 U1337 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n1511), .Z(n1220) );
  MUX2_X1 U1338 ( .A(n1220), .B(n1219), .S(n1509), .Z(n1221) );
  MUX2_X1 U1339 ( .A(n1221), .B(n1218), .S(n1505), .Z(n1222) );
  MUX2_X1 U1340 ( .A(\mem[14][12] ), .B(\mem[15][12] ), .S(n1515), .Z(n1223)
         );
  MUX2_X1 U1341 ( .A(\mem[12][12] ), .B(\mem[13][12] ), .S(n1526), .Z(n1224)
         );
  MUX2_X1 U1342 ( .A(n1224), .B(n1223), .S(n1508), .Z(n1225) );
  MUX2_X1 U1343 ( .A(\mem[10][12] ), .B(\mem[11][12] ), .S(n1517), .Z(n1226)
         );
  MUX2_X1 U1344 ( .A(\mem[8][12] ), .B(\mem[9][12] ), .S(n1524), .Z(n1227) );
  MUX2_X1 U1345 ( .A(n1227), .B(n1226), .S(n1508), .Z(n1228) );
  MUX2_X1 U1346 ( .A(n1228), .B(n1225), .S(n1505), .Z(n1229) );
  MUX2_X1 U1347 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n1511), .Z(n1230) );
  MUX2_X1 U1348 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n1512), .Z(n1231) );
  MUX2_X1 U1349 ( .A(n1231), .B(n1230), .S(n1509), .Z(n1232) );
  MUX2_X1 U1350 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n1514), .Z(n1233) );
  MUX2_X1 U1351 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n1525), .Z(n1234) );
  MUX2_X1 U1352 ( .A(n1234), .B(n1233), .S(n1509), .Z(n1235) );
  MUX2_X1 U1353 ( .A(n1235), .B(n1232), .S(n1504), .Z(n1236) );
  MUX2_X1 U1354 ( .A(\mem[14][13] ), .B(\mem[15][13] ), .S(n1524), .Z(n1237)
         );
  MUX2_X1 U1355 ( .A(\mem[12][13] ), .B(\mem[13][13] ), .S(N10), .Z(n1238) );
  MUX2_X1 U1356 ( .A(n1238), .B(n1237), .S(n1506), .Z(n1239) );
  MUX2_X1 U1357 ( .A(\mem[10][13] ), .B(\mem[11][13] ), .S(N10), .Z(n1240) );
  MUX2_X1 U1358 ( .A(\mem[8][13] ), .B(\mem[9][13] ), .S(N10), .Z(n1241) );
  MUX2_X1 U1359 ( .A(n1241), .B(n1240), .S(n1507), .Z(n1242) );
  MUX2_X1 U1360 ( .A(n1242), .B(n1239), .S(n1503), .Z(n1243) );
  MUX2_X1 U1361 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n1517), .Z(n1244) );
  MUX2_X1 U1362 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n1511), .Z(n1245) );
  MUX2_X1 U1363 ( .A(n1245), .B(n1244), .S(n1509), .Z(n1246) );
  MUX2_X1 U1364 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n1516), .Z(n1247) );
  MUX2_X1 U1365 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n1526), .Z(n1248) );
  MUX2_X1 U1366 ( .A(n1248), .B(n1247), .S(n1509), .Z(n1249) );
  MUX2_X1 U1367 ( .A(n1249), .B(n1246), .S(n1504), .Z(n1250) );
  MUX2_X1 U1368 ( .A(\mem[14][14] ), .B(\mem[15][14] ), .S(n1525), .Z(n1251)
         );
  MUX2_X1 U1369 ( .A(\mem[12][14] ), .B(\mem[13][14] ), .S(n1524), .Z(n1252)
         );
  MUX2_X1 U1370 ( .A(n1252), .B(n1251), .S(n1508), .Z(n1253) );
  MUX2_X1 U1371 ( .A(\mem[10][14] ), .B(\mem[11][14] ), .S(n1524), .Z(n1254)
         );
  MUX2_X1 U1372 ( .A(\mem[8][14] ), .B(\mem[9][14] ), .S(n1524), .Z(n1255) );
  MUX2_X1 U1373 ( .A(n1255), .B(n1254), .S(n1508), .Z(n1256) );
  MUX2_X1 U1374 ( .A(n1256), .B(n1253), .S(n1504), .Z(n1257) );
  MUX2_X1 U1375 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n1511), .Z(n1258) );
  MUX2_X1 U1376 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n1511), .Z(n1259) );
  MUX2_X1 U1377 ( .A(n1259), .B(n1258), .S(n1509), .Z(n1260) );
  MUX2_X1 U1378 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n1512), .Z(n1261) );
  MUX2_X1 U1379 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n1511), .Z(n1262) );
  MUX2_X1 U1380 ( .A(n1262), .B(n1261), .S(n1509), .Z(n1263) );
  MUX2_X1 U1381 ( .A(n1263), .B(n1260), .S(n1503), .Z(n1264) );
  MUX2_X1 U1382 ( .A(\mem[14][15] ), .B(\mem[15][15] ), .S(n1525), .Z(n1265)
         );
  MUX2_X1 U1383 ( .A(\mem[12][15] ), .B(\mem[13][15] ), .S(n1524), .Z(n1266)
         );
  MUX2_X1 U1384 ( .A(n1266), .B(n1265), .S(n1510), .Z(n1267) );
  MUX2_X1 U1385 ( .A(\mem[10][15] ), .B(\mem[11][15] ), .S(n1524), .Z(n1268)
         );
  MUX2_X1 U1386 ( .A(\mem[8][15] ), .B(\mem[9][15] ), .S(n1524), .Z(n1269) );
  MUX2_X1 U1387 ( .A(n1269), .B(n1268), .S(n1506), .Z(n1270) );
  MUX2_X1 U1388 ( .A(n1270), .B(n1267), .S(n1505), .Z(n1271) );
  MUX2_X1 U1389 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n1513), .Z(n1272) );
  MUX2_X1 U1390 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n1513), .Z(n1273) );
  MUX2_X1 U1391 ( .A(n1273), .B(n1272), .S(n1508), .Z(n1274) );
  MUX2_X1 U1392 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(n1512), .Z(n1275) );
  MUX2_X1 U1393 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(n1512), .Z(n1276) );
  MUX2_X1 U1394 ( .A(n1276), .B(n1275), .S(n1508), .Z(n1277) );
  MUX2_X1 U1395 ( .A(n1277), .B(n1274), .S(n1503), .Z(n1278) );
  MUX2_X1 U1396 ( .A(\mem[14][16] ), .B(\mem[15][16] ), .S(n1512), .Z(n1279)
         );
  MUX2_X1 U1397 ( .A(\mem[12][16] ), .B(\mem[13][16] ), .S(n1513), .Z(n1280)
         );
  MUX2_X1 U1398 ( .A(n1280), .B(n1279), .S(n1506), .Z(n1281) );
  MUX2_X1 U1399 ( .A(\mem[10][16] ), .B(\mem[11][16] ), .S(n1512), .Z(n1282)
         );
  MUX2_X1 U1400 ( .A(\mem[8][16] ), .B(\mem[9][16] ), .S(n1512), .Z(n1283) );
  MUX2_X1 U1401 ( .A(n1283), .B(n1282), .S(n1506), .Z(n1284) );
  MUX2_X1 U1402 ( .A(n1284), .B(n1281), .S(n1503), .Z(n1285) );
  MUX2_X1 U1403 ( .A(\mem[6][16] ), .B(\mem[7][16] ), .S(n1512), .Z(n1286) );
  MUX2_X1 U1404 ( .A(\mem[4][16] ), .B(\mem[5][16] ), .S(n1513), .Z(n1287) );
  MUX2_X1 U1405 ( .A(n1287), .B(n1286), .S(n1506), .Z(n1288) );
  MUX2_X1 U1406 ( .A(\mem[2][16] ), .B(\mem[3][16] ), .S(n1512), .Z(n1289) );
  MUX2_X1 U1407 ( .A(\mem[0][16] ), .B(\mem[1][16] ), .S(n1511), .Z(n1290) );
  MUX2_X1 U1408 ( .A(n1290), .B(n1289), .S(n1510), .Z(n1291) );
  MUX2_X1 U1409 ( .A(n1291), .B(n1288), .S(n1503), .Z(n1292) );
  MUX2_X1 U1410 ( .A(n1292), .B(n1285), .S(N13), .Z(N29) );
  MUX2_X1 U1411 ( .A(\mem[14][17] ), .B(\mem[15][17] ), .S(n1514), .Z(n1293)
         );
  MUX2_X1 U1412 ( .A(\mem[12][17] ), .B(\mem[13][17] ), .S(n1514), .Z(n1294)
         );
  MUX2_X1 U1413 ( .A(n1294), .B(n1293), .S(n1508), .Z(n1295) );
  MUX2_X1 U1414 ( .A(\mem[10][17] ), .B(\mem[11][17] ), .S(n1514), .Z(n1296)
         );
  MUX2_X1 U1415 ( .A(\mem[8][17] ), .B(\mem[9][17] ), .S(n1514), .Z(n1297) );
  MUX2_X1 U1416 ( .A(n1297), .B(n1296), .S(n1508), .Z(n1298) );
  MUX2_X1 U1417 ( .A(n1298), .B(n1295), .S(n1504), .Z(n1299) );
  MUX2_X1 U1418 ( .A(\mem[6][17] ), .B(\mem[7][17] ), .S(n1514), .Z(n1300) );
  MUX2_X1 U1419 ( .A(\mem[4][17] ), .B(\mem[5][17] ), .S(n1514), .Z(n1301) );
  MUX2_X1 U1420 ( .A(n1301), .B(n1300), .S(n1508), .Z(n1302) );
  MUX2_X1 U1421 ( .A(\mem[2][17] ), .B(\mem[3][17] ), .S(n1514), .Z(n1303) );
  MUX2_X1 U1422 ( .A(\mem[0][17] ), .B(\mem[1][17] ), .S(n1514), .Z(n1304) );
  MUX2_X1 U1423 ( .A(n1304), .B(n1303), .S(n1508), .Z(n1305) );
  MUX2_X1 U1424 ( .A(n1305), .B(n1302), .S(n1503), .Z(n1306) );
  MUX2_X1 U1425 ( .A(\mem[14][18] ), .B(\mem[15][18] ), .S(n1514), .Z(n1307)
         );
  MUX2_X1 U1426 ( .A(\mem[12][18] ), .B(\mem[13][18] ), .S(n1514), .Z(n1308)
         );
  MUX2_X1 U1427 ( .A(n1308), .B(n1307), .S(n1508), .Z(n1309) );
  MUX2_X1 U1428 ( .A(\mem[10][18] ), .B(\mem[11][18] ), .S(n1514), .Z(n1310)
         );
  MUX2_X1 U1429 ( .A(\mem[8][18] ), .B(\mem[9][18] ), .S(n1514), .Z(n1311) );
  MUX2_X1 U1430 ( .A(n1311), .B(n1310), .S(n1508), .Z(n1312) );
  MUX2_X1 U1431 ( .A(n1312), .B(n1309), .S(n1505), .Z(n1313) );
  MUX2_X1 U1432 ( .A(\mem[6][18] ), .B(\mem[7][18] ), .S(n1515), .Z(n1314) );
  MUX2_X1 U1433 ( .A(\mem[4][18] ), .B(\mem[5][18] ), .S(n1515), .Z(n1315) );
  MUX2_X1 U1434 ( .A(n1315), .B(n1314), .S(n1508), .Z(n1316) );
  MUX2_X1 U1435 ( .A(\mem[2][18] ), .B(\mem[3][18] ), .S(n1515), .Z(n1317) );
  MUX2_X1 U1436 ( .A(\mem[0][18] ), .B(\mem[1][18] ), .S(n1515), .Z(n1318) );
  MUX2_X1 U1437 ( .A(n1318), .B(n1317), .S(n1508), .Z(n1319) );
  MUX2_X1 U1438 ( .A(n1319), .B(n1316), .S(n1503), .Z(n1320) );
  MUX2_X1 U1439 ( .A(\mem[14][19] ), .B(\mem[15][19] ), .S(n1515), .Z(n1321)
         );
  MUX2_X1 U1440 ( .A(\mem[12][19] ), .B(\mem[13][19] ), .S(n1515), .Z(n1322)
         );
  MUX2_X1 U1441 ( .A(n1322), .B(n1321), .S(n1508), .Z(n1323) );
  MUX2_X1 U1442 ( .A(\mem[10][19] ), .B(\mem[11][19] ), .S(n1515), .Z(n1324)
         );
  MUX2_X1 U1443 ( .A(\mem[8][19] ), .B(\mem[9][19] ), .S(n1515), .Z(n1325) );
  MUX2_X1 U1444 ( .A(n1325), .B(n1324), .S(n1508), .Z(n1326) );
  MUX2_X1 U1445 ( .A(n1326), .B(n1323), .S(n1503), .Z(n1327) );
  MUX2_X1 U1446 ( .A(\mem[6][19] ), .B(\mem[7][19] ), .S(n1515), .Z(n1328) );
  MUX2_X1 U1447 ( .A(\mem[4][19] ), .B(\mem[5][19] ), .S(n1515), .Z(n1329) );
  MUX2_X1 U1448 ( .A(n1329), .B(n1328), .S(n1508), .Z(n1330) );
  MUX2_X1 U1449 ( .A(\mem[2][19] ), .B(\mem[3][19] ), .S(n1515), .Z(n1331) );
  MUX2_X1 U1450 ( .A(\mem[0][19] ), .B(\mem[1][19] ), .S(n1515), .Z(n1332) );
  MUX2_X1 U1451 ( .A(n1332), .B(n1331), .S(n1508), .Z(n1333) );
  MUX2_X1 U1452 ( .A(n1333), .B(n1330), .S(n1503), .Z(n1334) );
  MUX2_X1 U1453 ( .A(\mem[14][20] ), .B(\mem[15][20] ), .S(n1516), .Z(n1335)
         );
  MUX2_X1 U1454 ( .A(\mem[12][20] ), .B(\mem[13][20] ), .S(n1516), .Z(n1336)
         );
  MUX2_X1 U1455 ( .A(n1336), .B(n1335), .S(n1509), .Z(n1337) );
  MUX2_X1 U1456 ( .A(\mem[10][20] ), .B(\mem[11][20] ), .S(n1516), .Z(n1338)
         );
  MUX2_X1 U1457 ( .A(\mem[8][20] ), .B(\mem[9][20] ), .S(n1516), .Z(n1339) );
  MUX2_X1 U1458 ( .A(n1339), .B(n1338), .S(n1509), .Z(n1340) );
  MUX2_X1 U1459 ( .A(n1340), .B(n1337), .S(n1504), .Z(n1341) );
  MUX2_X1 U1460 ( .A(\mem[6][20] ), .B(\mem[7][20] ), .S(n1516), .Z(n1342) );
  MUX2_X1 U1461 ( .A(\mem[4][20] ), .B(\mem[5][20] ), .S(n1516), .Z(n1343) );
  MUX2_X1 U1462 ( .A(n1343), .B(n1342), .S(n1509), .Z(n1344) );
  MUX2_X1 U1463 ( .A(\mem[2][20] ), .B(\mem[3][20] ), .S(n1516), .Z(n1345) );
  MUX2_X1 U1464 ( .A(\mem[0][20] ), .B(\mem[1][20] ), .S(n1516), .Z(n1346) );
  MUX2_X1 U1465 ( .A(n1346), .B(n1345), .S(n1509), .Z(n1347) );
  MUX2_X1 U1466 ( .A(n1347), .B(n1344), .S(n1504), .Z(n1348) );
  MUX2_X1 U1467 ( .A(n1348), .B(n1341), .S(N13), .Z(N25) );
  MUX2_X1 U1468 ( .A(\mem[14][21] ), .B(\mem[15][21] ), .S(n1516), .Z(n1349)
         );
  MUX2_X1 U1469 ( .A(\mem[12][21] ), .B(\mem[13][21] ), .S(n1516), .Z(n1350)
         );
  MUX2_X1 U1470 ( .A(n1350), .B(n1349), .S(n1509), .Z(n1351) );
  MUX2_X1 U1471 ( .A(\mem[10][21] ), .B(\mem[11][21] ), .S(n1516), .Z(n1352)
         );
  MUX2_X1 U1472 ( .A(\mem[8][21] ), .B(\mem[9][21] ), .S(n1516), .Z(n1353) );
  MUX2_X1 U1473 ( .A(n1353), .B(n1352), .S(n1509), .Z(n1354) );
  MUX2_X1 U1474 ( .A(n1354), .B(n1351), .S(n1504), .Z(n1355) );
  MUX2_X1 U1475 ( .A(\mem[6][21] ), .B(\mem[7][21] ), .S(n1517), .Z(n1356) );
  MUX2_X1 U1476 ( .A(\mem[4][21] ), .B(\mem[5][21] ), .S(n1517), .Z(n1357) );
  MUX2_X1 U1477 ( .A(n1357), .B(n1356), .S(n1509), .Z(n1358) );
  MUX2_X1 U1478 ( .A(\mem[2][21] ), .B(\mem[3][21] ), .S(n1517), .Z(n1359) );
  MUX2_X1 U1479 ( .A(\mem[0][21] ), .B(\mem[1][21] ), .S(n1517), .Z(n1360) );
  MUX2_X1 U1480 ( .A(n1360), .B(n1359), .S(n1509), .Z(n1361) );
  MUX2_X1 U1481 ( .A(n1361), .B(n1358), .S(n1504), .Z(n1362) );
  MUX2_X1 U1482 ( .A(\mem[14][22] ), .B(\mem[15][22] ), .S(n1517), .Z(n1363)
         );
  MUX2_X1 U1483 ( .A(\mem[12][22] ), .B(\mem[13][22] ), .S(n1517), .Z(n1364)
         );
  MUX2_X1 U1484 ( .A(n1364), .B(n1363), .S(n1509), .Z(n1365) );
  MUX2_X1 U1485 ( .A(\mem[10][22] ), .B(\mem[11][22] ), .S(n1517), .Z(n1366)
         );
  MUX2_X1 U1486 ( .A(\mem[8][22] ), .B(\mem[9][22] ), .S(n1517), .Z(n1367) );
  MUX2_X1 U1487 ( .A(n1367), .B(n1366), .S(n1509), .Z(n1368) );
  MUX2_X1 U1488 ( .A(n1368), .B(n1365), .S(n1504), .Z(n1369) );
  MUX2_X1 U1489 ( .A(\mem[6][22] ), .B(\mem[7][22] ), .S(n1517), .Z(n1370) );
  MUX2_X1 U1490 ( .A(\mem[4][22] ), .B(\mem[5][22] ), .S(n1517), .Z(n1371) );
  MUX2_X1 U1491 ( .A(n1371), .B(n1370), .S(n1509), .Z(n1372) );
  MUX2_X1 U1492 ( .A(\mem[2][22] ), .B(\mem[3][22] ), .S(n1517), .Z(n1373) );
  MUX2_X1 U1493 ( .A(\mem[0][22] ), .B(\mem[1][22] ), .S(n1517), .Z(n1374) );
  MUX2_X1 U1494 ( .A(n1374), .B(n1373), .S(n1509), .Z(n1375) );
  MUX2_X1 U1495 ( .A(n1375), .B(n1372), .S(n1504), .Z(n1376) );
  MUX2_X1 U1496 ( .A(\mem[14][23] ), .B(\mem[15][23] ), .S(n1518), .Z(n1377)
         );
  MUX2_X1 U1497 ( .A(\mem[12][23] ), .B(\mem[13][23] ), .S(n1518), .Z(n1378)
         );
  MUX2_X1 U1498 ( .A(n1378), .B(n1377), .S(N11), .Z(n1379) );
  MUX2_X1 U1499 ( .A(\mem[10][23] ), .B(\mem[11][23] ), .S(n1518), .Z(n1380)
         );
  MUX2_X1 U1500 ( .A(\mem[8][23] ), .B(\mem[9][23] ), .S(n1518), .Z(n1381) );
  MUX2_X1 U1501 ( .A(n1381), .B(n1380), .S(N11), .Z(n1382) );
  MUX2_X1 U1502 ( .A(n1382), .B(n1379), .S(n1504), .Z(n1383) );
  MUX2_X1 U1503 ( .A(\mem[6][23] ), .B(\mem[7][23] ), .S(n1518), .Z(n1384) );
  MUX2_X1 U1504 ( .A(\mem[4][23] ), .B(\mem[5][23] ), .S(n1518), .Z(n1385) );
  MUX2_X1 U1505 ( .A(n1385), .B(n1384), .S(n1509), .Z(n1386) );
  MUX2_X1 U1506 ( .A(\mem[2][23] ), .B(\mem[3][23] ), .S(n1518), .Z(n1387) );
  MUX2_X1 U1507 ( .A(\mem[0][23] ), .B(\mem[1][23] ), .S(n1518), .Z(n1388) );
  MUX2_X1 U1508 ( .A(n1388), .B(n1387), .S(N11), .Z(n1389) );
  MUX2_X1 U1509 ( .A(n1389), .B(n1386), .S(n1504), .Z(n1390) );
  MUX2_X1 U1510 ( .A(\mem[14][24] ), .B(\mem[15][24] ), .S(n1518), .Z(n1391)
         );
  MUX2_X1 U1511 ( .A(\mem[12][24] ), .B(\mem[13][24] ), .S(n1518), .Z(n1392)
         );
  MUX2_X1 U1512 ( .A(n1392), .B(n1391), .S(n1510), .Z(n1393) );
  MUX2_X1 U1513 ( .A(\mem[10][24] ), .B(\mem[11][24] ), .S(n1518), .Z(n1394)
         );
  MUX2_X1 U1514 ( .A(\mem[8][24] ), .B(\mem[9][24] ), .S(n1518), .Z(n1395) );
  MUX2_X1 U1515 ( .A(n1395), .B(n1394), .S(n1506), .Z(n1396) );
  MUX2_X1 U1516 ( .A(n1396), .B(n1393), .S(n1504), .Z(n1397) );
  MUX2_X1 U1517 ( .A(\mem[6][24] ), .B(\mem[7][24] ), .S(n1519), .Z(n1398) );
  MUX2_X1 U1518 ( .A(\mem[4][24] ), .B(\mem[5][24] ), .S(n1519), .Z(n1399) );
  MUX2_X1 U1519 ( .A(n1399), .B(n1398), .S(n1507), .Z(n1400) );
  MUX2_X1 U1520 ( .A(\mem[2][24] ), .B(\mem[3][24] ), .S(n1519), .Z(n1401) );
  MUX2_X1 U1521 ( .A(\mem[0][24] ), .B(\mem[1][24] ), .S(n1519), .Z(n1402) );
  MUX2_X1 U1522 ( .A(n1402), .B(n1401), .S(N11), .Z(n1403) );
  MUX2_X1 U1523 ( .A(n1403), .B(n1400), .S(n1504), .Z(n1404) );
  MUX2_X1 U1524 ( .A(n1404), .B(n1397), .S(N13), .Z(N21) );
  MUX2_X1 U1525 ( .A(\mem[14][25] ), .B(\mem[15][25] ), .S(n1519), .Z(n1405)
         );
  MUX2_X1 U1526 ( .A(\mem[12][25] ), .B(\mem[13][25] ), .S(n1519), .Z(n1406)
         );
  MUX2_X1 U1527 ( .A(n1406), .B(n1405), .S(N11), .Z(n1407) );
  MUX2_X1 U1528 ( .A(\mem[10][25] ), .B(\mem[11][25] ), .S(n1519), .Z(n1408)
         );
  MUX2_X1 U1529 ( .A(\mem[8][25] ), .B(\mem[9][25] ), .S(n1519), .Z(n1409) );
  MUX2_X1 U1530 ( .A(n1409), .B(n1408), .S(n1507), .Z(n1410) );
  MUX2_X1 U1531 ( .A(n1410), .B(n1407), .S(n1504), .Z(n1411) );
  MUX2_X1 U1532 ( .A(\mem[6][25] ), .B(\mem[7][25] ), .S(n1519), .Z(n1412) );
  MUX2_X1 U1533 ( .A(\mem[4][25] ), .B(\mem[5][25] ), .S(n1519), .Z(n1413) );
  MUX2_X1 U1534 ( .A(n1413), .B(n1412), .S(N11), .Z(n1414) );
  MUX2_X1 U1535 ( .A(\mem[2][25] ), .B(\mem[3][25] ), .S(n1519), .Z(n1415) );
  MUX2_X1 U1536 ( .A(\mem[0][25] ), .B(\mem[1][25] ), .S(n1519), .Z(n1416) );
  MUX2_X1 U1537 ( .A(n1416), .B(n1415), .S(N11), .Z(n1417) );
  MUX2_X1 U1538 ( .A(n1417), .B(n1414), .S(n1504), .Z(n1418) );
  MUX2_X1 U1539 ( .A(\mem[14][26] ), .B(\mem[15][26] ), .S(n1520), .Z(n1419)
         );
  MUX2_X1 U1540 ( .A(\mem[12][26] ), .B(\mem[13][26] ), .S(n1520), .Z(n1420)
         );
  MUX2_X1 U1541 ( .A(n1420), .B(n1419), .S(n1507), .Z(n1421) );
  MUX2_X1 U1542 ( .A(\mem[10][26] ), .B(\mem[11][26] ), .S(n1520), .Z(n1422)
         );
  MUX2_X1 U1543 ( .A(\mem[8][26] ), .B(\mem[9][26] ), .S(n1520), .Z(n1423) );
  MUX2_X1 U1544 ( .A(n1423), .B(n1422), .S(N11), .Z(n1424) );
  MUX2_X1 U1545 ( .A(n1424), .B(n1421), .S(n1505), .Z(n1425) );
  MUX2_X1 U1546 ( .A(\mem[6][26] ), .B(\mem[7][26] ), .S(n1520), .Z(n1426) );
  MUX2_X1 U1547 ( .A(\mem[4][26] ), .B(\mem[5][26] ), .S(n1520), .Z(n1427) );
  MUX2_X1 U1548 ( .A(n1427), .B(n1426), .S(n1510), .Z(n1428) );
  MUX2_X1 U1549 ( .A(\mem[2][26] ), .B(\mem[3][26] ), .S(n1520), .Z(n1429) );
  MUX2_X1 U1550 ( .A(\mem[0][26] ), .B(\mem[1][26] ), .S(n1520), .Z(n1430) );
  MUX2_X1 U1551 ( .A(n1430), .B(n1429), .S(N11), .Z(n1431) );
  MUX2_X1 U1552 ( .A(n1431), .B(n1428), .S(n1505), .Z(n1432) );
  MUX2_X1 U1553 ( .A(n1432), .B(n1425), .S(N13), .Z(N19) );
  MUX2_X1 U1554 ( .A(\mem[14][27] ), .B(\mem[15][27] ), .S(n1520), .Z(n1433)
         );
  MUX2_X1 U1555 ( .A(\mem[12][27] ), .B(\mem[13][27] ), .S(n1520), .Z(n1434)
         );
  MUX2_X1 U1556 ( .A(n1434), .B(n1433), .S(N11), .Z(n1435) );
  MUX2_X1 U1557 ( .A(\mem[10][27] ), .B(\mem[11][27] ), .S(n1520), .Z(n1436)
         );
  MUX2_X1 U1558 ( .A(\mem[8][27] ), .B(\mem[9][27] ), .S(n1520), .Z(n1437) );
  MUX2_X1 U1559 ( .A(n1437), .B(n1436), .S(N11), .Z(n1438) );
  MUX2_X1 U1560 ( .A(n1438), .B(n1435), .S(n1505), .Z(n1439) );
  MUX2_X1 U1561 ( .A(\mem[6][27] ), .B(\mem[7][27] ), .S(n1521), .Z(n1440) );
  MUX2_X1 U1562 ( .A(\mem[4][27] ), .B(\mem[5][27] ), .S(n1521), .Z(n1441) );
  MUX2_X1 U1563 ( .A(n1441), .B(n1440), .S(N11), .Z(n1442) );
  MUX2_X1 U1564 ( .A(\mem[2][27] ), .B(\mem[3][27] ), .S(n1521), .Z(n1443) );
  MUX2_X1 U1565 ( .A(\mem[0][27] ), .B(\mem[1][27] ), .S(n1521), .Z(n1444) );
  MUX2_X1 U1566 ( .A(n1444), .B(n1443), .S(N11), .Z(n1445) );
  MUX2_X1 U1567 ( .A(n1445), .B(n1442), .S(n1505), .Z(n1446) );
  MUX2_X1 U1568 ( .A(\mem[14][28] ), .B(\mem[15][28] ), .S(n1521), .Z(n1447)
         );
  MUX2_X1 U1569 ( .A(\mem[12][28] ), .B(\mem[13][28] ), .S(n1521), .Z(n1448)
         );
  MUX2_X1 U1570 ( .A(n1448), .B(n1447), .S(n1506), .Z(n1449) );
  MUX2_X1 U1571 ( .A(\mem[10][28] ), .B(\mem[11][28] ), .S(n1521), .Z(n1450)
         );
  MUX2_X1 U1572 ( .A(\mem[8][28] ), .B(\mem[9][28] ), .S(n1521), .Z(n1451) );
  MUX2_X1 U1573 ( .A(n1451), .B(n1450), .S(N11), .Z(n1452) );
  MUX2_X1 U1574 ( .A(n1452), .B(n1449), .S(n1505), .Z(n1453) );
  MUX2_X1 U1575 ( .A(\mem[6][28] ), .B(\mem[7][28] ), .S(n1521), .Z(n1454) );
  MUX2_X1 U1576 ( .A(\mem[4][28] ), .B(\mem[5][28] ), .S(n1521), .Z(n1455) );
  MUX2_X1 U1577 ( .A(n1455), .B(n1454), .S(n1510), .Z(n1456) );
  MUX2_X1 U1578 ( .A(\mem[2][28] ), .B(\mem[3][28] ), .S(n1521), .Z(n1457) );
  MUX2_X1 U1579 ( .A(\mem[0][28] ), .B(\mem[1][28] ), .S(n1521), .Z(n1458) );
  MUX2_X1 U1580 ( .A(n1458), .B(n1457), .S(N11), .Z(n1459) );
  MUX2_X1 U1581 ( .A(n1459), .B(n1456), .S(n1505), .Z(n1460) );
  MUX2_X1 U1582 ( .A(n1460), .B(n1453), .S(N13), .Z(N17) );
  MUX2_X1 U1583 ( .A(\mem[14][29] ), .B(\mem[15][29] ), .S(n1522), .Z(n1461)
         );
  MUX2_X1 U1584 ( .A(\mem[12][29] ), .B(\mem[13][29] ), .S(n1522), .Z(n1462)
         );
  MUX2_X1 U1585 ( .A(n1462), .B(n1461), .S(n1506), .Z(n1463) );
  MUX2_X1 U1586 ( .A(\mem[10][29] ), .B(\mem[11][29] ), .S(n1522), .Z(n1464)
         );
  MUX2_X1 U1587 ( .A(\mem[8][29] ), .B(\mem[9][29] ), .S(n1522), .Z(n1465) );
  MUX2_X1 U1588 ( .A(n1465), .B(n1464), .S(n1509), .Z(n1466) );
  MUX2_X1 U1589 ( .A(n1466), .B(n1463), .S(n1505), .Z(n1467) );
  MUX2_X1 U1590 ( .A(\mem[6][29] ), .B(\mem[7][29] ), .S(n1522), .Z(n1468) );
  MUX2_X1 U1591 ( .A(\mem[4][29] ), .B(\mem[5][29] ), .S(n1522), .Z(n1469) );
  MUX2_X1 U1592 ( .A(n1469), .B(n1468), .S(n1507), .Z(n1470) );
  MUX2_X1 U1593 ( .A(\mem[2][29] ), .B(\mem[3][29] ), .S(n1522), .Z(n1471) );
  MUX2_X1 U1594 ( .A(\mem[0][29] ), .B(\mem[1][29] ), .S(n1522), .Z(n1472) );
  MUX2_X1 U1595 ( .A(n1472), .B(n1471), .S(N11), .Z(n1473) );
  MUX2_X1 U1596 ( .A(n1473), .B(n1470), .S(n1505), .Z(n1474) );
  MUX2_X1 U1597 ( .A(n1474), .B(n1467), .S(N13), .Z(N16) );
  MUX2_X1 U1598 ( .A(\mem[14][30] ), .B(\mem[15][30] ), .S(n1522), .Z(n1475)
         );
  MUX2_X1 U1599 ( .A(\mem[12][30] ), .B(\mem[13][30] ), .S(n1522), .Z(n1476)
         );
  MUX2_X1 U1600 ( .A(n1476), .B(n1475), .S(n1509), .Z(n1477) );
  MUX2_X1 U1601 ( .A(\mem[10][30] ), .B(\mem[11][30] ), .S(n1522), .Z(n1478)
         );
  MUX2_X1 U1602 ( .A(\mem[8][30] ), .B(\mem[9][30] ), .S(n1522), .Z(n1479) );
  MUX2_X1 U1603 ( .A(n1479), .B(n1478), .S(n1510), .Z(n1480) );
  MUX2_X1 U1604 ( .A(n1480), .B(n1477), .S(n1505), .Z(n1481) );
  MUX2_X1 U1605 ( .A(\mem[6][30] ), .B(\mem[7][30] ), .S(n1523), .Z(n1482) );
  MUX2_X1 U1606 ( .A(\mem[4][30] ), .B(\mem[5][30] ), .S(n1523), .Z(n1483) );
  MUX2_X1 U1607 ( .A(n1483), .B(n1482), .S(n1508), .Z(n1484) );
  MUX2_X1 U1608 ( .A(\mem[2][30] ), .B(\mem[3][30] ), .S(n1523), .Z(n1485) );
  MUX2_X1 U1609 ( .A(\mem[0][30] ), .B(\mem[1][30] ), .S(n1523), .Z(n1486) );
  MUX2_X1 U1610 ( .A(n1486), .B(n1485), .S(n1510), .Z(n1487) );
  MUX2_X1 U1611 ( .A(n1487), .B(n1484), .S(n1505), .Z(n1488) );
  MUX2_X1 U1612 ( .A(\mem[14][31] ), .B(\mem[15][31] ), .S(n1523), .Z(n1489)
         );
  MUX2_X1 U1613 ( .A(\mem[12][31] ), .B(\mem[13][31] ), .S(n1523), .Z(n1490)
         );
  MUX2_X1 U1614 ( .A(n1490), .B(n1489), .S(n1510), .Z(n1491) );
  MUX2_X1 U1615 ( .A(\mem[10][31] ), .B(\mem[11][31] ), .S(n1523), .Z(n1492)
         );
  MUX2_X1 U1616 ( .A(\mem[8][31] ), .B(\mem[9][31] ), .S(n1523), .Z(n1493) );
  MUX2_X1 U1617 ( .A(n1493), .B(n1492), .S(N11), .Z(n1494) );
  MUX2_X1 U1618 ( .A(n1494), .B(n1491), .S(n1505), .Z(n1495) );
  MUX2_X1 U1619 ( .A(\mem[6][31] ), .B(\mem[7][31] ), .S(n1523), .Z(n1496) );
  MUX2_X1 U1620 ( .A(\mem[4][31] ), .B(\mem[5][31] ), .S(n1523), .Z(n1497) );
  MUX2_X1 U1621 ( .A(n1497), .B(n1496), .S(n1510), .Z(n1498) );
  MUX2_X1 U1622 ( .A(\mem[2][31] ), .B(\mem[3][31] ), .S(n1523), .Z(n1499) );
  MUX2_X1 U1623 ( .A(\mem[0][31] ), .B(\mem[1][31] ), .S(n1523), .Z(n1500) );
  MUX2_X1 U1624 ( .A(n1500), .B(n1499), .S(n1510), .Z(n1501) );
  MUX2_X1 U1625 ( .A(n1501), .B(n1498), .S(n1505), .Z(n1502) );
  MUX2_X1 U1626 ( .A(n1502), .B(n1495), .S(N13), .Z(N14) );
  CLKBUF_X1 U1627 ( .A(N12), .Z(n1503) );
  CLKBUF_X1 U1628 ( .A(n543), .Z(n1530) );
  CLKBUF_X1 U1629 ( .A(n443), .Z(n1542) );
  CLKBUF_X1 U1630 ( .A(n410), .Z(n1546) );
  CLKBUF_X1 U1631 ( .A(n207), .Z(n1570) );
  CLKBUF_X1 U1632 ( .A(n106), .Z(n1582) );
  CLKBUF_X1 U1633 ( .A(n72), .Z(n1586) );
  INV_X1 U1634 ( .A(N10), .ZN(n1591) );
  INV_X1 U1635 ( .A(N11), .ZN(n1592) );
  INV_X1 U1636 ( .A(N13), .ZN(n1593) );
endmodule


module layer_13_16_1_32_W_rom ( clk, addr, z );
  input [7:0] addr;
  output [31:0] z;
  input clk;
  wire   n796, n797, n798, n799, n800, n801, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n19, n21, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n204, n207,
         n208, n209, n210, n211, n213, n214, n215, n220, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n262, n263, n264,
         n265, n266, n267, n268, n273, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n291, n292, n293, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n391, n392, n393, n394, n395, n396, n398, n399, n400,
         n405, n406, n407, n408, n409, n410, n411, n412, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n482, n483, n484, n485, n486,
         n487, n488, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n662, n663, n664, n667, n668, n669, n670, n672, n673, n674,
         n675, n676, n677, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n18, n23, n25, n26, n27, n28, n29, n30,
         n31, n32, n34, n36, n37, n38, n39, n40, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n180, n181, n182, n183,
         n202, n203, n205, n206, n212, n216, n217, n218, n219, n221, n222,
         n223, n224, n225, n226, n260, n261, n269, n270, n271, n272, n274,
         n275, n276, n277, n290, n294, n295, n296, n297, n331, n332, n333,
         n334, n360, n361, n362, n363, n387, n388, n389, n390, n397, n401,
         n402, n403, n404, n413, n435, n479, n480, n481, n489, n490, n535,
         n536, n537, n538, n595, n625, n661, n665, n666, n671, n678, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795;

  DFF_X1 \z_reg[29]  ( .D(n744), .CK(clk), .Q(z[29]), .QN(n3) );
  DFF_X1 \z_reg[28]  ( .D(n743), .CK(clk), .Q(z[28]), .QN(n4) );
  DFF_X1 \z_reg[27]  ( .D(n742), .CK(clk), .Q(z[27]), .QN(n5) );
  DFF_X1 \z_reg[26]  ( .D(n741), .CK(clk), .Q(z[26]), .QN(n6) );
  DFF_X1 \z_reg[25]  ( .D(n740), .CK(clk), .Q(z[25]), .QN(n7) );
  DFF_X1 \z_reg[24]  ( .D(n739), .CK(clk), .Q(z[24]), .QN(n8) );
  DFF_X1 \z_reg[23]  ( .D(n738), .CK(clk), .Q(z[23]), .QN(n9) );
  DFF_X1 \z_reg[22]  ( .D(n737), .CK(clk), .Q(z[22]), .QN(n10) );
  DFF_X1 \z_reg[21]  ( .D(n736), .CK(clk), .Q(z[21]), .QN(n11) );
  DFF_X1 \z_reg[20]  ( .D(n735), .CK(clk), .Q(z[20]), .QN(n12) );
  DFF_X1 \z_reg[19]  ( .D(n734), .CK(clk), .Q(z[19]), .QN(n13) );
  DFF_X1 \z_reg[18]  ( .D(n733), .CK(clk), .Q(z[18]), .QN(n14) );
  DFF_X1 \z_reg[17]  ( .D(n732), .CK(clk), .Q(z[17]), .QN(n15) );
  DFF_X1 \z_reg[16]  ( .D(n731), .CK(clk), .Q(z[16]), .QN(n16) );
  DFF_X1 \z_reg[15]  ( .D(n730), .CK(clk), .Q(z[15]), .QN(n17) );
  DFF_X1 \z_reg[14]  ( .D(n729), .CK(clk), .Q(z[14]) );
  DFF_X1 \z_reg[13]  ( .D(n728), .CK(clk), .Q(z[13]) );
  DFF_X1 \z_reg[12]  ( .D(n727), .CK(clk), .Q(z[12]) );
  DFF_X1 \z_reg[10]  ( .D(n725), .CK(clk), .Q(z[10]) );
  DFF_X1 \z_reg[5]  ( .D(n720), .CK(clk), .Q(n797), .QN(n40) );
  DFF_X1 \z_reg[0]  ( .D(n715), .CK(clk), .Q(z[0]), .QN(n36) );
  AND2_X2 U524 ( .A1(addr[7]), .A2(n795), .ZN(n714) );
  NAND3_X1 U679 ( .A1(n168), .A2(n169), .A3(n170), .ZN(n166) );
  NAND3_X1 U680 ( .A1(n171), .A2(n172), .A3(n173), .ZN(n165) );
  NAND3_X1 U681 ( .A1(n188), .A2(n189), .A3(n190), .ZN(n185) );
  NAND3_X1 U683 ( .A1(n235), .A2(n236), .A3(n237), .ZN(n177) );
  NAND3_X1 U684 ( .A1(n281), .A2(n243), .A3(n264), .ZN(n279) );
  NAND3_X1 U685 ( .A1(n302), .A2(n303), .A3(n251), .ZN(n299) );
  NAND3_X1 U686 ( .A1(n324), .A2(n194), .A3(n325), .ZN(n322) );
  NAND3_X1 U687 ( .A1(n339), .A2(n340), .A3(n267), .ZN(n336) );
  NAND3_X1 U688 ( .A1(n345), .A2(n346), .A3(n215), .ZN(n287) );
  NAND3_X1 U689 ( .A1(n358), .A2(n315), .A3(n359), .ZN(n248) );
  NAND3_X1 U690 ( .A1(n168), .A2(n172), .A3(n349), .ZN(n209) );
  NAND3_X1 U691 ( .A1(n459), .A2(n379), .A3(n460), .ZN(n293) );
  NAND3_X1 U692 ( .A1(n464), .A2(n465), .A3(n280), .ZN(n463) );
  NAND3_X1 U694 ( .A1(n472), .A2(n473), .A3(n474), .ZN(n286) );
  NAND3_X1 U696 ( .A1(n281), .A2(n189), .A3(n303), .ZN(n483) );
  NAND3_X1 U697 ( .A1(n439), .A2(n244), .A3(n436), .ZN(n510) );
  NAND3_X1 U698 ( .A1(n526), .A2(n434), .A3(n527), .ZN(n525) );
  NAND3_X1 U699 ( .A1(n301), .A2(n493), .A3(n405), .ZN(n540) );
  NAND3_X1 U700 ( .A1(n551), .A2(n512), .A3(n532), .ZN(n200) );
  NAND3_X1 U701 ( .A1(n559), .A2(n560), .A3(n561), .ZN(n446) );
  NAND3_X1 U702 ( .A1(n521), .A2(n451), .A3(n393), .ZN(n208) );
  NAND3_X1 U703 ( .A1(n313), .A2(n364), .A3(n564), .ZN(n246) );
  NAND3_X1 U704 ( .A1(n571), .A2(n572), .A3(n573), .ZN(n210) );
  NAND3_X1 U705 ( .A1(n578), .A2(n579), .A3(n580), .ZN(n327) );
  NAND3_X1 U706 ( .A1(n592), .A2(n394), .A3(n228), .ZN(n488) );
  NAND3_X1 U707 ( .A1(n593), .A2(n594), .A3(n515), .ZN(n245) );
  NAND3_X1 U708 ( .A1(n610), .A2(n576), .A3(n324), .ZN(n384) );
  NAND3_X1 U709 ( .A1(n612), .A2(n613), .A3(n614), .ZN(n198) );
  NAND3_X1 U710 ( .A1(n621), .A2(n379), .A3(n624), .ZN(n627) );
  NAND3_X1 U711 ( .A1(n191), .A2(n484), .A3(n575), .ZN(n651) );
  NAND3_X1 U712 ( .A1(n326), .A2(n440), .A3(n233), .ZN(n622) );
  NAND3_X1 U713 ( .A1(n467), .A2(n358), .A3(n654), .ZN(n604) );
  NAND3_X1 U715 ( .A1(n314), .A2(n300), .A3(n676), .ZN(n617) );
  NAND3_X1 U716 ( .A1(n444), .A2(n559), .A3(n623), .ZN(n329) );
  NAND3_X1 U717 ( .A1(n263), .A2(n249), .A3(n353), .ZN(n514) );
  NAND3_X1 U718 ( .A1(n439), .A2(n323), .A3(n473), .ZN(n616) );
  NAND3_X1 U719 ( .A1(n303), .A2(n412), .A3(n686), .ZN(n608) );
  NAND3_X1 U720 ( .A1(n451), .A2(n188), .A3(n504), .ZN(n600) );
  NAND3_X1 U721 ( .A1(n553), .A2(n511), .A3(n366), .ZN(n690) );
  NAND3_X1 U722 ( .A1(n691), .A2(n692), .A3(n693), .ZN(n220) );
  NAND3_X1 U723 ( .A1(n545), .A2(n264), .A3(n464), .ZN(n694) );
  NAND3_X1 U724 ( .A1(n588), .A2(n593), .A3(n570), .ZN(n371) );
  NAND3_X1 U725 ( .A1(n517), .A2(n557), .A3(n280), .ZN(n701) );
  NAND3_X1 U726 ( .A1(n592), .A2(n493), .A3(n534), .ZN(n317) );
  NAND3_X1 U727 ( .A1(n472), .A2(n512), .A3(n227), .ZN(n712) );
  NAND3_X1 U728 ( .A1(n494), .A2(n228), .A3(n170), .ZN(n291) );
  NAND3_X1 U729 ( .A1(n242), .A2(n229), .A3(n579), .ZN(n372) );
  DFF_X2 \z_reg[6]  ( .D(n721), .CK(clk), .Q(z[6]), .QN(n38) );
  DFF_X1 \z_reg[1]  ( .D(n716), .CK(clk), .Q(n801), .QN(n34) );
  DFF_X1 \z_reg[4]  ( .D(n719), .CK(clk), .Q(n798), .QN(n19) );
  DFF_X2 \z_reg[9]  ( .D(n724), .CK(clk), .Q(z[9]) );
  DFF_X2 \z_reg[8]  ( .D(n723), .CK(clk), .Q(z[8]), .QN(n32) );
  DFF_X2 \z_reg[11]  ( .D(n726), .CK(clk), .Q(z[11]) );
  DFF_X1 \z_reg[31]  ( .D(n746), .CK(clk), .Q(z[31]), .QN(n1) );
  DFF_X1 \z_reg[30]  ( .D(n745), .CK(clk), .Q(z[30]), .QN(n2) );
  DFF_X1 \z_reg[3]  ( .D(n718), .CK(clk), .Q(n799), .QN(n23) );
  DFF_X1 \z_reg[2]  ( .D(n717), .CK(clk), .Q(n800), .QN(n21) );
  DFF_X1 \z_reg[7]  ( .D(n722), .CK(clk), .Q(n796), .QN(n18) );
  INV_X2 U3 ( .A(n18), .ZN(z[7]) );
  NOR4_X2 U4 ( .A1(n481), .A2(n767), .A3(n582), .A4(n707), .ZN(n601) );
  AND2_X2 U5 ( .A1(n58), .A2(n57), .ZN(n45) );
  INV_X1 U6 ( .A(n34), .ZN(z[1]) );
  BUF_X4 U7 ( .A(n800), .Z(z[2]) );
  INV_X2 U8 ( .A(n23), .ZN(z[3]) );
  AND4_X1 U9 ( .A1(n301), .A2(n436), .A3(n437), .A4(n438), .ZN(n25) );
  AND3_X1 U10 ( .A1(n469), .A2(n470), .A3(n471), .ZN(n26) );
  AND3_X1 U11 ( .A1(n392), .A2(n555), .A3(n527), .ZN(n27) );
  AND4_X2 U12 ( .A1(n598), .A2(n599), .A3(n596), .A4(n597), .ZN(n28) );
  AND4_X1 U13 ( .A1(n276), .A2(n281), .A3(n681), .A4(n682), .ZN(n29) );
  AND4_X1 U14 ( .A1(n655), .A2(n656), .A3(n338), .A4(n515), .ZN(n30) );
  AND4_X1 U15 ( .A1(n522), .A2(n348), .A3(n523), .A4(n524), .ZN(n31) );
  NAND4_X2 U16 ( .A1(n626), .A2(n45), .A3(n63), .A4(n62), .ZN(n213) );
  INV_X2 U17 ( .A(n213), .ZN(n156) );
  AOI211_X4 U18 ( .C1(n799), .C2(n156), .A(n80), .B(n220), .ZN(n81) );
  INV_X2 U19 ( .A(n668), .ZN(n790) );
  INV_X2 U20 ( .A(n419), .ZN(n791) );
  NOR3_X2 U21 ( .A1(n400), .A2(n609), .A3(n94), .ZN(n62) );
  BUF_X4 U22 ( .A(n798), .Z(z[4]) );
  INV_X1 U23 ( .A(n36), .ZN(n37) );
  INV_X1 U24 ( .A(n38), .ZN(n39) );
  INV_X2 U25 ( .A(n40), .ZN(z[5]) );
  AND2_X2 U26 ( .A1(n684), .A2(n705), .ZN(n642) );
  AND2_X2 U27 ( .A1(n708), .A2(n695), .ZN(n638) );
  AND2_X1 U28 ( .A1(n697), .A2(n698), .ZN(n637) );
  AND2_X1 U29 ( .A1(n708), .A2(n709), .ZN(n485) );
  AND2_X1 U30 ( .A1(n709), .A2(n684), .ZN(n634) );
  AND2_X1 U31 ( .A1(n710), .A2(n685), .ZN(n652) );
  AND2_X1 U32 ( .A1(n695), .A2(n710), .ZN(n653) );
  AND2_X1 U33 ( .A1(n710), .A2(n705), .ZN(n640) );
  AND3_X1 U34 ( .A1(addr[6]), .A2(n698), .A3(addr[7]), .ZN(n632) );
  NOR4_X1 U35 ( .A1(n752), .A2(n198), .A3(n554), .A4(n395), .ZN(n596) );
  INV_X1 U36 ( .A(n624), .ZN(n752) );
  NOR3_X1 U37 ( .A1(n528), .A2(n179), .A3(n468), .ZN(n523) );
  NOR3_X1 U38 ( .A1(n203), .A2(n360), .A3(n202), .ZN(n374) );
  NOR2_X1 U39 ( .A1(n600), .A2(n608), .ZN(n677) );
  INV_X1 U40 ( .A(n354), .ZN(n202) );
  INV_X1 U41 ( .A(n318), .ZN(n759) );
  INV_X1 U42 ( .A(n405), .ZN(n360) );
  INV_X1 U43 ( .A(n257), .ZN(n180) );
  INV_X1 U44 ( .A(n554), .ZN(n161) );
  INV_X1 U45 ( .A(n230), .ZN(n331) );
  INV_X1 U46 ( .A(n220), .ZN(n217) );
  NAND2_X1 U47 ( .A1(n256), .A2(n257), .ZN(n234) );
  INV_X1 U48 ( .A(n312), .ZN(n763) );
  INV_X1 U49 ( .A(n358), .ZN(n780) );
  NAND4_X1 U50 ( .A1(n251), .A2(n312), .A3(n345), .A4(n169), .ZN(n707) );
  NOR4_X1 U51 ( .A1(n775), .A2(n310), .A3(n294), .A4(n781), .ZN(n599) );
  NOR4_X1 U52 ( .A1(n602), .A2(n603), .A3(n372), .A4(n604), .ZN(n597) );
  NOR4_X1 U53 ( .A1(n463), .A2(n167), .A3(n332), .A4(n766), .ZN(n462) );
  INV_X1 U54 ( .A(n170), .ZN(n766) );
  NAND4_X1 U55 ( .A1(n562), .A2(n285), .A3(n476), .A4(n563), .ZN(n259) );
  NOR4_X1 U56 ( .A1(n377), .A2(n224), .A3(n411), .A4(n222), .ZN(n563) );
  INV_X1 U57 ( .A(n281), .ZN(n224) );
  INV_X1 U58 ( .A(n366), .ZN(n222) );
  NOR4_X1 U59 ( .A1(n680), .A2(n490), .A3(n226), .A4(n402), .ZN(n679) );
  NAND4_X1 U60 ( .A1(n341), .A2(n491), .A3(n506), .A4(n594), .ZN(n680) );
  INV_X1 U61 ( .A(n455), .ZN(n490) );
  NAND2_X1 U62 ( .A1(n497), .A2(n498), .ZN(n386) );
  NOR4_X1 U63 ( .A1(n499), .A2(n239), .A3(n403), .A4(n254), .ZN(n498) );
  NOR4_X1 U64 ( .A1(n500), .A2(n501), .A3(n288), .A4(n305), .ZN(n497) );
  NAND4_X1 U65 ( .A1(n194), .A2(n433), .A3(n465), .A4(n453), .ZN(n499) );
  NOR3_X1 U66 ( .A1(n356), .A2(n382), .A3(n671), .ZN(n257) );
  NOR3_X1 U67 ( .A1(n271), .A2(n758), .A3(n566), .ZN(n621) );
  NOR2_X1 U68 ( .A1(n43), .A2(n44), .ZN(n42) );
  NAND3_X1 U69 ( .A1(n381), .A2(n470), .A3(n581), .ZN(n43) );
  OR4_X1 U70 ( .A1(n667), .A2(n261), .A3(n403), .A4(n355), .ZN(n44) );
  NOR4_X1 U71 ( .A1(n167), .A2(n388), .A3(n202), .A4(n770), .ZN(n664) );
  INV_X1 U72 ( .A(n610), .ZN(n388) );
  AOI22_X1 U73 ( .A1(n779), .A2(n790), .B1(n361), .B2(n791), .ZN(n359) );
  NOR4_X1 U74 ( .A1(n260), .A2(n356), .A3(n600), .A4(n216), .ZN(n598) );
  INV_X1 U75 ( .A(n527), .ZN(n260) );
  INV_X1 U76 ( .A(n601), .ZN(n216) );
  NAND4_X1 U77 ( .A1(n346), .A2(n455), .A3(n456), .A4(n457), .ZN(n383) );
  NOR3_X1 U78 ( .A1(n223), .A2(n458), .A3(n770), .ZN(n457) );
  NAND4_X1 U79 ( .A1(n303), .A2(n341), .A3(n263), .A4(n342), .ZN(n335) );
  NOR3_X1 U80 ( .A1(n767), .A2(n311), .A3(n187), .ZN(n342) );
  INV_X1 U81 ( .A(n636), .ZN(n361) );
  AND3_X1 U82 ( .A1(n380), .A2(n409), .A3(n394), .ZN(n136) );
  NOR3_X1 U83 ( .A1(n316), .A2(n759), .A3(n317), .ZN(n306) );
  AOI21_X1 U84 ( .B1(n786), .B2(n792), .A(n253), .ZN(n624) );
  NAND4_X1 U85 ( .A1(n601), .A2(n219), .A3(n699), .A4(n700), .ZN(n273) );
  INV_X1 U86 ( .A(n317), .ZN(n219) );
  AND3_X1 U87 ( .A1(n359), .A2(n265), .A3(n171), .ZN(n699) );
  NOR4_X1 U88 ( .A1(n701), .A2(n333), .A3(n187), .A4(n362), .ZN(n700) );
  NOR4_X1 U89 ( .A1(n239), .A2(n163), .A3(n181), .A4(n382), .ZN(n613) );
  NOR4_X1 U90 ( .A1(n615), .A2(n331), .A3(n206), .A4(n443), .ZN(n614) );
  NOR3_X1 U91 ( .A1(n396), .A2(n616), .A3(n617), .ZN(n612) );
  NOR3_X1 U92 ( .A1(n290), .A2(n458), .A3(n782), .ZN(n676) );
  INV_X1 U93 ( .A(n460), .ZN(n290) );
  NOR3_X1 U94 ( .A1(n232), .A2(n536), .A3(n231), .ZN(n654) );
  AND3_X1 U95 ( .A1(n436), .A2(n352), .A3(n465), .ZN(n686) );
  NOR3_X1 U96 ( .A1(n755), .A2(n756), .A3(n239), .ZN(n646) );
  NOR4_X1 U97 ( .A1(n648), .A2(n760), .A3(n772), .A4(n178), .ZN(n647) );
  NAND4_X1 U98 ( .A1(n369), .A2(n365), .A3(n445), .A4(n611), .ZN(n554) );
  NOR4_X1 U99 ( .A1(n162), .A2(n413), .A3(n769), .A4(n401), .ZN(n611) );
  NAND4_X1 U100 ( .A1(n555), .A2(n241), .A3(n556), .A4(n557), .ZN(n501) );
  NOR2_X1 U101 ( .A1(n558), .A2(n186), .ZN(n556) );
  NAND4_X1 U102 ( .A1(n313), .A2(n255), .A3(n434), .A4(n453), .ZN(n602) );
  NAND4_X1 U103 ( .A1(n225), .A2(n507), .A3(n508), .A4(n509), .ZN(n288) );
  NOR3_X1 U104 ( .A1(n754), .A2(n625), .A3(n167), .ZN(n508) );
  INV_X1 U105 ( .A(n514), .ZN(n225) );
  NOR4_X1 U106 ( .A1(n510), .A2(n417), .A3(n411), .A4(n785), .ZN(n509) );
  NAND4_X1 U107 ( .A1(n283), .A2(n565), .A3(n454), .A4(n426), .ZN(n528) );
  NOR4_X1 U108 ( .A1(n574), .A2(n269), .A3(n458), .A4(n751), .ZN(n573) );
  NOR3_X1 U109 ( .A1(n582), .A2(n347), .A3(n583), .ZN(n571) );
  NOR4_X1 U110 ( .A1(n232), .A2(n328), .A3(n327), .A4(n496), .ZN(n572) );
  NAND2_X1 U111 ( .A1(n790), .A2(n361), .ZN(n230) );
  NAND4_X1 U112 ( .A1(n605), .A2(n513), .A3(n606), .A4(n607), .ZN(n395) );
  NOR3_X1 U113 ( .A1(n254), .A2(n558), .A3(n770), .ZN(n606) );
  NOR4_X1 U114 ( .A1(n296), .A2(n608), .A3(n609), .A4(n384), .ZN(n607) );
  NOR4_X1 U115 ( .A1(n694), .A2(n186), .A3(n417), .A4(n311), .ZN(n693) );
  NOR3_X1 U116 ( .A1(n363), .A2(n748), .A3(n407), .ZN(n692) );
  NOR3_X1 U117 ( .A1(n273), .A2(n371), .A3(n602), .ZN(n691) );
  NAND4_X1 U118 ( .A1(n26), .A2(n205), .A3(n461), .A4(n462), .ZN(n196) );
  INV_X1 U119 ( .A(n468), .ZN(n205) );
  AND3_X1 U120 ( .A1(n368), .A2(n466), .A3(n467), .ZN(n461) );
  NAND4_X1 U121 ( .A1(n421), .A2(n169), .A3(n338), .A4(n422), .ZN(n304) );
  NOR3_X1 U122 ( .A1(n363), .A2(n665), .A3(n423), .ZN(n422) );
  NAND2_X1 U123 ( .A1(n212), .A2(n791), .ZN(n285) );
  NAND4_X1 U124 ( .A1(n264), .A2(n323), .A3(n280), .A4(n577), .ZN(n496) );
  NOR3_X1 U125 ( .A1(n199), .A2(n782), .A3(n755), .ZN(n577) );
  NAND4_X1 U126 ( .A1(n368), .A2(n428), .A3(n476), .A4(n318), .ZN(n609) );
  NAND4_X1 U127 ( .A1(n618), .A2(n249), .A3(n619), .A4(n620), .ZN(n396) );
  NOR3_X1 U128 ( .A1(n387), .A2(n535), .A3(n226), .ZN(n619) );
  AND4_X1 U129 ( .A1(n520), .A2(n578), .A3(n295), .A4(n621), .ZN(n620) );
  INV_X1 U130 ( .A(n622), .ZN(n295) );
  NAND4_X1 U131 ( .A1(n297), .A2(n495), .A3(n370), .A4(n378), .ZN(n201) );
  INV_X1 U132 ( .A(n246), .ZN(n297) );
  NAND2_X1 U133 ( .A1(n790), .A2(n765), .ZN(n312) );
  NAND4_X1 U134 ( .A1(n306), .A2(n307), .A3(n308), .A4(n309), .ZN(n289) );
  AND4_X1 U135 ( .A1(n313), .A2(n227), .A3(n314), .A4(n315), .ZN(n307) );
  NOR4_X1 U136 ( .A1(n413), .A2(n277), .A3(n402), .A4(n310), .ZN(n309) );
  NOR4_X1 U137 ( .A1(n274), .A2(n311), .A3(n763), .A4(n481), .ZN(n308) );
  NAND4_X1 U138 ( .A1(n469), .A2(n513), .A3(n230), .A4(n520), .ZN(n583) );
  AND4_X1 U139 ( .A1(n189), .A2(n250), .A3(n576), .A4(n505), .ZN(n674) );
  NOR4_X1 U140 ( .A1(n413), .A2(n769), .A3(n535), .A4(n558), .ZN(n673) );
  AOI211_X1 U141 ( .C1(n765), .C2(n791), .A(n675), .B(n617), .ZN(n672) );
  NAND4_X1 U142 ( .A1(n591), .A2(n214), .A3(n349), .A4(n589), .ZN(n399) );
  NAND4_X1 U143 ( .A1(n547), .A2(n161), .A3(n548), .A4(n549), .ZN(n344) );
  AND4_X1 U144 ( .A1(n550), .A2(n494), .A3(n492), .A4(n534), .ZN(n549) );
  NOR2_X1 U145 ( .A1(n446), .A2(n501), .ZN(n547) );
  NOR4_X1 U146 ( .A1(n760), .A2(n747), .A3(n468), .A4(n200), .ZN(n548) );
  NAND4_X1 U147 ( .A1(n373), .A2(n374), .A3(n375), .A4(n376), .ZN(n207) );
  AND3_X1 U148 ( .A1(n285), .A2(n380), .A3(n227), .ZN(n375) );
  NOR3_X1 U149 ( .A1(n780), .A2(n435), .A3(n382), .ZN(n373) );
  NOR4_X1 U150 ( .A1(n538), .A2(n277), .A3(n775), .A4(n377), .ZN(n376) );
  NAND4_X1 U151 ( .A1(n319), .A2(n182), .A3(n320), .A4(n321), .ZN(n258) );
  INV_X1 U152 ( .A(n327), .ZN(n182) );
  AOI211_X1 U153 ( .C1(n792), .C2(n786), .A(n389), .B(n390), .ZN(n320) );
  NOR4_X1 U154 ( .A1(n322), .A2(n333), .A3(n749), .A4(n186), .ZN(n321) );
  NAND2_X1 U155 ( .A1(n552), .A2(n553), .ZN(n468) );
  NAND4_X1 U156 ( .A1(n489), .A2(n440), .A3(n441), .A4(n442), .ZN(n385) );
  NOR2_X1 U157 ( .A1(n678), .A2(n536), .ZN(n441) );
  INV_X1 U158 ( .A(n446), .ZN(n489) );
  NOR4_X1 U159 ( .A1(n750), .A2(n774), .A3(n355), .A4(n443), .ZN(n442) );
  NAND2_X1 U160 ( .A1(n765), .A2(n792), .ZN(n318) );
  NAND4_X1 U161 ( .A1(n475), .A2(n215), .A3(n495), .A4(n639), .ZN(n400) );
  AND3_X1 U162 ( .A1(n424), .A2(n283), .A3(n357), .ZN(n639) );
  NAND2_X1 U163 ( .A1(n791), .A2(n779), .ZN(n192) );
  NAND4_X1 U164 ( .A1(n532), .A2(n533), .A3(n534), .A4(n312), .ZN(n174) );
  NAND2_X1 U165 ( .A1(n212), .A2(n792), .ZN(n354) );
  NAND4_X1 U166 ( .A1(n348), .A2(n349), .A3(n350), .A4(n351), .ZN(n176) );
  NOR2_X1 U167 ( .A1(n355), .A2(n203), .ZN(n350) );
  AND4_X1 U168 ( .A1(n189), .A2(n352), .A3(n353), .A4(n354), .ZN(n351) );
  INV_X1 U169 ( .A(n616), .ZN(n276) );
  NOR3_X1 U170 ( .A1(n761), .A2(n310), .A3(n776), .ZN(n681) );
  NOR2_X1 U171 ( .A1(n196), .A2(n293), .ZN(n447) );
  INV_X1 U172 ( .A(n452), .ZN(n769) );
  INV_X1 U173 ( .A(n618), .ZN(n403) );
  OR4_X1 U174 ( .A1(n316), .A2(n253), .A3(n773), .A4(n269), .ZN(n500) );
  INV_X1 U175 ( .A(n282), .ZN(n271) );
  INV_X1 U176 ( .A(n339), .ZN(n261) );
  NAND4_X1 U177 ( .A1(n451), .A2(n352), .A3(n452), .A4(n453), .ZN(n450) );
  INV_X1 U178 ( .A(n541), .ZN(n768) );
  NAND4_X1 U179 ( .A1(n241), .A2(n242), .A3(n243), .A4(n244), .ZN(n238) );
  NAND2_X1 U180 ( .A1(n791), .A2(n786), .ZN(n358) );
  INV_X1 U181 ( .A(n190), .ZN(n274) );
  INV_X1 U182 ( .A(n516), .ZN(n767) );
  NAND4_X1 U183 ( .A1(n432), .A2(n511), .A3(n188), .A4(n576), .ZN(n574) );
  INV_X1 U184 ( .A(n409), .ZN(n413) );
  NAND2_X1 U185 ( .A1(n361), .A2(n793), .ZN(n405) );
  NAND4_X1 U186 ( .A1(n282), .A2(n283), .A3(n284), .A4(n285), .ZN(n278) );
  NAND4_X1 U187 ( .A1(n191), .A2(n192), .A3(n193), .A4(n194), .ZN(n184) );
  INV_X1 U188 ( .A(n381), .ZN(n203) );
  NAND2_X1 U189 ( .A1(n786), .A2(n793), .ZN(n504) );
  INV_X1 U190 ( .A(n471), .ZN(n760) );
  INV_X1 U191 ( .A(n394), .ZN(n402) );
  INV_X1 U192 ( .A(n484), .ZN(n163) );
  OR3_X1 U193 ( .A1(n187), .A2(n186), .A3(n199), .ZN(n68) );
  NOR3_X1 U194 ( .A1(n404), .A2(n435), .A3(n389), .ZN(n655) );
  NOR4_X1 U195 ( .A1(n199), .A2(n657), .A3(n181), .A4(n180), .ZN(n656) );
  NAND2_X1 U196 ( .A1(n191), .A2(n581), .ZN(n328) );
  OR3_X1 U197 ( .A1(n178), .A2(n179), .A3(n176), .ZN(n64) );
  INV_X1 U198 ( .A(n243), .ZN(n226) );
  INV_X1 U199 ( .A(n511), .ZN(n785) );
  INV_X1 U200 ( .A(n193), .ZN(n666) );
  INV_X1 U201 ( .A(n341), .ZN(n665) );
  NOR3_X1 U202 ( .A1(n275), .A2(n768), .A3(n310), .ZN(n437) );
  NOR4_X1 U203 ( .A1(n261), .A2(n239), .A3(n231), .A4(n271), .ZN(n438) );
  INV_X1 U204 ( .A(n244), .ZN(n162) );
  INV_X1 U205 ( .A(n370), .ZN(n333) );
  INV_X1 U206 ( .A(n492), .ZN(n481) );
  INV_X1 U207 ( .A(n506), .ZN(n401) );
  INV_X1 U208 ( .A(n533), .ZN(n781) );
  INV_X1 U209 ( .A(n267), .ZN(n772) );
  INV_X1 U210 ( .A(n378), .ZN(n277) );
  OR2_X1 U211 ( .A1(n46), .A2(n47), .ZN(n247) );
  NAND4_X1 U212 ( .A1(n494), .A2(n340), .A3(n357), .A4(n495), .ZN(n46) );
  NAND4_X1 U213 ( .A1(n491), .A2(n345), .A3(n492), .A4(n493), .ZN(n47) );
  INV_X1 U214 ( .A(n542), .ZN(n535) );
  INV_X1 U215 ( .A(n605), .ZN(n755) );
  INV_X1 U216 ( .A(n562), .ZN(n536) );
  OR3_X1 U217 ( .A1(n274), .A2(n423), .A3(n407), .ZN(n179) );
  INV_X1 U218 ( .A(n459), .ZN(n782) );
  INV_X1 U219 ( .A(n623), .ZN(n387) );
  INV_X1 U220 ( .A(n590), .ZN(n223) );
  AND4_X1 U221 ( .A1(n27), .A2(n428), .A3(n429), .A4(n430), .ZN(n256) );
  AND2_X1 U222 ( .A1(n214), .A2(n283), .ZN(n429) );
  AND4_X1 U223 ( .A1(n431), .A2(n432), .A3(n433), .A4(n434), .ZN(n430) );
  OR3_X1 U224 ( .A1(n223), .A2(n254), .A3(n781), .ZN(n667) );
  NAND2_X1 U225 ( .A1(n445), .A2(n324), .ZN(n648) );
  OR3_X1 U226 ( .A1(n528), .A2(n201), .A3(n208), .ZN(n546) );
  INV_X1 U227 ( .A(n515), .ZN(n773) );
  NAND2_X1 U228 ( .A1(n337), .A2(n268), .ZN(n657) );
  AND4_X1 U229 ( .A1(n447), .A2(n218), .A3(n448), .A4(n449), .ZN(n319) );
  NOR4_X1 U230 ( .A1(n403), .A2(n178), .A3(n270), .A4(n163), .ZN(n448) );
  NOR4_X1 U231 ( .A1(n450), .A2(n202), .A3(n785), .A4(n661), .ZN(n449) );
  INV_X1 U232 ( .A(n383), .ZN(n218) );
  NOR4_X1 U233 ( .A1(n423), .A2(n683), .A3(n753), .A4(n377), .ZN(n682) );
  INV_X1 U234 ( .A(n543), .ZN(n753) );
  NAND2_X1 U235 ( .A1(n365), .A2(n364), .ZN(n683) );
  INV_X1 U236 ( .A(n575), .ZN(n269) );
  OR2_X1 U237 ( .A1(n48), .A2(n49), .ZN(n195) );
  NAND4_X1 U238 ( .A1(n266), .A2(n267), .A3(n268), .A4(n215), .ZN(n48) );
  NAND4_X1 U239 ( .A1(n262), .A2(n263), .A3(n264), .A4(n265), .ZN(n49) );
  AND3_X1 U240 ( .A1(n397), .A2(n591), .A3(n424), .ZN(n584) );
  INV_X1 U241 ( .A(n488), .ZN(n397) );
  INV_X1 U242 ( .A(n265), .ZN(n762) );
  INV_X1 U243 ( .A(n474), .ZN(n294) );
  AND4_X1 U244 ( .A1(n265), .A2(n436), .A3(n380), .A4(n505), .ZN(n550) );
  INV_X1 U245 ( .A(n324), .ZN(n747) );
  NAND2_X1 U246 ( .A1(n369), .A2(n370), .ZN(n367) );
  INV_X1 U247 ( .A(n380), .ZN(n776) );
  NAND4_X1 U248 ( .A1(n249), .A2(n250), .A3(n251), .A4(n252), .ZN(n211) );
  NOR3_X1 U249 ( .A1(n253), .A2(n778), .A3(n254), .ZN(n252) );
  INV_X1 U250 ( .A(n255), .ZN(n778) );
  INV_X1 U251 ( .A(n353), .ZN(n783) );
  INV_X1 U252 ( .A(n314), .ZN(n774) );
  INV_X1 U253 ( .A(n346), .ZN(n784) );
  INV_X1 U254 ( .A(n432), .ZN(n748) );
  INV_X1 U255 ( .A(n454), .ZN(n270) );
  INV_X1 U256 ( .A(n412), .ZN(n777) );
  INV_X1 U257 ( .A(n323), .ZN(n749) );
  INV_X1 U258 ( .A(n171), .ZN(n661) );
  INV_X1 U259 ( .A(n444), .ZN(n750) );
  INV_X1 U260 ( .A(n578), .ZN(n756) );
  INV_X1 U261 ( .A(n470), .ZN(n751) );
  INV_X1 U262 ( .A(n512), .ZN(n625) );
  AND4_X1 U263 ( .A1(n393), .A2(n474), .A3(n315), .A4(n193), .ZN(n662) );
  INV_X1 U264 ( .A(n439), .ZN(n275) );
  AND4_X1 U265 ( .A1(n194), .A2(n552), .A3(n340), .A4(n426), .ZN(n663) );
  AND3_X1 U266 ( .A1(n412), .A2(n465), .A3(n504), .ZN(n569) );
  INV_X1 U267 ( .A(n326), .ZN(n390) );
  OR2_X1 U268 ( .A1(n176), .A2(n347), .ZN(n343) );
  NOR4_X1 U269 ( .A1(n627), .A2(n771), .A3(n757), .A4(n162), .ZN(n626) );
  INV_X1 U270 ( .A(n262), .ZN(n757) );
  INV_X1 U271 ( .A(n420), .ZN(n765) );
  INV_X1 U272 ( .A(n660), .ZN(n779) );
  INV_X1 U273 ( .A(n669), .ZN(n212) );
  NOR2_X1 U274 ( .A1(n668), .A2(n669), .ZN(n254) );
  INV_X1 U275 ( .A(n635), .ZN(n792) );
  NOR2_X1 U276 ( .A1(n659), .A2(n660), .ZN(n199) );
  NOR2_X1 U277 ( .A1(n635), .A2(n660), .ZN(n458) );
  NOR2_X1 U278 ( .A1(n420), .A2(n659), .ZN(n407) );
  OAI211_X1 U279 ( .C1(n659), .C2(n669), .A(n433), .B(n266), .ZN(n582) );
  INV_X1 U280 ( .A(n659), .ZN(n793) );
  NOR2_X1 U281 ( .A1(n668), .A2(n696), .ZN(n187) );
  INV_X1 U282 ( .A(n696), .ZN(n786) );
  AND2_X1 U283 ( .A1(n643), .A2(n631), .ZN(n239) );
  NOR3_X1 U284 ( .A1(n651), .A2(n537), .A3(n240), .ZN(n650) );
  NOR3_X1 U285 ( .A1(n399), .A2(n296), .A3(n622), .ZN(n649) );
  INV_X1 U286 ( .A(n604), .ZN(n164) );
  NAND2_X1 U287 ( .A1(n633), .A2(n637), .ZN(n453) );
  NOR3_X1 U288 ( .A1(n232), .A2(n478), .A3(n773), .ZN(n477) );
  NAND4_X1 U289 ( .A1(n255), .A2(n408), .A3(n502), .A4(n503), .ZN(n305) );
  AND3_X1 U290 ( .A1(n504), .A2(n505), .A3(n506), .ZN(n502) );
  NOR4_X1 U291 ( .A1(n764), .A2(n666), .A3(n261), .A4(n296), .ZN(n503) );
  AND2_X1 U292 ( .A1(n629), .A2(n645), .ZN(n310) );
  AND2_X1 U293 ( .A1(n641), .A2(n786), .ZN(n417) );
  AND2_X1 U294 ( .A1(n640), .A2(n645), .ZN(n411) );
  NAND2_X1 U295 ( .A1(n486), .A2(n765), .ZN(n265) );
  NOR2_X1 U296 ( .A1(n635), .A2(n636), .ZN(n566) );
  NAND4_X1 U297 ( .A1(n424), .A2(n393), .A3(n359), .A4(n425), .ZN(n292) );
  AND3_X1 U298 ( .A1(n426), .A2(n427), .A3(n242), .ZN(n425) );
  NAND4_X1 U299 ( .A1(n584), .A2(n585), .A3(n586), .A4(n587), .ZN(n347) );
  AND3_X1 U300 ( .A1(n408), .A2(n453), .A3(n262), .ZN(n587) );
  AND3_X1 U301 ( .A1(n589), .A2(n590), .A3(n268), .ZN(n585) );
  NOR3_X1 U302 ( .A1(n666), .A2(n417), .A3(n332), .ZN(n586) );
  NAND2_X1 U303 ( .A1(n645), .A2(n631), .ZN(n475) );
  NAND2_X1 U304 ( .A1(n644), .A2(n485), .ZN(n474) );
  NAND2_X1 U305 ( .A1(n644), .A2(n633), .ZN(n393) );
  NAND2_X1 U306 ( .A1(n792), .A2(n642), .ZN(n194) );
  NAND4_X1 U307 ( .A1(n526), .A2(n456), .A3(n301), .A4(n713), .ZN(n603) );
  NOR3_X1 U308 ( .A1(n291), .A2(n360), .A3(n595), .ZN(n713) );
  INV_X1 U309 ( .A(n168), .ZN(n595) );
  AND2_X1 U310 ( .A1(n765), .A2(n643), .ZN(n186) );
  AND2_X1 U311 ( .A1(n637), .A2(n786), .ZN(n167) );
  NAND2_X1 U312 ( .A1(n645), .A2(n779), .ZN(n380) );
  NAND2_X1 U313 ( .A1(n765), .A2(n630), .ZN(n471) );
  NAND4_X1 U314 ( .A1(n516), .A2(n517), .A3(n518), .A4(n519), .ZN(n316) );
  NOR3_X1 U315 ( .A1(n221), .A2(n768), .A3(n418), .ZN(n518) );
  AND4_X1 U316 ( .A1(n266), .A2(n520), .A3(n230), .A4(n475), .ZN(n519) );
  INV_X1 U317 ( .A(n521), .ZN(n221) );
  AND2_X1 U318 ( .A1(n645), .A2(n786), .ZN(n232) );
  OAI21_X1 U319 ( .B1(n419), .B2(n420), .A(n337), .ZN(n416) );
  NAND2_X1 U320 ( .A1(n645), .A2(n652), .ZN(n394) );
  NAND2_X1 U321 ( .A1(n629), .A2(n628), .ZN(n340) );
  NAND2_X1 U322 ( .A1(n644), .A2(n640), .ZN(n215) );
  NAND2_X1 U323 ( .A1(n641), .A2(n212), .ZN(n436) );
  NAND2_X1 U324 ( .A1(n485), .A2(n645), .ZN(n378) );
  NAND2_X1 U325 ( .A1(n645), .A2(n638), .ZN(n243) );
  NAND2_X1 U326 ( .A1(n486), .A2(n633), .ZN(n495) );
  NAND2_X1 U327 ( .A1(n486), .A2(n642), .ZN(n193) );
  NAND2_X1 U328 ( .A1(n628), .A2(n642), .ZN(n324) );
  NAND2_X1 U329 ( .A1(n644), .A2(n629), .ZN(n513) );
  NAND4_X1 U330 ( .A1(n256), .A2(n334), .A3(n414), .A4(n415), .ZN(n197) );
  NOR4_X1 U331 ( .A1(n416), .A2(n417), .A3(n418), .A4(n783), .ZN(n415) );
  INV_X1 U332 ( .A(n292), .ZN(n334) );
  NOR2_X1 U333 ( .A1(n209), .A2(n304), .ZN(n414) );
  NAND4_X1 U334 ( .A1(n217), .A2(n687), .A3(n688), .A4(n689), .ZN(n398) );
  NAND2_X1 U335 ( .A1(n485), .A2(n486), .ZN(n687) );
  AND3_X1 U336 ( .A1(n408), .A2(n172), .A3(n521), .ZN(n688) );
  NOR4_X1 U337 ( .A1(n690), .A2(n411), .A3(n274), .A4(n784), .ZN(n689) );
  NAND2_X1 U338 ( .A1(n486), .A2(n638), .ZN(n281) );
  NAND2_X1 U339 ( .A1(n634), .A2(n793), .ZN(n492) );
  NAND2_X1 U340 ( .A1(n791), .A2(n652), .ZN(n241) );
  NAND2_X1 U341 ( .A1(n658), .A2(n791), .ZN(n301) );
  NAND2_X1 U342 ( .A1(n637), .A2(n642), .ZN(n520) );
  NAND2_X1 U343 ( .A1(n486), .A2(n640), .ZN(n433) );
  NAND2_X1 U344 ( .A1(n790), .A2(n658), .ZN(n264) );
  NAND2_X1 U345 ( .A1(n641), .A2(n361), .ZN(n370) );
  NAND2_X1 U346 ( .A1(n630), .A2(n779), .ZN(n255) );
  NAND2_X1 U347 ( .A1(n637), .A2(n631), .ZN(n189) );
  NAND2_X1 U348 ( .A1(n790), .A2(n642), .ZN(n283) );
  NAND2_X1 U349 ( .A1(n212), .A2(n637), .ZN(n484) );
  NAND2_X1 U350 ( .A1(n709), .A2(n710), .ZN(n636) );
  AND2_X1 U351 ( .A1(n765), .A2(n641), .ZN(n377) );
  AND2_X1 U352 ( .A1(n644), .A2(n212), .ZN(n231) );
  NAND2_X1 U353 ( .A1(n644), .A2(n765), .ZN(n476) );
  NAND2_X1 U354 ( .A1(n629), .A2(n793), .ZN(n428) );
  NAND2_X1 U355 ( .A1(n644), .A2(n642), .ZN(n341) );
  NAND2_X1 U356 ( .A1(n628), .A2(n631), .ZN(n576) );
  NAND2_X1 U357 ( .A1(n633), .A2(n793), .ZN(n432) );
  NAND2_X1 U358 ( .A1(n629), .A2(n637), .ZN(n594) );
  NAND2_X1 U359 ( .A1(n638), .A2(n637), .ZN(n369) );
  NAND2_X1 U360 ( .A1(n634), .A2(n628), .ZN(n426) );
  NAND2_X1 U361 ( .A1(n658), .A2(n628), .ZN(n505) );
  AND2_X1 U362 ( .A1(n793), .A2(n652), .ZN(n443) );
  NAND2_X1 U363 ( .A1(n486), .A2(n653), .ZN(n280) );
  AND2_X1 U364 ( .A1(n792), .A2(n652), .ZN(n355) );
  AND2_X1 U365 ( .A1(n790), .A2(n653), .ZN(n382) );
  AND2_X1 U366 ( .A1(n644), .A2(n779), .ZN(n558) );
  AND2_X1 U367 ( .A1(n653), .A2(n643), .ZN(n311) );
  NAND2_X1 U368 ( .A1(n628), .A2(n212), .ZN(n244) );
  NAND2_X1 U369 ( .A1(n645), .A2(n361), .ZN(n266) );
  NAND4_X1 U370 ( .A1(n532), .A2(n369), .A3(n192), .A4(n670), .ZN(n330) );
  NOR2_X1 U371 ( .A1(n443), .A2(n478), .ZN(n670) );
  NAND4_X1 U372 ( .A1(n183), .A2(n475), .A3(n567), .A4(n568), .ZN(n175) );
  AND3_X1 U373 ( .A1(n300), .A2(n456), .A3(n460), .ZN(n567) );
  AND3_X1 U374 ( .A1(n569), .A2(n517), .A3(n570), .ZN(n568) );
  INV_X1 U375 ( .A(n210), .ZN(n183) );
  NAND2_X1 U376 ( .A1(n486), .A2(n779), .ZN(n314) );
  AND2_X1 U377 ( .A1(n640), .A2(n630), .ZN(n423) );
  NAND2_X1 U378 ( .A1(n640), .A2(n637), .ZN(n434) );
  NAND2_X1 U379 ( .A1(n638), .A2(n628), .ZN(n227) );
  NAND2_X1 U380 ( .A1(n485), .A2(n792), .ZN(n465) );
  NAND2_X1 U381 ( .A1(n486), .A2(n786), .ZN(n511) );
  NAND2_X1 U382 ( .A1(n658), .A2(n645), .ZN(n534) );
  NAND2_X1 U383 ( .A1(n637), .A2(n779), .ZN(n267) );
  NAND2_X1 U384 ( .A1(n634), .A2(n791), .ZN(n315) );
  NAND2_X1 U385 ( .A1(n641), .A2(n652), .ZN(n263) );
  NOR3_X1 U386 ( .A1(n245), .A2(n271), .A3(n246), .ZN(n236) );
  NOR4_X1 U387 ( .A1(n238), .A2(n759), .A3(n239), .A4(n240), .ZN(n237) );
  NOR3_X1 U388 ( .A1(n247), .A2(n248), .A3(n211), .ZN(n235) );
  NAND2_X1 U389 ( .A1(n765), .A2(n628), .ZN(n464) );
  NAND2_X1 U390 ( .A1(n361), .A2(n630), .ZN(n169) );
  NAND2_X1 U391 ( .A1(n485), .A2(n793), .ZN(n467) );
  NAND2_X1 U392 ( .A1(n791), .A2(n631), .ZN(n532) );
  NAND2_X1 U393 ( .A1(n641), .A2(n642), .ZN(n445) );
  NAND2_X1 U394 ( .A1(n630), .A2(n652), .ZN(n506) );
  NAND2_X1 U395 ( .A1(n644), .A2(n652), .ZN(n268) );
  NAND2_X1 U396 ( .A1(n765), .A2(n637), .ZN(n507) );
  INV_X1 U397 ( .A(n427), .ZN(n775) );
  NAND2_X1 U398 ( .A1(n765), .A2(n645), .ZN(n431) );
  NAND2_X1 U399 ( .A1(n658), .A2(n792), .ZN(n456) );
  NAND2_X1 U400 ( .A1(n643), .A2(n652), .ZN(n349) );
  NAND2_X1 U401 ( .A1(n638), .A2(n630), .ZN(n345) );
  NAND2_X1 U402 ( .A1(n638), .A2(n793), .ZN(n454) );
  NAND2_X1 U403 ( .A1(n485), .A2(n637), .ZN(n352) );
  NAND2_X1 U404 ( .A1(n643), .A2(n786), .ZN(n353) );
  NAND2_X1 U405 ( .A1(n633), .A2(n645), .ZN(n444) );
  NAND2_X1 U406 ( .A1(n633), .A2(n791), .ZN(n466) );
  NAND2_X1 U407 ( .A1(n658), .A2(n643), .ZN(n303) );
  NAND2_X1 U408 ( .A1(n628), .A2(n652), .ZN(n529) );
  NAND2_X1 U409 ( .A1(n628), .A2(n361), .ZN(n242) );
  NAND2_X1 U410 ( .A1(n633), .A2(n792), .ZN(n323) );
  NAND2_X1 U411 ( .A1(n629), .A2(n643), .ZN(n578) );
  NAND2_X1 U412 ( .A1(n644), .A2(n786), .ZN(n346) );
  NAND2_X1 U413 ( .A1(n790), .A2(n638), .ZN(n339) );
  NAND2_X1 U414 ( .A1(n485), .A2(n790), .ZN(n251) );
  NAND2_X1 U415 ( .A1(n790), .A2(n631), .ZN(n365) );
  INV_X1 U416 ( .A(n564), .ZN(n296) );
  NAND2_X1 U417 ( .A1(n629), .A2(n630), .ZN(n262) );
  NAND2_X1 U418 ( .A1(n658), .A2(n793), .ZN(n337) );
  NAND2_X1 U419 ( .A1(n628), .A2(n779), .ZN(n515) );
  NAND2_X1 U420 ( .A1(n638), .A2(n641), .ZN(n249) );
  NAND2_X1 U421 ( .A1(n486), .A2(n634), .ZN(n421) );
  NAND2_X1 U422 ( .A1(n486), .A2(n658), .ZN(n366) );
  AND2_X1 U423 ( .A1(n212), .A2(n630), .ZN(n178) );
  NAND2_X1 U424 ( .A1(n653), .A2(n645), .ZN(n494) );
  NAND4_X1 U425 ( .A1(n570), .A2(n545), .A3(n444), .A4(n594), .ZN(n615) );
  NAND2_X1 U426 ( .A1(n628), .A2(n786), .ZN(n533) );
  NAND2_X1 U427 ( .A1(n641), .A2(n779), .ZN(n412) );
  NAND2_X1 U428 ( .A1(n633), .A2(n641), .ZN(n313) );
  NAND2_X1 U429 ( .A1(n629), .A2(n792), .ZN(n191) );
  AND2_X1 U430 ( .A1(n643), .A2(n212), .ZN(n356) );
  NAND2_X1 U431 ( .A1(n643), .A2(n642), .ZN(n493) );
  NAND2_X1 U432 ( .A1(n486), .A2(n629), .ZN(n605) );
  NAND2_X1 U433 ( .A1(n486), .A2(n631), .ZN(n541) );
  NAND2_X1 U434 ( .A1(n630), .A2(n631), .ZN(n250) );
  NAND2_X1 U435 ( .A1(n637), .A2(n652), .ZN(n618) );
  NAND2_X1 U436 ( .A1(n641), .A2(n631), .ZN(n452) );
  NAND2_X1 U437 ( .A1(n643), .A2(n361), .ZN(n338) );
  NAND2_X1 U438 ( .A1(n644), .A2(n638), .ZN(n517) );
  NAND2_X1 U439 ( .A1(n644), .A2(n653), .ZN(n214) );
  OR4_X1 U440 ( .A1(n479), .A2(n199), .A3(n240), .A4(n203), .ZN(n298) );
  NAND2_X1 U441 ( .A1(n653), .A2(n628), .ZN(n302) );
  AND2_X1 U442 ( .A1(n633), .A2(n630), .ZN(n253) );
  NAND2_X1 U443 ( .A1(n640), .A2(n641), .ZN(n357) );
  NAND2_X1 U444 ( .A1(n486), .A2(n652), .ZN(n233) );
  NAND2_X1 U445 ( .A1(n653), .A2(n637), .ZN(n188) );
  NAND2_X1 U446 ( .A1(n791), .A2(n642), .ZN(n561) );
  NAND2_X1 U447 ( .A1(n644), .A2(n631), .ZN(n516) );
  NAND2_X1 U448 ( .A1(n790), .A2(n633), .ZN(n364) );
  NAND2_X1 U449 ( .A1(n485), .A2(n641), .ZN(n460) );
  NAND2_X1 U450 ( .A1(n486), .A2(n212), .ZN(n553) );
  NAND2_X1 U451 ( .A1(n642), .A2(n793), .ZN(n171) );
  NAND2_X1 U452 ( .A1(n653), .A2(n630), .ZN(n565) );
  NAND2_X1 U453 ( .A1(n642), .A2(n630), .ZN(n512) );
  NAND2_X1 U454 ( .A1(n638), .A2(n791), .ZN(n527) );
  NAND2_X1 U455 ( .A1(n793), .A2(n631), .ZN(n170) );
  NAND2_X1 U456 ( .A1(n485), .A2(n630), .ZN(n439) );
  NAND2_X1 U457 ( .A1(n633), .A2(n643), .ZN(n470) );
  NAND2_X1 U458 ( .A1(n790), .A2(n640), .ZN(n545) );
  NAND2_X1 U459 ( .A1(n645), .A2(n642), .ZN(n472) );
  NAND2_X1 U460 ( .A1(n629), .A2(n641), .ZN(n543) );
  NAND2_X1 U461 ( .A1(n634), .A2(n637), .ZN(n451) );
  NAND2_X1 U462 ( .A1(n640), .A2(n643), .ZN(n424) );
  NAND2_X1 U463 ( .A1(n640), .A2(n793), .ZN(n368) );
  NAND2_X1 U464 ( .A1(n643), .A2(n779), .ZN(n557) );
  NAND2_X1 U465 ( .A1(n634), .A2(n645), .ZN(n455) );
  NAND2_X1 U466 ( .A1(n634), .A2(n643), .ZN(n542) );
  NAND2_X1 U467 ( .A1(n792), .A2(n631), .ZN(n284) );
  NAND2_X1 U468 ( .A1(n658), .A2(n641), .ZN(n491) );
  NAND2_X1 U469 ( .A1(n790), .A2(n629), .ZN(n552) );
  NAND2_X1 U470 ( .A1(n644), .A2(n361), .ZN(n581) );
  NAND2_X1 U471 ( .A1(n645), .A2(n212), .ZN(n381) );
  NAND2_X1 U472 ( .A1(n634), .A2(n630), .ZN(n562) );
  NAND2_X1 U473 ( .A1(n644), .A2(n658), .ZN(n392) );
  NAND2_X1 U474 ( .A1(n638), .A2(n792), .ZN(n282) );
  NAND2_X1 U475 ( .A1(n643), .A2(n638), .ZN(n575) );
  NAND2_X1 U476 ( .A1(n637), .A2(n361), .ZN(n588) );
  NAND2_X1 U477 ( .A1(n486), .A2(n361), .ZN(n579) );
  NAND2_X1 U478 ( .A1(n634), .A2(n792), .ZN(n589) );
  NAND2_X1 U479 ( .A1(n790), .A2(n652), .ZN(n228) );
  NAND2_X1 U480 ( .A1(n485), .A2(n628), .ZN(n440) );
  NAND2_X1 U481 ( .A1(n485), .A2(n791), .ZN(n469) );
  NAND2_X1 U482 ( .A1(n485), .A2(n643), .ZN(n190) );
  NAND2_X1 U483 ( .A1(n629), .A2(n791), .ZN(n300) );
  NAND2_X1 U484 ( .A1(n640), .A2(n628), .ZN(n409) );
  NAND2_X1 U485 ( .A1(n658), .A2(n630), .ZN(n590) );
  NAND2_X1 U486 ( .A1(n644), .A2(n634), .ZN(n592) );
  NAND2_X1 U487 ( .A1(n633), .A2(n628), .ZN(n555) );
  NAND2_X1 U488 ( .A1(n653), .A2(n641), .ZN(n326) );
  NAND2_X1 U489 ( .A1(n786), .A2(n630), .ZN(n459) );
  NAND2_X1 U490 ( .A1(n653), .A2(n793), .ZN(n623) );
  NAND2_X1 U491 ( .A1(n653), .A2(n792), .ZN(n610) );
  NAND2_X1 U492 ( .A1(n653), .A2(n791), .ZN(n526) );
  NAND2_X1 U493 ( .A1(n640), .A2(n791), .ZN(n591) );
  NOR3_X1 U494 ( .A1(n401), .A2(n771), .A3(n775), .ZN(n173) );
  NOR2_X1 U495 ( .A1(n772), .A2(n240), .ZN(n522) );
  NOR4_X1 U496 ( .A1(n525), .A2(n762), .A3(n769), .A4(n665), .ZN(n524) );
  INV_X1 U497 ( .A(n580), .ZN(n181) );
  OR4_X1 U498 ( .A1(n768), .A2(n418), .A3(n514), .A4(n329), .ZN(n50) );
  INV_X1 U499 ( .A(n560), .ZN(n771) );
  NAND2_X1 U500 ( .A1(n790), .A2(n634), .ZN(n229) );
  NAND2_X1 U501 ( .A1(n634), .A2(n641), .ZN(n559) );
  NAND2_X1 U502 ( .A1(n658), .A2(n637), .ZN(n593) );
  INV_X1 U503 ( .A(n531), .ZN(n363) );
  NAND2_X1 U504 ( .A1(n640), .A2(n792), .ZN(n325) );
  NAND4_X1 U505 ( .A1(n541), .A2(n542), .A3(n543), .A4(n544), .ZN(n539) );
  AND3_X1 U506 ( .A1(n302), .A2(n473), .A3(n545), .ZN(n544) );
  AND4_X1 U507 ( .A1(n466), .A2(n474), .A3(n529), .A4(n530), .ZN(n348) );
  AND3_X1 U508 ( .A1(n472), .A2(n464), .A3(n531), .ZN(n530) );
  NOR3_X1 U509 ( .A1(n767), .A2(n272), .A3(n407), .ZN(n406) );
  NOR3_X1 U510 ( .A1(n411), .A2(n777), .A3(n387), .ZN(n410) );
  INV_X1 U511 ( .A(n408), .ZN(n272) );
  NAND2_X1 U512 ( .A1(n427), .A2(n378), .ZN(n675) );
  INV_X1 U513 ( .A(n379), .ZN(n538) );
  NOR2_X1 U514 ( .A1(n480), .A2(n787), .ZN(n710) );
  NOR2_X1 U515 ( .A1(n789), .A2(n788), .ZN(n709) );
  AND2_X2 U516 ( .A1(n703), .A2(n698), .ZN(n628) );
  AND2_X2 U517 ( .A1(n706), .A2(n714), .ZN(n486) );
  AND2_X1 U518 ( .A1(n703), .A2(n704), .ZN(n641) );
  AND2_X1 U519 ( .A1(n697), .A2(n711), .ZN(n630) );
  AND2_X2 U520 ( .A1(n714), .A2(n698), .ZN(n645) );
  AND2_X1 U521 ( .A1(n703), .A2(n711), .ZN(n644) );
  AND2_X1 U522 ( .A1(n706), .A2(n703), .ZN(n643) );
  AND2_X1 U523 ( .A1(n685), .A2(n702), .ZN(n631) );
  AND2_X1 U525 ( .A1(n708), .A2(n705), .ZN(n658) );
  AND2_X1 U526 ( .A1(n695), .A2(n684), .ZN(n633) );
  AND2_X1 U527 ( .A1(n684), .A2(n685), .ZN(n629) );
  NAND2_X1 U528 ( .A1(n714), .A2(n711), .ZN(n659) );
  NAND2_X1 U529 ( .A1(n706), .A2(n697), .ZN(n668) );
  NAND2_X1 U530 ( .A1(n704), .A2(n697), .ZN(n635) );
  AND2_X1 U531 ( .A1(n640), .A2(n632), .ZN(n240) );
  NAND2_X1 U532 ( .A1(n705), .A2(n702), .ZN(n660) );
  NAND2_X1 U533 ( .A1(n779), .A2(n632), .ZN(n427) );
  NAND2_X1 U534 ( .A1(n708), .A2(n685), .ZN(n669) );
  NAND2_X1 U535 ( .A1(n485), .A2(n632), .ZN(n408) );
  NAND2_X1 U536 ( .A1(n709), .A2(n702), .ZN(n420) );
  NAND2_X1 U537 ( .A1(n695), .A2(n702), .ZN(n696) );
  AND2_X1 U538 ( .A1(n638), .A2(n632), .ZN(n418) );
  NAND2_X1 U539 ( .A1(n704), .A2(n714), .ZN(n419) );
  NAND4_X1 U540 ( .A1(n392), .A2(n339), .A3(n393), .A4(n394), .ZN(n391) );
  NAND4_X1 U541 ( .A1(n428), .A2(n467), .A3(n484), .A4(n471), .ZN(n482) );
  OR2_X1 U542 ( .A1(n488), .A2(n247), .ZN(n487) );
  OR4_X1 U543 ( .A1(n208), .A2(n209), .A3(n210), .A4(n211), .ZN(n204) );
  NAND2_X1 U544 ( .A1(n212), .A2(n632), .ZN(n580) );
  NAND2_X1 U545 ( .A1(n765), .A2(n632), .ZN(n551) );
  NAND2_X1 U546 ( .A1(n658), .A2(n632), .ZN(n521) );
  AND2_X1 U547 ( .A1(n629), .A2(n632), .ZN(n478) );
  NAND2_X1 U548 ( .A1(n634), .A2(n632), .ZN(n379) );
  NAND2_X1 U549 ( .A1(n642), .A2(n632), .ZN(n168) );
  NAND2_X1 U550 ( .A1(n786), .A2(n632), .ZN(n570) );
  NAND2_X1 U551 ( .A1(n652), .A2(n632), .ZN(n172) );
  NAND2_X1 U552 ( .A1(n633), .A2(n632), .ZN(n473) );
  NAND2_X1 U553 ( .A1(n631), .A2(n632), .ZN(n560) );
  NAND2_X1 U554 ( .A1(n653), .A2(n632), .ZN(n531) );
  NAND2_X1 U555 ( .A1(n361), .A2(n632), .ZN(n564) );
  NOR2_X1 U556 ( .A1(addr[5]), .A2(addr[4]), .ZN(n698) );
  NOR2_X1 U557 ( .A1(n787), .A2(addr[0]), .ZN(n702) );
  NOR2_X1 U558 ( .A1(n788), .A2(addr[3]), .ZN(n685) );
  NOR2_X1 U559 ( .A1(n789), .A2(addr[2]), .ZN(n705) );
  NOR2_X1 U560 ( .A1(addr[1]), .A2(addr[0]), .ZN(n684) );
  NOR2_X1 U561 ( .A1(addr[7]), .A2(addr[6]), .ZN(n697) );
  NOR2_X1 U562 ( .A1(n795), .A2(addr[7]), .ZN(n703) );
  NOR2_X1 U563 ( .A1(addr[3]), .A2(addr[2]), .ZN(n695) );
  NOR2_X1 U564 ( .A1(n480), .A2(addr[1]), .ZN(n708) );
  NOR2_X1 U565 ( .A1(n794), .A2(addr[4]), .ZN(n706) );
  OAI21_X1 U566 ( .B1(n51), .B2(n2), .A(n28), .ZN(n745) );
  OAI21_X1 U567 ( .B1(n52), .B2(n3), .A(n28), .ZN(n744) );
  OAI21_X1 U568 ( .B1(n213), .B2(n1), .A(n28), .ZN(n746) );
  AND2_X1 U569 ( .A1(addr[5]), .A2(addr[4]), .ZN(n711) );
  AND2_X1 U570 ( .A1(addr[4]), .A2(n794), .ZN(n704) );
  INV_X1 U571 ( .A(addr[0]), .ZN(n480) );
  INV_X1 U572 ( .A(addr[2]), .ZN(n788) );
  INV_X1 U573 ( .A(addr[1]), .ZN(n787) );
  INV_X1 U574 ( .A(addr[3]), .ZN(n789) );
  INV_X1 U575 ( .A(addr[6]), .ZN(n795) );
  INV_X1 U576 ( .A(addr[5]), .ZN(n794) );
  NAND4_X1 U577 ( .A1(n626), .A2(n45), .A3(n63), .A4(n62), .ZN(n51) );
  NAND4_X1 U578 ( .A1(n626), .A2(n45), .A3(n63), .A4(n62), .ZN(n52) );
  NAND4_X1 U579 ( .A1(n673), .A2(n674), .A3(n679), .A4(n672), .ZN(n54) );
  INV_X1 U580 ( .A(n285), .ZN(n206) );
  INV_X1 U581 ( .A(n677), .ZN(n53) );
  NOR4_X1 U582 ( .A1(n54), .A2(n206), .A3(n50), .A4(n53), .ZN(n58) );
  INV_X1 U583 ( .A(n603), .ZN(n79) );
  INV_X1 U584 ( .A(n398), .ZN(n55) );
  NAND3_X1 U585 ( .A1(n79), .A2(n55), .A3(n29), .ZN(n56) );
  INV_X1 U586 ( .A(n551), .ZN(n764) );
  NOR4_X1 U587 ( .A1(n56), .A2(n712), .A3(n372), .A4(n764), .ZN(n57) );
  NAND3_X1 U588 ( .A1(n241), .A2(n466), .A3(n27), .ZN(n60) );
  NAND4_X1 U589 ( .A1(n663), .A2(n664), .A3(n662), .A4(n42), .ZN(n59) );
  OR4_X1 U590 ( .A1(n330), .A2(n583), .A3(n60), .A4(n59), .ZN(n78) );
  INV_X1 U591 ( .A(n78), .ZN(n63) );
  NAND4_X1 U592 ( .A1(n649), .A2(n650), .A3(n164), .A4(n30), .ZN(n100) );
  INV_X1 U593 ( .A(n100), .ZN(n61) );
  NAND4_X1 U594 ( .A1(n646), .A2(n647), .A3(n454), .A4(n61), .ZN(n94) );
  INV_X1 U595 ( .A(n192), .ZN(n73) );
  INV_X1 U596 ( .A(n445), .ZN(n678) );
  INV_X1 U597 ( .A(n284), .ZN(n770) );
  NOR4_X1 U598 ( .A1(n175), .A2(n73), .A3(n678), .A4(n770), .ZN(n67) );
  AOI211_X1 U599 ( .C1(n37), .C2(n156), .A(n177), .B(n174), .ZN(n66) );
  NOR4_X1 U600 ( .A1(n64), .A2(n167), .A3(n166), .A4(n165), .ZN(n65) );
  NAND3_X1 U601 ( .A1(n67), .A2(n66), .A3(n65), .ZN(n715) );
  INV_X1 U602 ( .A(n529), .ZN(n404) );
  NOR4_X1 U603 ( .A1(n195), .A2(n198), .A3(n197), .A4(n404), .ZN(n71) );
  AOI211_X1 U604 ( .C1(n801), .C2(n156), .A(n185), .B(n200), .ZN(n70) );
  NOR4_X1 U605 ( .A1(n68), .A2(n184), .A3(n196), .A4(n201), .ZN(n69) );
  NAND3_X1 U606 ( .A1(n71), .A2(n70), .A3(n69), .ZN(n716) );
  NOR2_X1 U607 ( .A1(n21), .A2(n51), .ZN(n77) );
  INV_X1 U608 ( .A(n207), .ZN(n72) );
  NAND3_X1 U609 ( .A1(n31), .A2(n25), .A3(n72), .ZN(n76) );
  INV_X1 U610 ( .A(n431), .ZN(n761) );
  INV_X1 U611 ( .A(n338), .ZN(n113) );
  NOR3_X1 U612 ( .A1(n761), .A2(n113), .A3(n73), .ZN(n74) );
  NAND4_X1 U613 ( .A1(n215), .A2(n421), .A3(n214), .A4(n74), .ZN(n75) );
  OR4_X1 U614 ( .A1(n204), .A2(n77), .A3(n76), .A4(n75), .ZN(n717) );
  INV_X1 U615 ( .A(n712), .ZN(n83) );
  NOR3_X1 U616 ( .A1(n78), .A2(n764), .A3(n206), .ZN(n82) );
  NAND2_X1 U617 ( .A1(n79), .A2(n29), .ZN(n80) );
  NAND4_X1 U618 ( .A1(n30), .A2(n83), .A3(n82), .A4(n81), .ZN(n718) );
  OAI21_X1 U619 ( .B1(n19), .B2(n51), .A(n45), .ZN(n719) );
  NAND4_X1 U620 ( .A1(n230), .A2(n233), .A3(n227), .A4(n513), .ZN(n86) );
  INV_X1 U621 ( .A(n228), .ZN(n85) );
  INV_X1 U622 ( .A(n229), .ZN(n84) );
  NOR4_X1 U623 ( .A1(n86), .A2(n259), .A3(n85), .A4(n84), .ZN(n92) );
  INV_X1 U624 ( .A(n231), .ZN(n89) );
  INV_X1 U625 ( .A(n258), .ZN(n88) );
  AOI21_X1 U626 ( .B1(n797), .B2(n156), .A(n177), .ZN(n87) );
  NAND3_X1 U627 ( .A1(n89), .A2(n88), .A3(n87), .ZN(n90) );
  NOR4_X1 U628 ( .A1(n90), .A2(n234), .A3(n232), .A4(n195), .ZN(n91) );
  NAND2_X1 U629 ( .A1(n92), .A2(n91), .ZN(n720) );
  INV_X1 U630 ( .A(n679), .ZN(n93) );
  INV_X1 U631 ( .A(n241), .ZN(n141) );
  NOR3_X1 U632 ( .A1(n50), .A2(n93), .A3(n141), .ZN(n98) );
  INV_X1 U633 ( .A(n94), .ZN(n95) );
  NAND3_X1 U634 ( .A1(n95), .A2(n677), .A3(n29), .ZN(n96) );
  AOI211_X1 U635 ( .C1(n39), .C2(n156), .A(n96), .B(n273), .ZN(n97) );
  NAND4_X1 U636 ( .A1(n466), .A2(n42), .A3(n98), .A4(n97), .ZN(n721) );
  INV_X1 U637 ( .A(n588), .ZN(n332) );
  INV_X1 U638 ( .A(n280), .ZN(n99) );
  NOR4_X1 U639 ( .A1(n286), .A2(n100), .A3(n332), .A4(n99), .ZN(n104) );
  AOI211_X1 U640 ( .C1(n796), .C2(n156), .A(n289), .B(n287), .ZN(n103) );
  NOR3_X1 U641 ( .A1(n279), .A2(n293), .A3(n291), .ZN(n102) );
  NOR3_X1 U642 ( .A1(n278), .A2(n292), .A3(n288), .ZN(n101) );
  NAND4_X1 U643 ( .A1(n104), .A2(n103), .A3(n102), .A4(n101), .ZN(n722) );
  NOR3_X1 U644 ( .A1(n304), .A2(n305), .A3(n299), .ZN(n111) );
  NOR3_X1 U645 ( .A1(n298), .A2(n289), .A3(n258), .ZN(n110) );
  INV_X1 U646 ( .A(n328), .ZN(n123) );
  INV_X1 U647 ( .A(n329), .ZN(n105) );
  OAI211_X1 U648 ( .C1(n52), .C2(n32), .A(n123), .B(n105), .ZN(n108) );
  INV_X1 U649 ( .A(n300), .ZN(n107) );
  INV_X1 U650 ( .A(n301), .ZN(n106) );
  NOR4_X1 U651 ( .A1(n108), .A2(n330), .A3(n107), .A4(n106), .ZN(n109) );
  NAND3_X1 U652 ( .A1(n111), .A2(n110), .A3(n109), .ZN(n723) );
  INV_X1 U653 ( .A(n357), .ZN(n479) );
  INV_X1 U654 ( .A(n337), .ZN(n112) );
  NOR4_X1 U655 ( .A1(n344), .A2(n113), .A3(n479), .A4(n112), .ZN(n117) );
  AOI211_X1 U656 ( .C1(z[9]), .C2(n156), .A(n248), .B(n198), .ZN(n116) );
  NOR3_X1 U657 ( .A1(n356), .A2(n336), .A3(n287), .ZN(n115) );
  NOR3_X1 U658 ( .A1(n335), .A2(n343), .A3(n231), .ZN(n114) );
  NAND4_X1 U659 ( .A1(n117), .A2(n116), .A3(n115), .A4(n114), .ZN(n724) );
  INV_X1 U660 ( .A(n364), .ZN(n120) );
  INV_X1 U661 ( .A(n365), .ZN(n119) );
  INV_X1 U662 ( .A(n368), .ZN(n118) );
  NOR4_X1 U663 ( .A1(n120), .A2(n119), .A3(n118), .A4(n226), .ZN(n127) );
  NOR4_X1 U664 ( .A1(n385), .A2(n386), .A3(n372), .A4(n222), .ZN(n126) );
  INV_X1 U665 ( .A(n384), .ZN(n122) );
  AOI21_X1 U666 ( .B1(z[10]), .B2(n156), .A(n371), .ZN(n121) );
  NAND3_X1 U667 ( .A1(n123), .A2(n122), .A3(n121), .ZN(n124) );
  NOR4_X1 U668 ( .A1(n124), .A2(n367), .A3(n383), .A4(n207), .ZN(n125) );
  NAND3_X1 U669 ( .A1(n127), .A2(n126), .A3(n125), .ZN(n725) );
  INV_X1 U670 ( .A(n399), .ZN(n129) );
  INV_X1 U671 ( .A(n396), .ZN(n128) );
  NAND3_X1 U672 ( .A1(n26), .A2(n129), .A3(n128), .ZN(n132) );
  AOI211_X1 U673 ( .C1(z[11]), .C2(n156), .A(n400), .B(n398), .ZN(n130) );
  NAND4_X1 U674 ( .A1(n561), .A2(n565), .A3(n529), .A4(n130), .ZN(n131) );
  OR4_X1 U675 ( .A1(n391), .A2(n395), .A3(n132), .A4(n131), .ZN(n726) );
  INV_X1 U676 ( .A(n286), .ZN(n135) );
  INV_X1 U677 ( .A(n385), .ZN(n134) );
  INV_X1 U678 ( .A(n197), .ZN(n133) );
  NAND4_X1 U682 ( .A1(n135), .A2(n134), .A3(n133), .A4(n25), .ZN(n146) );
  INV_X1 U693 ( .A(z[12]), .ZN(n137) );
  OAI211_X1 U695 ( .C1(n213), .C2(n137), .A(n405), .B(n136), .ZN(n145) );
  AND3_X1 U714 ( .A1(n410), .A2(n406), .A3(n319), .ZN(n143) );
  INV_X1 U730 ( .A(n340), .ZN(n140) );
  INV_X1 U731 ( .A(n233), .ZN(n139) );
  INV_X1 U732 ( .A(n476), .ZN(n138) );
  NOR4_X1 U733 ( .A1(n141), .A2(n140), .A3(n139), .A4(n138), .ZN(n142) );
  NAND4_X1 U734 ( .A1(n475), .A2(n477), .A3(n143), .A4(n142), .ZN(n144) );
  OR3_X1 U735 ( .A1(n146), .A2(n145), .A3(n144), .ZN(n727) );
  INV_X1 U736 ( .A(n174), .ZN(n148) );
  INV_X1 U737 ( .A(n386), .ZN(n147) );
  NAND3_X1 U738 ( .A1(n148), .A2(n31), .A3(n147), .ZN(n154) );
  INV_X1 U739 ( .A(z[13]), .ZN(n151) );
  INV_X1 U740 ( .A(n485), .ZN(n150) );
  INV_X1 U741 ( .A(n486), .ZN(n149) );
  OAI221_X1 U742 ( .B1(n52), .B2(n151), .C1(n150), .C2(n149), .A(n302), .ZN(
        n152) );
  OR4_X1 U743 ( .A1(n478), .A2(n483), .A3(n496), .A4(n152), .ZN(n153) );
  OR4_X1 U744 ( .A1(n482), .A2(n487), .A3(n154), .A4(n153), .ZN(n728) );
  INV_X1 U745 ( .A(n325), .ZN(n435) );
  INV_X1 U746 ( .A(n507), .ZN(n758) );
  INV_X1 U747 ( .A(n467), .ZN(n155) );
  NOR3_X1 U748 ( .A1(n435), .A2(n758), .A3(n155), .ZN(n160) );
  AOI211_X1 U749 ( .C1(z[14]), .C2(n156), .A(n540), .B(n245), .ZN(n159) );
  NOR3_X1 U750 ( .A1(n546), .A2(n566), .A3(n175), .ZN(n158) );
  NOR3_X1 U751 ( .A1(n539), .A2(n344), .A3(n259), .ZN(n157) );
  NAND4_X1 U752 ( .A1(n160), .A2(n159), .A3(n158), .A4(n157), .ZN(n729) );
  OAI21_X1 U753 ( .B1(n17), .B2(n52), .A(n28), .ZN(n730) );
  OAI21_X1 U754 ( .B1(n16), .B2(n51), .A(n28), .ZN(n731) );
  OAI21_X1 U755 ( .B1(n15), .B2(n52), .A(n28), .ZN(n732) );
  OAI21_X1 U756 ( .B1(n14), .B2(n213), .A(n28), .ZN(n733) );
  OAI21_X1 U757 ( .B1(n13), .B2(n51), .A(n28), .ZN(n734) );
  OAI21_X1 U758 ( .B1(n12), .B2(n52), .A(n28), .ZN(n735) );
  OAI21_X1 U759 ( .B1(n11), .B2(n213), .A(n28), .ZN(n736) );
  OAI21_X1 U760 ( .B1(n10), .B2(n51), .A(n28), .ZN(n737) );
  OAI21_X1 U761 ( .B1(n9), .B2(n52), .A(n28), .ZN(n738) );
  OAI21_X1 U762 ( .B1(n8), .B2(n213), .A(n28), .ZN(n739) );
  OAI21_X1 U763 ( .B1(n7), .B2(n51), .A(n28), .ZN(n740) );
  OAI21_X1 U764 ( .B1(n6), .B2(n52), .A(n28), .ZN(n741) );
  OAI21_X1 U765 ( .B1(n5), .B2(n213), .A(n28), .ZN(n742) );
  OAI21_X1 U766 ( .B1(n4), .B2(n51), .A(n28), .ZN(n743) );
  INV_X1 U767 ( .A(n302), .ZN(n362) );
  INV_X1 U768 ( .A(n565), .ZN(n389) );
  INV_X1 U769 ( .A(n561), .ZN(n671) );
  INV_X1 U770 ( .A(n421), .ZN(n537) );
  INV_X1 U771 ( .A(n513), .ZN(n754) );
endmodule


module layer_13_16_1_32_B_rom ( clk, addr, z );
  input [3:0] addr;
  output [31:0] z;
  input clk;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n20, n21, n22, n23, n24, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n19,
         n25, n26, n27, n28, n29, n30, n31, n32, n33;

  NAND3_X1 U79 ( .A1(n49), .A2(n50), .A3(n44), .ZN(n35) );
  NAND3_X1 U80 ( .A1(n52), .A2(n53), .A3(n54), .ZN(n83) );
  NAND3_X1 U81 ( .A1(n64), .A2(n27), .A3(n65), .ZN(n88) );
  NAND3_X1 U82 ( .A1(n39), .A2(n55), .A3(n51), .ZN(n37) );
  NAND3_X1 U83 ( .A1(n77), .A2(addr[3]), .A3(addr[0]), .ZN(n67) );
  NAND3_X1 U84 ( .A1(addr[3]), .A2(n74), .A3(addr[0]), .ZN(n49) );
  NAND3_X1 U85 ( .A1(addr[2]), .A2(n75), .A3(addr[1]), .ZN(n59) );
  NAND3_X1 U86 ( .A1(addr[1]), .A2(addr[2]), .A3(n71), .ZN(n60) );
  DFF_X1 \z_reg[12]  ( .D(n25), .CK(clk), .Q(z[12]) );
  DFF_X1 \z_reg[3]  ( .D(n80), .CK(clk), .Q(z[3]) );
  DFF_X1 \z_reg[10]  ( .D(n87), .CK(clk), .Q(z[10]) );
  DFF_X1 \z_reg[11]  ( .D(n88), .CK(clk), .Q(z[11]) );
  DFF_X1 \z_reg[6]  ( .D(n83), .CK(clk), .Q(z[6]) );
  DFF_X1 \z_reg[7]  ( .D(n84), .CK(clk), .Q(z[7]) );
  DFF_X1 \z_reg[13]  ( .D(n89), .CK(clk), .Q(z[13]) );
  DFF_X1 \z_reg[0]  ( .D(n26), .CK(clk), .Q(z[0]) );
  DFF_X1 \z_reg[4]  ( .D(n81), .CK(clk), .Q(z[4]) );
  DFF_X1 \z_reg[30]  ( .D(n106), .CK(clk), .Q(z[30]), .QN(n2) );
  DFF_X1 \z_reg[29]  ( .D(n105), .CK(clk), .Q(z[29]), .QN(n3) );
  DFF_X1 \z_reg[28]  ( .D(n104), .CK(clk), .Q(z[28]), .QN(n4) );
  DFF_X1 \z_reg[27]  ( .D(n103), .CK(clk), .Q(z[27]), .QN(n5) );
  DFF_X1 \z_reg[26]  ( .D(n102), .CK(clk), .Q(z[26]), .QN(n6) );
  DFF_X1 \z_reg[25]  ( .D(n101), .CK(clk), .Q(z[25]), .QN(n7) );
  DFF_X1 \z_reg[14]  ( .D(n90), .CK(clk), .Q(z[14]), .QN(n18) );
  DFF_X1 \z_reg[9]  ( .D(n86), .CK(clk), .Q(z[9]), .QN(n20) );
  DFF_X1 \z_reg[8]  ( .D(n85), .CK(clk), .Q(z[8]), .QN(n21) );
  DFF_X1 \z_reg[2]  ( .D(n79), .CK(clk), .Q(z[2]), .QN(n23) );
  DFF_X1 \z_reg[1]  ( .D(n78), .CK(clk), .Q(z[1]), .QN(n24) );
  DFF_X1 \z_reg[31]  ( .D(n107), .CK(clk), .Q(z[31]), .QN(n1) );
  DFF_X1 \z_reg[24]  ( .D(n100), .CK(clk), .Q(z[24]), .QN(n8) );
  DFF_X1 \z_reg[23]  ( .D(n99), .CK(clk), .Q(z[23]), .QN(n9) );
  DFF_X1 \z_reg[22]  ( .D(n98), .CK(clk), .Q(z[22]), .QN(n10) );
  DFF_X1 \z_reg[21]  ( .D(n97), .CK(clk), .Q(z[21]), .QN(n11) );
  DFF_X1 \z_reg[20]  ( .D(n96), .CK(clk), .Q(z[20]), .QN(n12) );
  DFF_X1 \z_reg[19]  ( .D(n95), .CK(clk), .Q(z[19]), .QN(n13) );
  DFF_X1 \z_reg[18]  ( .D(n94), .CK(clk), .Q(z[18]), .QN(n14) );
  DFF_X1 \z_reg[17]  ( .D(n93), .CK(clk), .Q(z[17]), .QN(n15) );
  DFF_X1 \z_reg[16]  ( .D(n92), .CK(clk), .Q(z[16]), .QN(n16) );
  DFF_X1 \z_reg[15]  ( .D(n91), .CK(clk), .Q(z[15]), .QN(n17) );
  DFF_X1 \z_reg[5]  ( .D(n82), .CK(clk), .Q(z[5]), .QN(n22) );
  AND2_X1 U3 ( .A1(n68), .A2(n64), .ZN(n70) );
  NOR2_X1 U4 ( .A1(n28), .A2(n31), .ZN(n68) );
  AND2_X1 U5 ( .A1(n45), .A2(n40), .ZN(n53) );
  AND3_X1 U6 ( .A1(n38), .A2(n55), .A3(n40), .ZN(n42) );
  AND3_X1 U7 ( .A1(n40), .A2(n61), .A3(n56), .ZN(n64) );
  AND2_X1 U8 ( .A1(n58), .A2(n46), .ZN(n41) );
  AND4_X1 U9 ( .A1(n58), .A2(n53), .A3(n38), .A4(n62), .ZN(n51) );
  INV_X1 U10 ( .A(n48), .ZN(n27) );
  NAND2_X1 U11 ( .A1(n73), .A2(n74), .ZN(n38) );
  NAND2_X1 U12 ( .A1(n75), .A2(n74), .ZN(n45) );
  NAND4_X1 U13 ( .A1(n46), .A2(n59), .A3(n55), .A4(n45), .ZN(n36) );
  NAND2_X1 U14 ( .A1(n72), .A2(n75), .ZN(n55) );
  NAND2_X1 U15 ( .A1(n73), .A2(n72), .ZN(n46) );
  NAND2_X1 U16 ( .A1(n71), .A2(n72), .ZN(n62) );
  NAND2_X1 U17 ( .A1(n77), .A2(n73), .ZN(n61) );
  NAND2_X1 U18 ( .A1(n62), .A2(n67), .ZN(n48) );
  INV_X1 U19 ( .A(n60), .ZN(n28) );
  NAND2_X1 U20 ( .A1(n71), .A2(n74), .ZN(n40) );
  NAND2_X1 U21 ( .A1(n71), .A2(n77), .ZN(n44) );
  AND3_X1 U22 ( .A1(n59), .A2(n38), .A3(n44), .ZN(n56) );
  NAND2_X1 U23 ( .A1(n77), .A2(n75), .ZN(n50) );
  INV_X1 U24 ( .A(n49), .ZN(n31) );
  AND3_X1 U25 ( .A1(n60), .A2(n44), .A3(n46), .ZN(n39) );
  AND4_X1 U26 ( .A1(n59), .A2(n50), .A3(n49), .A4(n76), .ZN(n58) );
  AND2_X1 U27 ( .A1(n61), .A2(n67), .ZN(n76) );
  AND4_X1 U28 ( .A1(n46), .A2(n60), .A3(n61), .A4(n62), .ZN(n52) );
  NOR2_X1 U29 ( .A1(addr[2]), .A2(addr[1]), .ZN(n74) );
  NOR2_X1 U30 ( .A1(addr[3]), .A2(addr[0]), .ZN(n75) );
  NOR2_X1 U31 ( .A1(n32), .A2(addr[1]), .ZN(n72) );
  NOR2_X1 U32 ( .A1(n33), .A2(addr[0]), .ZN(n73) );
  OAI211_X1 U33 ( .C1(n37), .C2(n20), .A(n59), .B(n52), .ZN(n86) );
  NAND4_X1 U34 ( .A1(n42), .A2(n63), .A3(n60), .A4(n59), .ZN(n87) );
  NAND2_X1 U35 ( .A1(z[10]), .A2(n19), .ZN(n63) );
  AND2_X1 U36 ( .A1(addr[1]), .A2(n32), .ZN(n77) );
  AND2_X1 U37 ( .A1(addr[0]), .A2(n33), .ZN(n71) );
  OAI211_X1 U38 ( .C1(n37), .C2(n24), .A(n38), .B(n39), .ZN(n78) );
  OAI211_X1 U39 ( .C1(n37), .C2(n23), .A(n40), .B(n41), .ZN(n79) );
  OAI211_X1 U40 ( .C1(n37), .C2(n21), .A(n38), .B(n41), .ZN(n85) );
  OAI211_X1 U41 ( .C1(n37), .C2(n18), .A(n61), .B(n53), .ZN(n90) );
  OAI21_X1 U42 ( .B1(n37), .B2(n22), .A(n51), .ZN(n82) );
  OAI21_X1 U43 ( .B1(n37), .B2(n17), .A(n70), .ZN(n91) );
  OAI21_X1 U44 ( .B1(n37), .B2(n16), .A(n70), .ZN(n92) );
  OAI21_X1 U45 ( .B1(n37), .B2(n15), .A(n70), .ZN(n93) );
  OAI21_X1 U46 ( .B1(n37), .B2(n14), .A(n70), .ZN(n94) );
  OAI21_X1 U47 ( .B1(n37), .B2(n13), .A(n70), .ZN(n95) );
  OAI21_X1 U48 ( .B1(n37), .B2(n12), .A(n70), .ZN(n96) );
  OAI21_X1 U49 ( .B1(n37), .B2(n11), .A(n70), .ZN(n97) );
  OAI21_X1 U50 ( .B1(n37), .B2(n10), .A(n70), .ZN(n98) );
  OAI21_X1 U51 ( .B1(n37), .B2(n9), .A(n70), .ZN(n99) );
  OAI21_X1 U52 ( .B1(n37), .B2(n8), .A(n70), .ZN(n100) );
  OAI21_X1 U53 ( .B1(n37), .B2(n1), .A(n70), .ZN(n107) );
  NAND4_X1 U54 ( .A1(n38), .A2(n45), .A3(n46), .A4(n47), .ZN(n81) );
  AOI211_X1 U55 ( .C1(z[4]), .C2(n19), .A(n48), .B(n35), .ZN(n47) );
  OAI21_X1 U56 ( .B1(n37), .B2(n7), .A(n70), .ZN(n101) );
  OAI21_X1 U57 ( .B1(n37), .B2(n6), .A(n70), .ZN(n102) );
  OAI21_X1 U58 ( .B1(n37), .B2(n5), .A(n70), .ZN(n103) );
  OAI21_X1 U59 ( .B1(n37), .B2(n4), .A(n70), .ZN(n104) );
  OAI21_X1 U60 ( .B1(n37), .B2(n3), .A(n70), .ZN(n105) );
  OAI21_X1 U61 ( .B1(n37), .B2(n2), .A(n70), .ZN(n106) );
  NAND4_X1 U62 ( .A1(n68), .A2(n56), .A3(n69), .A4(n45), .ZN(n89) );
  NAND2_X1 U63 ( .A1(z[13]), .A2(n19), .ZN(n69) );
  NAND4_X1 U64 ( .A1(n42), .A2(n43), .A3(n44), .A4(n45), .ZN(n80) );
  NAND2_X1 U65 ( .A1(z[3]), .A2(n19), .ZN(n43) );
  NAND4_X1 U66 ( .A1(n56), .A2(n27), .A3(n57), .A4(n55), .ZN(n84) );
  NAND2_X1 U67 ( .A1(z[7]), .A2(n19), .ZN(n57) );
  INV_X1 U68 ( .A(addr[2]), .ZN(n32) );
  AOI211_X1 U69 ( .C1(z[11]), .C2(n19), .A(n30), .B(n28), .ZN(n65) );
  INV_X1 U70 ( .A(n50), .ZN(n30) );
  AOI211_X1 U71 ( .C1(z[6]), .C2(n19), .A(n29), .B(n31), .ZN(n54) );
  INV_X1 U72 ( .A(n55), .ZN(n29) );
  INV_X1 U73 ( .A(addr[3]), .ZN(n33) );
  INV_X1 U74 ( .A(n34), .ZN(n26) );
  AOI211_X1 U75 ( .C1(n19), .C2(z[0]), .A(n35), .B(n36), .ZN(n34) );
  INV_X1 U76 ( .A(n66), .ZN(n25) );
  AOI211_X1 U77 ( .C1(n19), .C2(z[12]), .A(n36), .B(n48), .ZN(n66) );
  INV_X1 U78 ( .A(n37), .ZN(n19) );
endmodule


module datapath_M13_N16_T32_DW_mult_tc_1 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n3, n6, n9, n12, n15, n18, n21, n24, n27, n30, n33, n36, n39, n42,
         n44, n48, n50, n53, n55, n58, n61, n63, n71, n74, n77, n79, n84, n86,
         n89, n91, n93, n95, n97, n99, n100, n102, n104, n105, n107, n109,
         n110, n112, n113, n114, n115, n116, n121, n127, n128, n130, n131,
         n132, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n151, n152, n154, n156, n158, n160,
         n161, n163, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n179, n180, n181, n182, n184, n187, n188, n189,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n203, n204,
         n205, n206, n213, n214, n215, n216, n217, n223, n224, n225, n226,
         n228, n231, n232, n233, n234, n238, n239, n240, n241, n242, n243,
         n244, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n261, n262, n263, n264, n269, n270, n271, n272, n274, n276,
         n277, n278, n279, n280, n281, n282, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n302, n304, n305, n306, n307, n308, n310, n312, n313, n314,
         n315, n316, n318, n320, n321, n322, n323, n324, n326, n328, n329,
         n331, n338, n344, n346, n350, n351, n352, n353, n354, n356, n358,
         n360, n363, n364, n365, n367, n369, n371, n372, n374, n375, n377,
         n378, n380, n382, n383, n384, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n824,
         n842, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1451, n1452, n1453, n1454, n1456, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1480, n1481, n1482, n1483,
         n1484, n1485, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938;
  assign n3 = a[1];
  assign n12 = a[3];
  assign n21 = a[5];
  assign n30 = a[7];
  assign n39 = a[9];
  assign n48 = a[11];
  assign n55 = a[13];
  assign n63 = a[15];
  assign n71 = a[17];
  assign n79 = a[19];
  assign n86 = a[21];
  assign n93 = a[23];
  assign n99 = a[25];
  assign n104 = a[27];
  assign n109 = a[29];
  assign n113 = a[31];
  assign n116 = b[0];
  assign n842 = a[0];
  assign n1427 = b[23];
  assign n1428 = b[22];
  assign n1429 = b[21];
  assign n1430 = b[20];
  assign n1431 = b[19];
  assign n1432 = b[18];
  assign n1433 = b[17];
  assign n1434 = b[16];
  assign n1435 = b[15];
  assign n1436 = b[14];
  assign n1437 = b[13];
  assign n1438 = b[12];
  assign n1439 = b[11];
  assign n1440 = b[10];
  assign n1441 = b[9];
  assign n1442 = b[8];
  assign n1443 = b[7];
  assign n1444 = b[6];
  assign n1445 = b[5];
  assign n1446 = b[4];
  assign n1447 = b[3];
  assign n1448 = b[2];
  assign n1449 = b[1];

  XOR2_X1 U378 ( .A(n378), .B(n371), .Z(n372) );
  XOR2_X1 U384 ( .A(n382), .B(n377), .Z(n378) );
  XOR2_X1 U390 ( .A(n970), .B(n383), .Z(n384) );
  XOR2_X1 U394 ( .A(n387), .B(n872), .Z(n388) );
  XOR2_X1 U396 ( .A(n860), .B(n389), .Z(n390) );
  FA_X1 U399 ( .A(n422), .B(n397), .CI(n395), .CO(n392), .S(n393) );
  FA_X1 U400 ( .A(n399), .B(n401), .CI(n424), .CO(n394), .S(n395) );
  FA_X1 U401 ( .A(n428), .B(n403), .CI(n426), .CO(n396), .S(n397) );
  FA_X1 U402 ( .A(n430), .B(n407), .CI(n405), .CO(n398), .S(n399) );
  FA_X1 U403 ( .A(n432), .B(n434), .CI(n409), .CO(n400), .S(n401) );
  FA_X1 U404 ( .A(n413), .B(n436), .CI(n411), .CO(n402), .S(n403) );
  FA_X1 U405 ( .A(n417), .B(n419), .CI(n415), .CO(n404), .S(n405) );
  FA_X1 U406 ( .A(n440), .B(n442), .CI(n438), .CO(n406), .S(n407) );
  FA_X1 U407 ( .A(n446), .B(n1017), .CI(n444), .CO(n408), .S(n409) );
  FA_X1 U408 ( .A(n1043), .B(n971), .CI(n1071), .CO(n410), .S(n411) );
  FA_X1 U409 ( .A(n993), .B(n917), .CI(n1101), .CO(n412), .S(n413) );
  FA_X1 U410 ( .A(n891), .B(n881), .CI(n951), .CO(n414), .S(n415) );
  FA_X1 U411 ( .A(n903), .B(n873), .CI(n933), .CO(n416), .S(n417) );
  FA_X1 U412 ( .A(n863), .B(n861), .CI(n867), .CO(n418), .S(n419) );
  FA_X1 U413 ( .A(n450), .B(n425), .CI(n423), .CO(n420), .S(n421) );
  FA_X1 U414 ( .A(n427), .B(n454), .CI(n452), .CO(n422), .S(n423) );
  FA_X1 U415 ( .A(n431), .B(n456), .CI(n429), .CO(n424), .S(n425) );
  FA_X1 U416 ( .A(n458), .B(n435), .CI(n433), .CO(n426), .S(n427) );
  FA_X1 U417 ( .A(n437), .B(n462), .CI(n460), .CO(n428), .S(n429) );
  FA_X1 U418 ( .A(n439), .B(n443), .CI(n441), .CO(n430), .S(n431) );
  FA_X1 U419 ( .A(n466), .B(n464), .CI(n445), .CO(n432), .S(n433) );
  FA_X1 U420 ( .A(n470), .B(n472), .CI(n468), .CO(n434), .S(n435) );
  FA_X1 U421 ( .A(n1018), .B(n972), .CI(n447), .CO(n436), .S(n437) );
  FA_X1 U422 ( .A(n1044), .B(n952), .CI(n1072), .CO(n438), .S(n439) );
  FA_X1 U423 ( .A(n918), .B(n994), .CI(n1102), .CO(n440), .S(n441) );
  FA_X1 U424 ( .A(n892), .B(n874), .CI(n934), .CO(n442), .S(n443) );
  FA_X1 U425 ( .A(n882), .B(n868), .CI(n904), .CO(n444), .S(n445) );
  HA_X1 U426 ( .A(n864), .B(n845), .CO(n446), .S(n447) );
  FA_X1 U428 ( .A(n455), .B(n457), .CI(n478), .CO(n450), .S(n451) );
  FA_X1 U429 ( .A(n459), .B(n482), .CI(n480), .CO(n452), .S(n453) );
  FA_X1 U430 ( .A(n484), .B(n463), .CI(n461), .CO(n454), .S(n455) );
  FA_X1 U431 ( .A(n488), .B(n465), .CI(n486), .CO(n456), .S(n457) );
  FA_X1 U432 ( .A(n469), .B(n471), .CI(n467), .CO(n458), .S(n459) );
  FA_X1 U433 ( .A(n490), .B(n492), .CI(n473), .CO(n460), .S(n461) );
  FA_X1 U434 ( .A(n494), .B(n498), .CI(n496), .CO(n462), .S(n463) );
  FA_X1 U435 ( .A(n1019), .B(n973), .CI(n1073), .CO(n464), .S(n465) );
  FA_X1 U436 ( .A(n1045), .B(n935), .CI(n1103), .CO(n466), .S(n467) );
  FA_X1 U437 ( .A(n919), .B(n893), .CI(n995), .CO(n468), .S(n469) );
  FA_X1 U438 ( .A(n905), .B(n883), .CI(n953), .CO(n470), .S(n471) );
  FA_X1 U439 ( .A(n875), .B(n865), .CI(n869), .CO(n472), .S(n473) );
  FA_X1 U440 ( .A(n502), .B(n479), .CI(n477), .CO(n474), .S(n475) );
  FA_X1 U441 ( .A(n483), .B(n481), .CI(n504), .CO(n476), .S(n477) );
  FA_X1 U443 ( .A(n510), .B(n489), .CI(n487), .CO(n480), .S(n481) );
  FA_X1 U444 ( .A(n491), .B(n493), .CI(n512), .CO(n482), .S(n483) );
  FA_X1 U445 ( .A(n497), .B(n514), .CI(n495), .CO(n484), .S(n485) );
  FA_X1 U446 ( .A(n518), .B(n520), .CI(n516), .CO(n486), .S(n487) );
  FA_X1 U447 ( .A(n522), .B(n1020), .CI(n499), .CO(n488), .S(n489) );
  FA_X1 U448 ( .A(n1074), .B(n1046), .CI(n974), .CO(n490), .S(n491) );
  FA_X1 U449 ( .A(n1104), .B(n920), .CI(n996), .CO(n492), .S(n493) );
  FA_X1 U450 ( .A(n894), .B(n884), .CI(n954), .CO(n494), .S(n495) );
  FA_X1 U451 ( .A(n906), .B(n876), .CI(n936), .CO(n496), .S(n497) );
  HA_X1 U452 ( .A(n870), .B(n846), .CO(n498), .S(n499) );
  FA_X1 U454 ( .A(n507), .B(n530), .CI(n528), .CO(n502), .S(n503) );
  FA_X1 U455 ( .A(n511), .B(n532), .CI(n509), .CO(n504), .S(n505) );
  FA_X1 U456 ( .A(n513), .B(n536), .CI(n534), .CO(n506), .S(n507) );
  FA_X1 U457 ( .A(n517), .B(n519), .CI(n515), .CO(n508), .S(n509) );
  FA_X1 U458 ( .A(n523), .B(n538), .CI(n521), .CO(n510), .S(n511) );
  FA_X1 U459 ( .A(n544), .B(n542), .CI(n540), .CO(n512), .S(n513) );
  FA_X1 U460 ( .A(n1021), .B(n546), .CI(n975), .CO(n514), .S(n515) );
  FA_X1 U461 ( .A(n1047), .B(n955), .CI(n1105), .CO(n516), .S(n517) );
  FA_X1 U462 ( .A(n907), .B(n937), .CI(n1075), .CO(n518), .S(n519) );
  FA_X1 U463 ( .A(n921), .B(n895), .CI(n997), .CO(n520), .S(n521) );
  FA_X1 U464 ( .A(n885), .B(n871), .CI(n877), .CO(n522), .S(n523) );
  FA_X1 U465 ( .A(n550), .B(n529), .CI(n527), .CO(n524), .S(n525) );
  FA_X1 U466 ( .A(n531), .B(n554), .CI(n552), .CO(n526), .S(n527) );
  FA_X1 U467 ( .A(n535), .B(n556), .CI(n533), .CO(n528), .S(n529) );
  FA_X1 U468 ( .A(n558), .B(n560), .CI(n537), .CO(n530), .S(n531) );
  FA_X1 U469 ( .A(n541), .B(n543), .CI(n539), .CO(n532), .S(n533) );
  FA_X1 U470 ( .A(n562), .B(n564), .CI(n545), .CO(n534), .S(n535) );
  FA_X1 U471 ( .A(n568), .B(n547), .CI(n566), .CO(n536), .S(n537) );
  FA_X1 U473 ( .A(n1048), .B(n938), .CI(n1106), .CO(n540), .S(n541) );
  FA_X1 U474 ( .A(n922), .B(n896), .CI(n998), .CO(n542), .S(n543) );
  FA_X1 U475 ( .A(n908), .B(n886), .CI(n956), .CO(n544), .S(n545) );
  HA_X1 U476 ( .A(n878), .B(n847), .CO(n546), .S(n547) );
  FA_X1 U478 ( .A(n555), .B(n557), .CI(n574), .CO(n550), .S(n551) );
  FA_X1 U479 ( .A(n559), .B(n578), .CI(n576), .CO(n552), .S(n553) );
  FA_X1 U480 ( .A(n580), .B(n582), .CI(n561), .CO(n554), .S(n555) );
  FA_X1 U481 ( .A(n565), .B(n567), .CI(n563), .CO(n556), .S(n557) );
  FA_X1 U482 ( .A(n584), .B(n586), .CI(n569), .CO(n558), .S(n559) );
  FA_X1 U483 ( .A(n590), .B(n977), .CI(n588), .CO(n560), .S(n561) );
  FA_X1 U484 ( .A(n1023), .B(n957), .CI(n1049), .CO(n562), .S(n563) );
  FA_X1 U485 ( .A(n999), .B(n923), .CI(n1107), .CO(n564), .S(n565) );
  FA_X1 U486 ( .A(n939), .B(n909), .CI(n1077), .CO(n566), .S(n567) );
  FA_X1 U487 ( .A(n887), .B(n879), .CI(n897), .CO(n568), .S(n569) );
  FA_X1 U490 ( .A(n581), .B(n600), .CI(n598), .CO(n574), .S(n575) );
  FA_X1 U491 ( .A(n602), .B(n585), .CI(n583), .CO(n576), .S(n577) );
  FA_X1 U492 ( .A(n589), .B(n606), .CI(n587), .CO(n578), .S(n579) );
  FA_X1 U493 ( .A(n608), .B(n610), .CI(n604), .CO(n580), .S(n581) );
  FA_X1 U494 ( .A(n1024), .B(n978), .CI(n591), .CO(n582), .S(n583) );
  FA_X1 U495 ( .A(n958), .B(n1050), .CI(n1108), .CO(n584), .S(n585) );
  FA_X1 U496 ( .A(n940), .B(n910), .CI(n1078), .CO(n586), .S(n587) );
  FA_X1 U497 ( .A(n924), .B(n898), .CI(n1000), .CO(n588), .S(n589) );
  HA_X1 U498 ( .A(n888), .B(n848), .CO(n590), .S(n591) );
  FA_X1 U499 ( .A(n614), .B(n597), .CI(n595), .CO(n592), .S(n593) );
  FA_X1 U500 ( .A(n599), .B(n601), .CI(n616), .CO(n594), .S(n595) );
  FA_X1 U501 ( .A(n620), .B(n603), .CI(n618), .CO(n596), .S(n597) );
  FA_X1 U502 ( .A(n605), .B(n607), .CI(n622), .CO(n598), .S(n599) );
  FA_X1 U503 ( .A(n611), .B(n624), .CI(n609), .CO(n600), .S(n601) );
  FA_X1 U505 ( .A(n979), .B(n959), .CI(n1025), .CO(n604), .S(n605) );
  FA_X1 U506 ( .A(n1051), .B(n941), .CI(n1079), .CO(n606), .S(n607) );
  FA_X1 U507 ( .A(n1001), .B(n925), .CI(n1109), .CO(n608), .S(n609) );
  FA_X1 U508 ( .A(n899), .B(n889), .CI(n911), .CO(n610), .S(n611) );
  FA_X1 U510 ( .A(n619), .B(n621), .CI(n636), .CO(n614), .S(n615) );
  FA_X1 U511 ( .A(n623), .B(n640), .CI(n638), .CO(n616), .S(n617) );
  FA_X1 U513 ( .A(n646), .B(n644), .CI(n642), .CO(n620), .S(n621) );
  FA_X1 U514 ( .A(n631), .B(n980), .CI(n648), .CO(n622), .S(n623) );
  FA_X1 U515 ( .A(n1026), .B(n1052), .CI(n960), .CO(n624), .S(n625) );
  FA_X1 U516 ( .A(n1110), .B(n926), .CI(n1002), .CO(n626), .S(n627) );
  HA_X1 U518 ( .A(n900), .B(n849), .CO(n630), .S(n631) );
  FA_X1 U520 ( .A(n639), .B(n641), .CI(n654), .CO(n634), .S(n635) );
  FA_X1 U521 ( .A(n658), .B(n643), .CI(n656), .CO(n636), .S(n637) );
  FA_X1 U524 ( .A(n981), .B(n1003), .CI(n666), .CO(n642), .S(n643) );
  FA_X1 U525 ( .A(n1027), .B(n961), .CI(n1081), .CO(n644), .S(n645) );
  FA_X1 U526 ( .A(n1111), .B(n943), .CI(n1053), .CO(n646), .S(n647) );
  FA_X1 U529 ( .A(n657), .B(n659), .CI(n672), .CO(n652), .S(n653) );
  FA_X1 U530 ( .A(n676), .B(n661), .CI(n674), .CO(n654), .S(n655) );
  FA_X1 U531 ( .A(n663), .B(n680), .CI(n665), .CO(n656), .S(n657) );
  FA_X1 U532 ( .A(n682), .B(n667), .CI(n678), .CO(n658), .S(n659) );
  FA_X1 U533 ( .A(n1028), .B(n962), .CI(n982), .CO(n660), .S(n661) );
  FA_X1 U534 ( .A(n1054), .B(n944), .CI(n1082), .CO(n662), .S(n663) );
  FA_X1 U535 ( .A(n928), .B(n1004), .CI(n1112), .CO(n664), .S(n665) );
  HA_X1 U536 ( .A(n850), .B(n914), .CO(n666), .S(n667) );
  FA_X1 U538 ( .A(n675), .B(n677), .CI(n688), .CO(n670), .S(n671) );
  FA_X1 U539 ( .A(n692), .B(n679), .CI(n690), .CO(n672), .S(n673) );
  FA_X1 U540 ( .A(n683), .B(n696), .CI(n681), .CO(n674), .S(n675) );
  FA_X1 U541 ( .A(n698), .B(n1005), .CI(n694), .CO(n676), .S(n677) );
  FA_X1 U542 ( .A(n1029), .B(n1055), .CI(n983), .CO(n678), .S(n679) );
  FA_X1 U543 ( .A(n1113), .B(n1083), .CI(n963), .CO(n680), .S(n681) );
  FA_X1 U544 ( .A(n929), .B(n915), .CI(n945), .CO(n682), .S(n683) );
  FA_X1 U545 ( .A(n689), .B(n702), .CI(n687), .CO(n684), .S(n685) );
  FA_X1 U546 ( .A(n691), .B(n693), .CI(n704), .CO(n686), .S(n687) );
  FA_X1 U547 ( .A(n695), .B(n697), .CI(n706), .CO(n688), .S(n689) );
  FA_X1 U548 ( .A(n712), .B(n708), .CI(n710), .CO(n690), .S(n691) );
  FA_X1 U549 ( .A(n1006), .B(n984), .CI(n699), .CO(n692), .S(n693) );
  FA_X1 U550 ( .A(n1030), .B(n964), .CI(n1084), .CO(n694), .S(n695) );
  FA_X1 U551 ( .A(n1056), .B(n946), .CI(n1114), .CO(n696), .S(n697) );
  HA_X1 U552 ( .A(n930), .B(n851), .CO(n698), .S(n699) );
  FA_X1 U553 ( .A(n716), .B(n705), .CI(n703), .CO(n700), .S(n701) );
  FA_X1 U554 ( .A(n707), .B(n720), .CI(n718), .CO(n702), .S(n703) );
  FA_X1 U555 ( .A(n711), .B(n713), .CI(n709), .CO(n704), .S(n705) );
  FA_X1 U556 ( .A(n722), .B(n726), .CI(n724), .CO(n706), .S(n707) );
  FA_X1 U557 ( .A(n1031), .B(n1057), .CI(n1007), .CO(n708), .S(n709) );
  FA_X1 U558 ( .A(n1085), .B(n1115), .CI(n985), .CO(n710), .S(n711) );
  FA_X1 U559 ( .A(n965), .B(n931), .CI(n947), .CO(n712), .S(n713) );
  FA_X1 U561 ( .A(n721), .B(n723), .CI(n732), .CO(n716), .S(n717) );
  FA_X1 U562 ( .A(n734), .B(n736), .CI(n725), .CO(n718), .S(n719) );
  FA_X1 U563 ( .A(n727), .B(n1008), .CI(n738), .CO(n720), .S(n721) );
  FA_X1 U565 ( .A(n1116), .B(n966), .CI(n1086), .CO(n724), .S(n725) );
  HA_X1 U566 ( .A(n948), .B(n852), .CO(n726), .S(n727) );
  FA_X1 U568 ( .A(n735), .B(n737), .CI(n744), .CO(n730), .S(n731) );
  FA_X1 U569 ( .A(n748), .B(n746), .CI(n739), .CO(n732), .S(n733) );
  FA_X1 U570 ( .A(n1059), .B(n1033), .CI(n750), .CO(n734), .S(n735) );
  FA_X1 U571 ( .A(n1117), .B(n1087), .CI(n1009), .CO(n736), .S(n737) );
  FA_X1 U572 ( .A(n967), .B(n949), .CI(n987), .CO(n738), .S(n739) );
  FA_X1 U573 ( .A(n754), .B(n745), .CI(n743), .CO(n740), .S(n741) );
  FA_X1 U574 ( .A(n747), .B(n749), .CI(n756), .CO(n742), .S(n743) );
  FA_X1 U575 ( .A(n760), .B(n751), .CI(n758), .CO(n744), .S(n745) );
  FA_X1 U576 ( .A(n1034), .B(n1060), .CI(n1010), .CO(n746), .S(n747) );
  FA_X1 U577 ( .A(n1088), .B(n1118), .CI(n988), .CO(n748), .S(n749) );
  HA_X1 U578 ( .A(n968), .B(n853), .CO(n750), .S(n751) );
  FA_X1 U579 ( .A(n757), .B(n764), .CI(n755), .CO(n752), .S(n753) );
  FA_X1 U580 ( .A(n759), .B(n761), .CI(n766), .CO(n754), .S(n755) );
  FA_X1 U581 ( .A(n770), .B(n1061), .CI(n768), .CO(n756), .S(n757) );
  FA_X1 U582 ( .A(n1089), .B(n1035), .CI(n1119), .CO(n758), .S(n759) );
  FA_X1 U583 ( .A(n1011), .B(n969), .CI(n989), .CO(n760), .S(n761) );
  FA_X1 U584 ( .A(n774), .B(n767), .CI(n765), .CO(n762), .S(n763) );
  FA_X1 U585 ( .A(n776), .B(n778), .CI(n769), .CO(n764), .S(n765) );
  FA_X1 U586 ( .A(n1062), .B(n1036), .CI(n771), .CO(n766), .S(n767) );
  FA_X1 U587 ( .A(n1090), .B(n1012), .CI(n1120), .CO(n768), .S(n769) );
  HA_X1 U588 ( .A(n990), .B(n854), .CO(n770), .S(n771) );
  FA_X1 U589 ( .A(n782), .B(n777), .CI(n775), .CO(n772), .S(n773) );
  FA_X1 U590 ( .A(n784), .B(n786), .CI(n779), .CO(n774), .S(n775) );
  FA_X1 U591 ( .A(n1091), .B(n1063), .CI(n1121), .CO(n776), .S(n777) );
  FA_X1 U592 ( .A(n1013), .B(n991), .CI(n1037), .CO(n778), .S(n779) );
  FA_X1 U593 ( .A(n785), .B(n790), .CI(n783), .CO(n780), .S(n781) );
  FA_X1 U594 ( .A(n787), .B(n1064), .CI(n792), .CO(n782), .S(n783) );
  FA_X1 U595 ( .A(n1092), .B(n1038), .CI(n1122), .CO(n784), .S(n785) );
  HA_X1 U596 ( .A(n1014), .B(n855), .CO(n786), .S(n787) );
  FA_X1 U597 ( .A(n793), .B(n796), .CI(n791), .CO(n788), .S(n789) );
  FA_X1 U598 ( .A(n1123), .B(n1093), .CI(n798), .CO(n790), .S(n791) );
  FA_X1 U599 ( .A(n1039), .B(n1015), .CI(n1065), .CO(n792), .S(n793) );
  FA_X1 U600 ( .A(n802), .B(n799), .CI(n797), .CO(n794), .S(n795) );
  FA_X1 U601 ( .A(n1094), .B(n1066), .CI(n1124), .CO(n796), .S(n797) );
  HA_X1 U602 ( .A(n1040), .B(n856), .CO(n798), .S(n799) );
  FA_X1 U603 ( .A(n806), .B(n1125), .CI(n803), .CO(n800), .S(n801) );
  FA_X1 U604 ( .A(n1067), .B(n1041), .CI(n1095), .CO(n802), .S(n803) );
  FA_X1 U605 ( .A(n1126), .B(n1096), .CI(n807), .CO(n804), .S(n805) );
  HA_X1 U606 ( .A(n1068), .B(n857), .CO(n806), .S(n807) );
  FA_X1 U607 ( .A(n1097), .B(n1069), .CI(n1127), .CO(n808), .S(n809) );
  HA_X1 U608 ( .A(n1098), .B(n858), .CO(n810), .S(n811) );
  OR2_X2 U1312 ( .A1(n1847), .A2(n1848), .ZN(n1722) );
  OAI21_X1 U1313 ( .B1(n193), .B2(n187), .A(n188), .ZN(n1588) );
  BUF_X1 U1314 ( .A(n1723), .Z(n1589) );
  CLKBUF_X1 U1315 ( .A(n1848), .Z(n1590) );
  CLKBUF_X3 U1316 ( .A(n1932), .Z(n1591) );
  CLKBUF_X3 U1317 ( .A(n1932), .Z(n1592) );
  INV_X1 U1318 ( .A(n818), .ZN(n1593) );
  CLKBUF_X1 U1319 ( .A(n1680), .Z(n1594) );
  NAND2_X1 U1320 ( .A1(n1790), .A2(n1791), .ZN(n1595) );
  INV_X1 U1321 ( .A(n1924), .ZN(n1596) );
  NOR2_X1 U1322 ( .A1(n741), .A2(n752), .ZN(n1597) );
  NOR2_X1 U1323 ( .A1(n741), .A2(n752), .ZN(n1598) );
  NOR2_X1 U1324 ( .A1(n741), .A2(n752), .ZN(n280) );
  CLKBUF_X1 U1325 ( .A(n278), .Z(n1727) );
  BUF_X2 U1326 ( .A(n9), .Z(n1913) );
  BUF_X2 U1327 ( .A(n9), .Z(n1717) );
  INV_X1 U1328 ( .A(n217), .ZN(n1599) );
  INV_X1 U1329 ( .A(n1766), .ZN(n1600) );
  OR2_X2 U1330 ( .A1(n633), .A2(n650), .ZN(n1662) );
  NAND2_X1 U1331 ( .A1(n1461), .A2(n1888), .ZN(n1601) );
  CLKBUF_X1 U1332 ( .A(n1449), .Z(n1602) );
  BUF_X4 U1333 ( .A(n1449), .Z(n1603) );
  XNOR2_X1 U1334 ( .A(n1604), .B(n596), .ZN(n573) );
  XNOR2_X1 U1335 ( .A(n577), .B(n579), .ZN(n1604) );
  XNOR2_X1 U1336 ( .A(n1605), .B(n573), .ZN(n571) );
  XNOR2_X1 U1337 ( .A(n594), .B(n575), .ZN(n1605) );
  XNOR2_X1 U1338 ( .A(n653), .B(n1606), .ZN(n651) );
  XNOR2_X1 U1339 ( .A(n670), .B(n655), .ZN(n1606) );
  FA_X1 U1340 ( .A(n502), .B(n479), .CI(n477), .S(n1607) );
  NAND2_X1 U1341 ( .A1(n1595), .A2(n100), .ZN(n1608) );
  NAND2_X1 U1342 ( .A1(n58), .A2(n1460), .ZN(n1609) );
  OAI22_X1 U1343 ( .A1(n1867), .A2(n1798), .B1(n1267), .B2(n1889), .ZN(n1610)
         );
  XOR2_X1 U1344 ( .A(n652), .B(n637), .Z(n1611) );
  XOR2_X1 U1345 ( .A(n635), .B(n1611), .Z(n633) );
  NAND2_X1 U1346 ( .A1(n635), .A2(n652), .ZN(n1612) );
  NAND2_X1 U1347 ( .A1(n635), .A2(n637), .ZN(n1613) );
  NAND2_X1 U1348 ( .A1(n652), .A2(n637), .ZN(n1614) );
  NAND3_X1 U1349 ( .A1(n1612), .A2(n1613), .A3(n1614), .ZN(n632) );
  INV_X1 U1350 ( .A(n223), .ZN(n1615) );
  CLKBUF_X1 U1351 ( .A(a[12]), .Z(n1721) );
  BUF_X1 U1352 ( .A(n77), .Z(n1758) );
  XNOR2_X1 U1353 ( .A(n1616), .B(n649), .ZN(n639) );
  XNOR2_X1 U1354 ( .A(n647), .B(n645), .ZN(n1616) );
  CLKBUF_X1 U1355 ( .A(n1877), .Z(n1617) );
  BUF_X1 U1356 ( .A(n1877), .Z(n1618) );
  CLKBUF_X1 U1357 ( .A(n1877), .Z(n1619) );
  XNOR2_X1 U1358 ( .A(n1935), .B(n1721), .ZN(n1877) );
  BUF_X4 U1359 ( .A(n36), .Z(n1896) );
  BUF_X1 U1360 ( .A(n179), .Z(n1620) );
  NAND2_X1 U1361 ( .A1(n577), .A2(n579), .ZN(n1621) );
  NAND2_X1 U1362 ( .A1(n577), .A2(n596), .ZN(n1622) );
  NAND2_X1 U1363 ( .A1(n579), .A2(n596), .ZN(n1623) );
  NAND3_X1 U1364 ( .A1(n1621), .A2(n1622), .A3(n1623), .ZN(n572) );
  NAND2_X1 U1365 ( .A1(n594), .A2(n575), .ZN(n1624) );
  NAND2_X1 U1366 ( .A1(n594), .A2(n573), .ZN(n1625) );
  NAND2_X1 U1367 ( .A1(n575), .A2(n573), .ZN(n1626) );
  NAND3_X1 U1368 ( .A1(n1624), .A2(n1625), .A3(n1626), .ZN(n570) );
  NAND2_X1 U1369 ( .A1(n1456), .A2(n1823), .ZN(n1627) );
  CLKBUF_X1 U1370 ( .A(n112), .Z(n1628) );
  NAND2_X2 U1371 ( .A1(n1453), .A2(n1703), .ZN(n107) );
  XOR2_X1 U1372 ( .A(n742), .B(n733), .Z(n1629) );
  XOR2_X1 U1373 ( .A(n731), .B(n1629), .Z(n729) );
  NAND2_X1 U1374 ( .A1(n731), .A2(n742), .ZN(n1630) );
  NAND2_X1 U1375 ( .A1(n731), .A2(n733), .ZN(n1631) );
  NAND2_X1 U1376 ( .A1(n742), .A2(n733), .ZN(n1632) );
  NAND3_X1 U1377 ( .A1(n1630), .A2(n1631), .A3(n1632), .ZN(n728) );
  CLKBUF_X1 U1378 ( .A(a[12]), .Z(n1633) );
  NAND2_X2 U1379 ( .A1(n1763), .A2(n1823), .ZN(n1787) );
  BUF_X2 U1380 ( .A(n1876), .Z(n1719) );
  INV_X1 U1381 ( .A(n1889), .ZN(n1634) );
  BUF_X2 U1382 ( .A(n55), .Z(n1858) );
  INV_X1 U1383 ( .A(n284), .ZN(n1635) );
  XOR2_X1 U1384 ( .A(n927), .B(n901), .Z(n1636) );
  XOR2_X1 U1385 ( .A(n1636), .B(n913), .Z(n649) );
  NAND2_X1 U1386 ( .A1(n927), .A2(n901), .ZN(n1637) );
  NAND2_X1 U1387 ( .A1(n927), .A2(n913), .ZN(n1638) );
  NAND2_X1 U1388 ( .A1(n901), .A2(n913), .ZN(n1639) );
  NAND3_X1 U1389 ( .A1(n1637), .A2(n1638), .A3(n1639), .ZN(n648) );
  NAND2_X1 U1390 ( .A1(n647), .A2(n645), .ZN(n1640) );
  NAND2_X1 U1391 ( .A1(n647), .A2(n649), .ZN(n1641) );
  NAND2_X1 U1392 ( .A1(n645), .A2(n649), .ZN(n1642) );
  NAND3_X1 U1393 ( .A1(n1640), .A2(n1641), .A3(n1642), .ZN(n638) );
  INV_X1 U1394 ( .A(n1762), .ZN(n1937) );
  XNOR2_X1 U1395 ( .A(n503), .B(n1643), .ZN(n501) );
  XNOR2_X1 U1396 ( .A(n526), .B(n505), .ZN(n1643) );
  INV_X1 U1397 ( .A(n1694), .ZN(n1644) );
  XOR2_X1 U1398 ( .A(n485), .B(n508), .Z(n1645) );
  XOR2_X1 U1399 ( .A(n506), .B(n1645), .Z(n479) );
  NAND2_X1 U1400 ( .A1(n506), .A2(n485), .ZN(n1646) );
  NAND2_X1 U1401 ( .A1(n506), .A2(n508), .ZN(n1647) );
  NAND2_X1 U1402 ( .A1(n485), .A2(n508), .ZN(n1648) );
  NAND3_X1 U1403 ( .A1(n1646), .A2(n1647), .A3(n1648), .ZN(n478) );
  CLKBUF_X1 U1404 ( .A(n986), .Z(n1731) );
  INV_X1 U1405 ( .A(n1714), .ZN(n1649) );
  AND2_X1 U1406 ( .A1(n571), .A2(n592), .ZN(n1833) );
  AND2_X1 U1407 ( .A1(n549), .A2(n570), .ZN(n1650) );
  INV_X4 U1408 ( .A(n1650), .ZN(n203) );
  NAND2_X1 U1409 ( .A1(n653), .A2(n670), .ZN(n1651) );
  NAND2_X1 U1410 ( .A1(n653), .A2(n655), .ZN(n1652) );
  NAND2_X1 U1411 ( .A1(n670), .A2(n655), .ZN(n1653) );
  NAND3_X1 U1412 ( .A1(n1651), .A2(n1652), .A3(n1653), .ZN(n650) );
  BUF_X1 U1413 ( .A(n1818), .Z(n1730) );
  BUF_X1 U1414 ( .A(n1601), .Z(n1867) );
  XOR2_X1 U1415 ( .A(n912), .B(n942), .Z(n1654) );
  XOR2_X1 U1416 ( .A(n1654), .B(n1080), .Z(n629) );
  XOR2_X1 U1417 ( .A(n627), .B(n625), .Z(n1655) );
  XOR2_X1 U1418 ( .A(n1655), .B(n629), .Z(n619) );
  NAND2_X1 U1419 ( .A1(n942), .A2(n912), .ZN(n1656) );
  NAND2_X1 U1420 ( .A1(n942), .A2(n1080), .ZN(n1657) );
  NAND2_X1 U1421 ( .A1(n912), .A2(n1080), .ZN(n1658) );
  NAND3_X1 U1422 ( .A1(n1656), .A2(n1657), .A3(n1658), .ZN(n628) );
  NAND2_X1 U1423 ( .A1(n627), .A2(n625), .ZN(n1659) );
  NAND2_X1 U1424 ( .A1(n627), .A2(n629), .ZN(n1660) );
  NAND2_X1 U1425 ( .A1(n625), .A2(n629), .ZN(n1661) );
  NAND3_X1 U1426 ( .A1(n1659), .A2(n1660), .A3(n1661), .ZN(n618) );
  CLKBUF_X3 U1427 ( .A(n27), .Z(n1902) );
  BUF_X1 U1428 ( .A(n61), .Z(n1855) );
  FA_X1 U1429 ( .A(n455), .B(n457), .CI(n478), .S(n1663) );
  INV_X1 U1430 ( .A(n1895), .ZN(n1664) );
  INV_X1 U1431 ( .A(n1895), .ZN(n1665) );
  INV_X1 U1432 ( .A(n1895), .ZN(n1893) );
  INV_X2 U1433 ( .A(n12), .ZN(n1924) );
  CLKBUF_X1 U1434 ( .A(a[18]), .Z(n1666) );
  CLKBUF_X1 U1435 ( .A(n93), .Z(n1667) );
  INV_X1 U1436 ( .A(n216), .ZN(n1668) );
  CLKBUF_X3 U1437 ( .A(n71), .Z(n1863) );
  CLKBUF_X3 U1438 ( .A(n55), .Z(n1859) );
  CLKBUF_X3 U1439 ( .A(n1932), .Z(n1860) );
  INV_X1 U1440 ( .A(n42), .ZN(n1669) );
  CLKBUF_X1 U1441 ( .A(n270), .Z(n1670) );
  CLKBUF_X3 U1442 ( .A(n44), .Z(n1733) );
  BUF_X1 U1443 ( .A(n95), .Z(n1706) );
  XOR2_X1 U1444 ( .A(n730), .B(n719), .Z(n1671) );
  XOR2_X1 U1445 ( .A(n717), .B(n1671), .Z(n715) );
  NAND2_X1 U1446 ( .A1(n717), .A2(n730), .ZN(n1672) );
  NAND2_X1 U1447 ( .A1(n717), .A2(n719), .ZN(n1673) );
  NAND2_X1 U1448 ( .A1(n730), .A2(n719), .ZN(n1674) );
  NAND3_X1 U1449 ( .A1(n1672), .A2(n1673), .A3(n1674), .ZN(n714) );
  NAND2_X1 U1450 ( .A1(n503), .A2(n526), .ZN(n1675) );
  NAND2_X1 U1451 ( .A1(n503), .A2(n505), .ZN(n1676) );
  NAND2_X1 U1452 ( .A1(n526), .A2(n505), .ZN(n1677) );
  NAND3_X1 U1453 ( .A1(n1675), .A2(n1676), .A3(n1677), .ZN(n500) );
  INV_X1 U1454 ( .A(n1911), .ZN(n1678) );
  INV_X1 U1455 ( .A(n1911), .ZN(n1910) );
  FA_X1 U1456 ( .A(n555), .B(n557), .CI(n574), .S(n1679) );
  XNOR2_X1 U1457 ( .A(n1767), .B(n1663), .ZN(n1680) );
  XOR2_X1 U1458 ( .A(n686), .B(n673), .Z(n1681) );
  XOR2_X1 U1459 ( .A(n671), .B(n1681), .Z(n669) );
  NAND2_X1 U1460 ( .A1(n671), .A2(n686), .ZN(n1682) );
  NAND2_X1 U1461 ( .A1(n671), .A2(n673), .ZN(n1683) );
  NAND2_X1 U1462 ( .A1(n686), .A2(n673), .ZN(n1684) );
  NAND3_X1 U1463 ( .A1(n1682), .A2(n1683), .A3(n1684), .ZN(n668) );
  XOR2_X1 U1464 ( .A(n664), .B(n662), .Z(n1685) );
  XOR2_X1 U1465 ( .A(n660), .B(n1685), .Z(n641) );
  NAND2_X1 U1466 ( .A1(n660), .A2(n664), .ZN(n1686) );
  NAND2_X1 U1467 ( .A1(n660), .A2(n662), .ZN(n1687) );
  NAND2_X1 U1468 ( .A1(n664), .A2(n662), .ZN(n1688) );
  NAND3_X1 U1469 ( .A1(n1686), .A2(n1687), .A3(n1688), .ZN(n640) );
  XNOR2_X1 U1470 ( .A(n615), .B(n1689), .ZN(n613) );
  XNOR2_X1 U1471 ( .A(n634), .B(n617), .ZN(n1689) );
  BUF_X1 U1472 ( .A(n18), .Z(n1909) );
  OR2_X1 U1473 ( .A1(n593), .A2(n612), .ZN(n1837) );
  BUF_X1 U1474 ( .A(a[14]), .Z(n1690) );
  BUF_X1 U1475 ( .A(n71), .Z(n1864) );
  CLKBUF_X1 U1476 ( .A(n1837), .Z(n1708) );
  XOR2_X1 U1477 ( .A(n12), .B(a[2]), .Z(n1465) );
  OR2_X1 U1478 ( .A1(n1811), .A2(n1812), .ZN(n1738) );
  XNOR2_X1 U1479 ( .A(n1870), .B(a[24]), .ZN(n100) );
  BUF_X1 U1480 ( .A(n44), .Z(n1892) );
  BUF_X2 U1481 ( .A(n1935), .Z(n1861) );
  BUF_X2 U1482 ( .A(n27), .Z(n1904) );
  BUF_X2 U1483 ( .A(n116), .Z(n1916) );
  INV_X1 U1484 ( .A(n1701), .ZN(n238) );
  OR2_X1 U1485 ( .A1(n613), .A2(n632), .ZN(n1788) );
  INV_X1 U1486 ( .A(n1788), .ZN(n225) );
  XNOR2_X1 U1487 ( .A(n1600), .B(n1691), .ZN(product[21]) );
  AND2_X1 U1488 ( .A1(n1788), .A2(n226), .ZN(n1691) );
  XNOR2_X1 U1489 ( .A(n180), .B(n1692), .ZN(product[27]) );
  AND2_X1 U1490 ( .A1(n1779), .A2(n1620), .ZN(n1692) );
  BUF_X2 U1491 ( .A(n53), .Z(n1693) );
  INV_X1 U1492 ( .A(n1806), .ZN(n1694) );
  INV_X1 U1493 ( .A(n1806), .ZN(n1695) );
  XNOR2_X1 U1494 ( .A(n173), .B(n1696), .ZN(product[28]) );
  AND2_X1 U1495 ( .A1(n1836), .A2(n172), .ZN(n1696) );
  CLKBUF_X1 U1496 ( .A(n701), .Z(n1697) );
  AND2_X1 U1497 ( .A1(n715), .A2(n728), .ZN(n1698) );
  INV_X1 U1498 ( .A(n1911), .ZN(n1699) );
  CLKBUF_X3 U1499 ( .A(n15), .Z(n1753) );
  BUF_X2 U1500 ( .A(n1724), .Z(n1907) );
  BUF_X2 U1501 ( .A(n63), .Z(n1777) );
  BUF_X2 U1502 ( .A(n63), .Z(n1776) );
  BUF_X2 U1503 ( .A(n1446), .Z(n1756) );
  CLKBUF_X3 U1504 ( .A(n9), .Z(n1912) );
  CLKBUF_X1 U1505 ( .A(n1834), .Z(n1700) );
  OR2_X1 U1506 ( .A1(n571), .A2(n592), .ZN(n1834) );
  AND2_X1 U1507 ( .A1(n633), .A2(n650), .ZN(n1701) );
  XNOR2_X1 U1508 ( .A(n1863), .B(a[18]), .ZN(n1702) );
  BUF_X1 U1509 ( .A(n105), .Z(n1703) );
  BUF_X1 U1510 ( .A(n105), .Z(n1704) );
  BUF_X1 U1511 ( .A(n105), .Z(n1705) );
  XNOR2_X1 U1512 ( .A(n99), .B(a[26]), .ZN(n105) );
  CLKBUF_X1 U1513 ( .A(a[10]), .Z(n1707) );
  OR2_X2 U1514 ( .A1(n1735), .A2(n1734), .ZN(n1709) );
  OR2_X2 U1515 ( .A1(n1735), .A2(n1734), .ZN(n1710) );
  OR2_X1 U1516 ( .A1(n1734), .A2(n1735), .ZN(n77) );
  BUF_X2 U1517 ( .A(n89), .Z(n1711) );
  BUF_X1 U1518 ( .A(n89), .Z(n1865) );
  INV_X1 U1519 ( .A(n261), .ZN(n1712) );
  INV_X1 U1520 ( .A(n1921), .ZN(n1713) );
  INV_X1 U1521 ( .A(n79), .ZN(n1714) );
  INV_X1 U1522 ( .A(n1714), .ZN(n1715) );
  NOR2_X1 U1523 ( .A1(n449), .A2(n474), .ZN(n1716) );
  BUF_X1 U1524 ( .A(n1932), .Z(n1718) );
  XOR2_X1 U1525 ( .A(n1482), .B(n1442), .Z(n1184) );
  BUF_X2 U1526 ( .A(n1876), .Z(n1720) );
  XNOR2_X1 U1527 ( .A(n1857), .B(n1690), .ZN(n1876) );
  OR2_X1 U1528 ( .A1(n1847), .A2(n1848), .ZN(n97) );
  OR2_X1 U1529 ( .A1(n701), .A2(n714), .ZN(n1723) );
  OR2_X1 U1530 ( .A1(n701), .A2(n714), .ZN(n1882) );
  NAND2_X1 U1531 ( .A1(n1465), .A2(n15), .ZN(n1724) );
  BUF_X2 U1532 ( .A(n1601), .Z(n1868) );
  INV_X1 U1533 ( .A(n1591), .ZN(n1725) );
  XNOR2_X1 U1534 ( .A(n30), .B(a[8]), .ZN(n1726) );
  INV_X1 U1535 ( .A(n1901), .ZN(n1728) );
  INV_X1 U1536 ( .A(n1901), .ZN(n1729) );
  INV_X1 U1537 ( .A(n1901), .ZN(n1900) );
  OR2_X2 U1538 ( .A1(n1816), .A2(n1815), .ZN(n84) );
  CLKBUF_X1 U1539 ( .A(n279), .Z(n1732) );
  XNOR2_X1 U1540 ( .A(n1862), .B(a[16]), .ZN(n1734) );
  XOR2_X1 U1541 ( .A(n63), .B(a[16]), .Z(n1735) );
  INV_X1 U1542 ( .A(n1931), .ZN(n1736) );
  INV_X1 U1543 ( .A(n1931), .ZN(n1737) );
  INV_X1 U1544 ( .A(n1931), .ZN(n1928) );
  OR2_X1 U1545 ( .A1(n1811), .A2(n1812), .ZN(n1814) );
  XNOR2_X2 U1546 ( .A(n1870), .B(a[24]), .ZN(n1739) );
  BUF_X2 U1547 ( .A(n99), .Z(n1866) );
  OR2_X1 U1548 ( .A1(n187), .A2(n192), .ZN(n1740) );
  CLKBUF_X1 U1549 ( .A(n241), .Z(n1741) );
  XOR2_X1 U1550 ( .A(n1917), .B(n1482), .Z(n1192) );
  INV_X1 U1551 ( .A(n1779), .ZN(n1742) );
  CLKBUF_X3 U1552 ( .A(n86), .Z(n1743) );
  CLKBUF_X1 U1553 ( .A(n86), .Z(n1856) );
  BUF_X2 U1554 ( .A(n24), .Z(n1744) );
  INV_X1 U1555 ( .A(n1926), .ZN(n1745) );
  INV_X1 U1556 ( .A(n1926), .ZN(n1746) );
  INV_X1 U1557 ( .A(n1926), .ZN(n1925) );
  INV_X1 U1558 ( .A(n50), .ZN(n1747) );
  INV_X2 U1559 ( .A(n1920), .ZN(n1748) );
  INV_X1 U1560 ( .A(n1919), .ZN(n1749) );
  INV_X2 U1561 ( .A(n1927), .ZN(n1750) );
  INV_X2 U1562 ( .A(n1927), .ZN(n1751) );
  CLKBUF_X1 U1563 ( .A(n55), .Z(n1857) );
  XNOR2_X1 U1564 ( .A(n1859), .B(n1690), .ZN(n1875) );
  AND2_X1 U1565 ( .A1(n701), .A2(n714), .ZN(n1752) );
  XNOR2_X1 U1566 ( .A(n104), .B(a[28]), .ZN(n1754) );
  NOR2_X1 U1567 ( .A1(n1730), .A2(n247), .ZN(n1755) );
  INV_X1 U1568 ( .A(n1924), .ZN(n1757) );
  INV_X1 U1569 ( .A(n1924), .ZN(n1922) );
  INV_X1 U1570 ( .A(n184), .ZN(n1759) );
  XNOR2_X1 U1571 ( .A(n626), .B(n1760), .ZN(n603) );
  XNOR2_X1 U1572 ( .A(n628), .B(n630), .ZN(n1760) );
  INV_X1 U1573 ( .A(n1740), .ZN(n1761) );
  NOR2_X1 U1574 ( .A1(n192), .A2(n187), .ZN(n181) );
  INV_X1 U1575 ( .A(n48), .ZN(n1762) );
  INV_X1 U1576 ( .A(n48), .ZN(n1938) );
  XOR2_X1 U1577 ( .A(n1856), .B(a[20]), .Z(n1763) );
  XNOR2_X1 U1578 ( .A(n1863), .B(n1666), .ZN(n1764) );
  XNOR2_X1 U1579 ( .A(n1863), .B(n1666), .ZN(n1873) );
  OR2_X1 U1580 ( .A1(n501), .A2(n524), .ZN(n1765) );
  CLKBUF_X1 U1581 ( .A(n232), .Z(n1766) );
  XNOR2_X1 U1582 ( .A(n1767), .B(n451), .ZN(n449) );
  XNOR2_X1 U1583 ( .A(n476), .B(n453), .ZN(n1767) );
  OR2_X1 U1584 ( .A1(n715), .A2(n728), .ZN(n1768) );
  BUF_X2 U1585 ( .A(n18), .Z(n1769) );
  XNOR2_X1 U1586 ( .A(n1592), .B(n1443), .ZN(n1770) );
  INV_X1 U1587 ( .A(n1920), .ZN(n1771) );
  INV_X1 U1588 ( .A(n1919), .ZN(n1772) );
  NAND2_X1 U1589 ( .A1(n615), .A2(n634), .ZN(n1773) );
  NAND2_X1 U1590 ( .A1(n615), .A2(n617), .ZN(n1774) );
  NAND2_X1 U1591 ( .A1(n634), .A2(n617), .ZN(n1775) );
  NAND3_X1 U1592 ( .A1(n1773), .A2(n1774), .A3(n1775), .ZN(n612) );
  NAND2_X1 U1593 ( .A1(n1595), .A2(n100), .ZN(n1778) );
  OR2_X1 U1594 ( .A1(n500), .A2(n1607), .ZN(n1779) );
  NAND2_X1 U1595 ( .A1(n1454), .A2(n100), .ZN(n102) );
  XNOR2_X1 U1596 ( .A(n12), .B(a[4]), .ZN(n24) );
  CLKBUF_X1 U1597 ( .A(n79), .Z(n1780) );
  NAND2_X1 U1598 ( .A1(n626), .A2(n628), .ZN(n1781) );
  NAND2_X1 U1599 ( .A1(n626), .A2(n630), .ZN(n1782) );
  NAND2_X1 U1600 ( .A1(n628), .A2(n630), .ZN(n1783) );
  NAND3_X1 U1601 ( .A1(n1781), .A2(n1782), .A3(n1783), .ZN(n602) );
  CLKBUF_X1 U1602 ( .A(n79), .Z(n1784) );
  INV_X1 U1603 ( .A(n1901), .ZN(n1785) );
  XNOR2_X1 U1604 ( .A(n21), .B(a[6]), .ZN(n33) );
  BUF_X1 U1605 ( .A(n71), .Z(n1862) );
  XNOR2_X1 U1606 ( .A(n1762), .B(n1707), .ZN(n1461) );
  INV_X1 U1607 ( .A(n1924), .ZN(n1786) );
  NOR2_X1 U1608 ( .A1(n501), .A2(n524), .ZN(n187) );
  NAND2_X1 U1609 ( .A1(n1456), .A2(n1823), .ZN(n91) );
  NAND2_X1 U1610 ( .A1(n99), .A2(n1789), .ZN(n1790) );
  NAND2_X1 U1611 ( .A1(n819), .A2(a[24]), .ZN(n1791) );
  NAND2_X1 U1612 ( .A1(n1790), .A2(n1791), .ZN(n1454) );
  INV_X1 U1613 ( .A(a[24]), .ZN(n1789) );
  INV_X1 U1614 ( .A(n1930), .ZN(n1792) );
  BUF_X2 U1615 ( .A(n61), .Z(n1854) );
  XNOR2_X1 U1616 ( .A(n1793), .B(n976), .ZN(n539) );
  XNOR2_X1 U1617 ( .A(n1022), .B(n1076), .ZN(n1793) );
  BUF_X1 U1618 ( .A(n93), .Z(n1870) );
  XOR2_X1 U1619 ( .A(n1058), .B(n1032), .Z(n1794) );
  XOR2_X1 U1620 ( .A(n1731), .B(n1794), .Z(n723) );
  NAND2_X1 U1621 ( .A1(n1610), .A2(n1032), .ZN(n1795) );
  NAND2_X1 U1622 ( .A1(n986), .A2(n1058), .ZN(n1796) );
  NAND2_X1 U1623 ( .A1(n1032), .A2(n1058), .ZN(n1797) );
  NAND3_X1 U1624 ( .A1(n1795), .A2(n1796), .A3(n1797), .ZN(n722) );
  XNOR2_X1 U1625 ( .A(n1861), .B(n1446), .ZN(n1798) );
  CLKBUF_X1 U1626 ( .A(n79), .Z(n1799) );
  INV_X1 U1627 ( .A(n1901), .ZN(n1899) );
  NAND2_X1 U1628 ( .A1(n976), .A2(n1022), .ZN(n1800) );
  NAND2_X1 U1629 ( .A1(n976), .A2(n1076), .ZN(n1801) );
  NAND2_X1 U1630 ( .A1(n1022), .A2(n1076), .ZN(n1802) );
  NAND3_X1 U1631 ( .A1(n1800), .A2(n1801), .A3(n1802), .ZN(n538) );
  INV_X1 U1632 ( .A(n1890), .ZN(n1888) );
  INV_X4 U1633 ( .A(n1747), .ZN(n1889) );
  XNOR2_X1 U1634 ( .A(n551), .B(n1803), .ZN(n549) );
  XNOR2_X1 U1635 ( .A(n572), .B(n553), .ZN(n1803) );
  INV_X1 U1636 ( .A(n1762), .ZN(n1936) );
  NOR2_X1 U1637 ( .A1(n1716), .A2(n176), .ZN(n1804) );
  CLKBUF_X1 U1638 ( .A(n250), .Z(n1805) );
  XNOR2_X1 U1639 ( .A(n1934), .B(a[8]), .ZN(n1462) );
  XNOR2_X1 U1640 ( .A(n1633), .B(n1762), .ZN(n1806) );
  AND2_X1 U1641 ( .A1(n669), .A2(n684), .ZN(n1807) );
  NAND2_X1 U1642 ( .A1(n1663), .A2(n476), .ZN(n1808) );
  NAND2_X1 U1643 ( .A1(n451), .A2(n453), .ZN(n1809) );
  NAND2_X1 U1644 ( .A1(n476), .A2(n453), .ZN(n1810) );
  NAND3_X1 U1645 ( .A1(n1808), .A2(n1809), .A3(n1810), .ZN(n448) );
  XNOR2_X1 U1646 ( .A(n63), .B(a[14]), .ZN(n1811) );
  XOR2_X1 U1647 ( .A(n55), .B(a[14]), .Z(n1812) );
  OR2_X2 U1648 ( .A1(n1811), .A2(n1812), .ZN(n1813) );
  XNOR2_X1 U1649 ( .A(n79), .B(a[18]), .ZN(n1815) );
  XOR2_X1 U1650 ( .A(n1862), .B(a[18]), .Z(n1816) );
  OR2_X2 U1651 ( .A1(n1816), .A2(n1815), .ZN(n1817) );
  NOR2_X1 U1652 ( .A1(n651), .A2(n668), .ZN(n1818) );
  INV_X1 U1653 ( .A(n1823), .ZN(n1819) );
  NAND2_X1 U1654 ( .A1(n1679), .A2(n572), .ZN(n1820) );
  NAND2_X1 U1655 ( .A1(n1679), .A2(n553), .ZN(n1821) );
  NAND2_X1 U1656 ( .A1(n572), .A2(n553), .ZN(n1822) );
  NAND3_X1 U1657 ( .A1(n1820), .A2(n1821), .A3(n1822), .ZN(n548) );
  XOR2_X1 U1658 ( .A(n1938), .B(a[12]), .Z(n58) );
  XNOR2_X1 U1659 ( .A(n79), .B(a[20]), .ZN(n1823) );
  OR2_X1 U1660 ( .A1(n421), .A2(n448), .ZN(n1831) );
  CLKBUF_X1 U1661 ( .A(n6), .Z(n1914) );
  BUF_X4 U1662 ( .A(n74), .Z(n1869) );
  BUF_X2 U1663 ( .A(n36), .Z(n1897) );
  XNOR2_X1 U1664 ( .A(n86), .B(a[22]), .ZN(n95) );
  XNOR2_X1 U1665 ( .A(n194), .B(n1824), .ZN(product[25]) );
  NAND2_X1 U1666 ( .A1(n338), .A2(n193), .ZN(n1824) );
  XOR2_X1 U1667 ( .A(n255), .B(n1825), .Z(product[17]) );
  AND2_X1 U1668 ( .A1(n346), .A2(n254), .ZN(n1825) );
  AND2_X1 U1669 ( .A1(n1845), .A2(n331), .ZN(product[1]) );
  AOI21_X1 U1670 ( .B1(n1708), .B2(n228), .A(n1615), .ZN(n1827) );
  BUF_X1 U1671 ( .A(n6), .Z(n1828) );
  BUF_X1 U1672 ( .A(n6), .Z(n1829) );
  OAI21_X1 U1673 ( .B1(n193), .B2(n187), .A(n188), .ZN(n182) );
  INV_X1 U1674 ( .A(n214), .ZN(n216) );
  INV_X1 U1675 ( .A(n165), .ZN(n163) );
  INV_X1 U1676 ( .A(n193), .ZN(n191) );
  AND2_X1 U1677 ( .A1(n1835), .A2(n1831), .ZN(n1830) );
  INV_X1 U1678 ( .A(n156), .ZN(n154) );
  INV_X1 U1679 ( .A(n160), .ZN(n158) );
  NAND2_X1 U1680 ( .A1(n525), .A2(n548), .ZN(n193) );
  AOI21_X1 U1681 ( .B1(n249), .B2(n1880), .A(n1807), .ZN(n244) );
  OR2_X1 U1682 ( .A1(n549), .A2(n570), .ZN(n1832) );
  NAND2_X1 U1683 ( .A1(n1607), .A2(n500), .ZN(n179) );
  NAND2_X1 U1684 ( .A1(n501), .A2(n524), .ZN(n188) );
  NAND2_X1 U1685 ( .A1(n421), .A2(n448), .ZN(n165) );
  NAND2_X1 U1686 ( .A1(n393), .A2(n420), .ZN(n160) );
  INV_X1 U1687 ( .A(n253), .ZN(n346) );
  OR2_X1 U1688 ( .A1(n393), .A2(n420), .ZN(n1835) );
  OR2_X1 U1689 ( .A1(n1594), .A2(n474), .ZN(n1836) );
  INV_X1 U1690 ( .A(n1698), .ZN(n264) );
  INV_X1 U1691 ( .A(n1881), .ZN(n223) );
  INV_X1 U1692 ( .A(n304), .ZN(n302) );
  AOI21_X1 U1693 ( .B1(n287), .B2(n351), .A(n284), .ZN(n282) );
  INV_X1 U1694 ( .A(n286), .ZN(n284) );
  NOR2_X1 U1695 ( .A1(n685), .A2(n700), .ZN(n253) );
  INV_X1 U1696 ( .A(n285), .ZN(n351) );
  NOR2_X1 U1697 ( .A1(n280), .A2(n285), .ZN(n278) );
  OAI21_X1 U1698 ( .B1(n296), .B2(n294), .A(n295), .ZN(n293) );
  OR2_X2 U1699 ( .A1(n729), .A2(n740), .ZN(n1838) );
  NAND2_X1 U1700 ( .A1(n685), .A2(n700), .ZN(n254) );
  NAND2_X1 U1701 ( .A1(n729), .A2(n740), .ZN(n276) );
  INV_X1 U1702 ( .A(n294), .ZN(n353) );
  INV_X1 U1703 ( .A(n298), .ZN(n354) );
  INV_X1 U1704 ( .A(n320), .ZN(n318) );
  OAI21_X1 U1705 ( .B1(n322), .B2(n324), .A(n323), .ZN(n321) );
  NAND2_X1 U1706 ( .A1(n773), .A2(n780), .ZN(n295) );
  AOI21_X1 U1707 ( .B1(n1843), .B2(n329), .A(n326), .ZN(n324) );
  INV_X1 U1708 ( .A(n328), .ZN(n326) );
  NOR2_X1 U1709 ( .A1(n763), .A2(n772), .ZN(n291) );
  NOR2_X1 U1710 ( .A1(n773), .A2(n780), .ZN(n294) );
  INV_X1 U1711 ( .A(n331), .ZN(n329) );
  NOR2_X1 U1712 ( .A1(n781), .A2(n788), .ZN(n298) );
  NAND2_X1 U1713 ( .A1(n781), .A2(n788), .ZN(n299) );
  NAND2_X1 U1714 ( .A1(n789), .A2(n794), .ZN(n304) );
  NAND2_X1 U1715 ( .A1(n763), .A2(n772), .ZN(n292) );
  OR2_X1 U1716 ( .A1(n789), .A2(n794), .ZN(n1839) );
  NAND2_X1 U1717 ( .A1(n741), .A2(n752), .ZN(n281) );
  INV_X1 U1718 ( .A(n314), .ZN(n358) );
  INV_X1 U1719 ( .A(n306), .ZN(n356) );
  INV_X1 U1720 ( .A(n322), .ZN(n360) );
  OR2_X1 U1721 ( .A1(n364), .A2(n392), .ZN(n1840) );
  XNOR2_X1 U1722 ( .A(n1841), .B(n363), .ZN(n364) );
  XNOR2_X1 U1723 ( .A(n365), .B(n400), .ZN(n1841) );
  OR2_X1 U1724 ( .A1(n801), .A2(n804), .ZN(n1842) );
  OR2_X1 U1725 ( .A1(n1129), .A2(n1099), .ZN(n1843) );
  NOR2_X1 U1726 ( .A1(n795), .A2(n800), .ZN(n306) );
  NAND2_X1 U1727 ( .A1(n795), .A2(n800), .ZN(n307) );
  OR2_X1 U1728 ( .A1(n809), .A2(n810), .ZN(n1844) );
  NAND2_X1 U1729 ( .A1(n801), .A2(n804), .ZN(n312) );
  NAND2_X1 U1730 ( .A1(n809), .A2(n810), .ZN(n320) );
  OR2_X1 U1731 ( .A1(n1130), .A2(n859), .ZN(n1845) );
  AND2_X1 U1732 ( .A1(n1916), .A2(n816), .ZN(n871) );
  AND2_X1 U1733 ( .A1(n1915), .A2(n1634), .ZN(n991) );
  AND2_X1 U1734 ( .A1(n1915), .A2(n814), .ZN(n865) );
  OAI22_X1 U1735 ( .A1(n1896), .A2(n1312), .B1(n1900), .B2(n1311), .ZN(n1028)
         );
  AND2_X1 U1736 ( .A1(n1915), .A2(n1644), .ZN(n969) );
  OAI22_X1 U1737 ( .A1(n1903), .A2(n1343), .B1(n1744), .B2(n1342), .ZN(n1058)
         );
  OAI22_X1 U1738 ( .A1(n1913), .A2(n1400), .B1(n1399), .B2(n1914), .ZN(n1113)
         );
  OR2_X1 U1739 ( .A1(n1915), .A2(n1920), .ZN(n1418) );
  XNOR2_X1 U1740 ( .A(n1917), .B(n1871), .ZN(n1164) );
  OR2_X1 U1741 ( .A1(n1916), .A2(n1725), .ZN(n1298) );
  OAI22_X1 U1742 ( .A1(n1912), .A2(n1417), .B1(n1416), .B2(n1828), .ZN(n1130)
         );
  OR2_X1 U1743 ( .A1(n1915), .A2(n817), .ZN(n1145) );
  AND2_X1 U1744 ( .A1(n1915), .A2(n1895), .ZN(n1015) );
  OAI22_X1 U1745 ( .A1(n1902), .A2(n1350), .B1(n1744), .B2(n1349), .ZN(n1065)
         );
  OAI22_X1 U1746 ( .A1(n1898), .A2(n1323), .B1(n1729), .B2(n1322), .ZN(n1039)
         );
  OAI22_X1 U1747 ( .A1(n1902), .A2(n1353), .B1(n1744), .B2(n1352), .ZN(n1068)
         );
  OR2_X1 U1748 ( .A1(n1916), .A2(n1927), .ZN(n1354) );
  OR2_X1 U1749 ( .A1(n1916), .A2(n1483), .ZN(n1210) );
  XOR2_X1 U1750 ( .A(n862), .B(n844), .Z(n391) );
  OAI22_X1 U1751 ( .A1(n115), .A2(n813), .B1(n1133), .B2(n114), .ZN(n844) );
  OAI22_X1 U1752 ( .A1(n1628), .A2(n1135), .B1(n1134), .B2(n1754), .ZN(n862)
         );
  XNOR2_X1 U1753 ( .A(n408), .B(n1846), .ZN(n371) );
  XNOR2_X1 U1754 ( .A(n384), .B(n375), .ZN(n1846) );
  BUF_X2 U1755 ( .A(n27), .Z(n1903) );
  AND2_X1 U1756 ( .A1(n1916), .A2(n1906), .ZN(n1069) );
  BUF_X2 U1757 ( .A(n44), .Z(n1891) );
  OAI22_X1 U1758 ( .A1(n115), .A2(n1132), .B1(n1131), .B2(n114), .ZN(n860) );
  OAI22_X1 U1759 ( .A1(n1717), .A2(n1399), .B1(n1398), .B2(n1828), .ZN(n1112)
         );
  OAI22_X1 U1760 ( .A1(n1913), .A2(n1398), .B1(n1397), .B2(n1914), .ZN(n1111)
         );
  AND2_X1 U1761 ( .A1(n1916), .A2(n1590), .ZN(n889) );
  AND2_X1 U1762 ( .A1(n1916), .A2(n824), .ZN(n915) );
  OAI22_X1 U1763 ( .A1(n1902), .A2(n1341), .B1(n1744), .B2(n1340), .ZN(n1056)
         );
  OAI22_X1 U1764 ( .A1(n1912), .A2(n1401), .B1(n1400), .B2(n1829), .ZN(n1114)
         );
  OAI22_X1 U1765 ( .A1(n1902), .A2(n1336), .B1(n1905), .B2(n1335), .ZN(n1051)
         );
  OAI22_X1 U1766 ( .A1(n1769), .A2(n1365), .B1(n1753), .B2(n1364), .ZN(n1079)
         );
  AND2_X1 U1767 ( .A1(n1916), .A2(n812), .ZN(n861) );
  OAI22_X1 U1768 ( .A1(n112), .A2(n1136), .B1(n1135), .B2(n1754), .ZN(n863) );
  OAI22_X1 U1769 ( .A1(n1902), .A2(n1335), .B1(n1905), .B2(n1334), .ZN(n1050)
         );
  OAI22_X1 U1770 ( .A1(n1717), .A2(n1405), .B1(n1404), .B2(n1829), .ZN(n1118)
         );
  OAI22_X1 U1771 ( .A1(n1904), .A2(n1334), .B1(n1905), .B2(n1333), .ZN(n1049)
         );
  OAI22_X1 U1772 ( .A1(n1896), .A2(n1307), .B1(n1729), .B2(n1306), .ZN(n1023)
         );
  OAI22_X1 U1773 ( .A1(n1903), .A2(n1342), .B1(n1744), .B2(n1341), .ZN(n1057)
         );
  OAI22_X1 U1774 ( .A1(n1902), .A2(n1348), .B1(n1744), .B2(n1347), .ZN(n1063)
         );
  OAI22_X1 U1775 ( .A1(n1912), .A2(n1408), .B1(n1407), .B2(n1828), .ZN(n1121)
         );
  OAI22_X1 U1776 ( .A1(n1896), .A2(n1322), .B1(n1785), .B2(n1321), .ZN(n1038)
         );
  OAI22_X1 U1777 ( .A1(n1902), .A2(n1344), .B1(n1744), .B2(n1343), .ZN(n1059)
         );
  OAI22_X1 U1778 ( .A1(n1898), .A2(n1305), .B1(n1728), .B2(n1304), .ZN(n1021)
         );
  OAI22_X1 U1779 ( .A1(n1904), .A2(n1351), .B1(n1744), .B2(n1350), .ZN(n1066)
         );
  OAI22_X1 U1780 ( .A1(n1902), .A2(n1349), .B1(n1744), .B2(n1348), .ZN(n1064)
         );
  AND2_X1 U1781 ( .A1(n1916), .A2(n1901), .ZN(n1041) );
  OAI22_X1 U1782 ( .A1(n1896), .A2(n1308), .B1(n1728), .B2(n1307), .ZN(n1024)
         );
  AND2_X1 U1783 ( .A1(n1915), .A2(n818), .ZN(n879) );
  OAI22_X1 U1784 ( .A1(n1897), .A2(n1310), .B1(n1899), .B2(n1309), .ZN(n1026)
         );
  OAI22_X1 U1785 ( .A1(n1909), .A2(n1367), .B1(n1910), .B2(n1366), .ZN(n1081)
         );
  OAI22_X1 U1786 ( .A1(n1897), .A2(n1311), .B1(n1728), .B2(n1310), .ZN(n1027)
         );
  OAI22_X1 U1787 ( .A1(n1904), .A2(n1339), .B1(n1905), .B2(n1338), .ZN(n1054)
         );
  OAI22_X1 U1788 ( .A1(n1908), .A2(n1368), .B1(n1678), .B2(n1367), .ZN(n1082)
         );
  OAI22_X1 U1789 ( .A1(n1896), .A2(n1306), .B1(n1785), .B2(n1305), .ZN(n1022)
         );
  OAI22_X1 U1790 ( .A1(n1912), .A2(n1404), .B1(n1403), .B2(n1828), .ZN(n1117)
         );
  AND2_X1 U1791 ( .A1(n1915), .A2(n1735), .ZN(n931) );
  XNOR2_X1 U1792 ( .A(n1917), .B(n1866), .ZN(n1153) );
  XNOR2_X1 U1793 ( .A(n1915), .B(n1864), .ZN(n1209) );
  OAI22_X1 U1794 ( .A1(n1898), .A2(n1309), .B1(n1785), .B2(n1308), .ZN(n1025)
         );
  OAI22_X1 U1795 ( .A1(n1902), .A2(n1332), .B1(n1744), .B2(n1331), .ZN(n1047)
         );
  OAI22_X1 U1796 ( .A1(n1913), .A2(n1403), .B1(n1402), .B2(n1829), .ZN(n1116)
         );
  OAI22_X1 U1797 ( .A1(n1913), .A2(n1402), .B1(n1401), .B2(n1829), .ZN(n1115)
         );
  OAI22_X1 U1798 ( .A1(n1904), .A2(n1340), .B1(n1744), .B2(n1339), .ZN(n1055)
         );
  OAI22_X1 U1799 ( .A1(n1896), .A2(n1313), .B1(n1900), .B2(n1312), .ZN(n1029)
         );
  OAI22_X1 U1800 ( .A1(n1912), .A2(n1407), .B1(n1406), .B2(n1829), .ZN(n1120)
         );
  OAI22_X1 U1801 ( .A1(n1912), .A2(n1406), .B1(n1405), .B2(n1914), .ZN(n1119)
         );
  INV_X1 U1802 ( .A(n1754), .ZN(n814) );
  OR2_X1 U1803 ( .A1(n1915), .A2(n1482), .ZN(n1193) );
  OR2_X1 U1804 ( .A1(n1917), .A2(n819), .ZN(n1154) );
  OAI22_X1 U1805 ( .A1(n1896), .A2(n1324), .B1(n1785), .B2(n1323), .ZN(n1040)
         );
  OR2_X1 U1806 ( .A1(n1916), .A2(n1931), .ZN(n1325) );
  INV_X1 U1807 ( .A(n114), .ZN(n812) );
  INV_X1 U1808 ( .A(n1871), .ZN(n1480) );
  AND2_X1 U1809 ( .A1(n1916), .A2(n1911), .ZN(n1099) );
  INV_X1 U1810 ( .A(n99), .ZN(n819) );
  INV_X1 U1811 ( .A(n1863), .ZN(n1483) );
  OR2_X1 U1812 ( .A1(n1916), .A2(n815), .ZN(n1138) );
  OR2_X1 U1813 ( .A1(n1915), .A2(n813), .ZN(n1133) );
  CLKBUF_X1 U1814 ( .A(n36), .Z(n1898) );
  OR2_X1 U1815 ( .A1(n1916), .A2(n1484), .ZN(n1229) );
  OR2_X1 U1816 ( .A1(n1917), .A2(n1480), .ZN(n1165) );
  OR2_X1 U1817 ( .A1(n1916), .A2(n1481), .ZN(n1178) );
  XNOR2_X1 U1818 ( .A(n104), .B(a[28]), .ZN(n110) );
  XNOR2_X1 U1819 ( .A(n109), .B(a[30]), .ZN(n114) );
  XNOR2_X1 U1820 ( .A(n1603), .B(n109), .ZN(n1136) );
  CLKBUF_X3 U1821 ( .A(n93), .Z(n1871) );
  XNOR2_X1 U1822 ( .A(n1448), .B(n109), .ZN(n1135) );
  XNOR2_X1 U1823 ( .A(n1863), .B(n1603), .ZN(n1208) );
  XNOR2_X1 U1824 ( .A(n1863), .B(n1445), .ZN(n1204) );
  XNOR2_X1 U1825 ( .A(n1861), .B(n1445), .ZN(n1267) );
  XNOR2_X1 U1826 ( .A(n1871), .B(n1445), .ZN(n1159) );
  XNOR2_X1 U1827 ( .A(n1596), .B(n1445), .ZN(n1379) );
  XNOR2_X1 U1828 ( .A(n1602), .B(n1871), .ZN(n1163) );
  XNOR2_X1 U1829 ( .A(n1866), .B(n1445), .ZN(n1148) );
  XNOR2_X1 U1830 ( .A(n1772), .B(n1445), .ZN(n1412) );
  XNOR2_X1 U1831 ( .A(n1737), .B(n1443), .ZN(n1317) );
  XNOR2_X1 U1832 ( .A(n1864), .B(n1443), .ZN(n1202) );
  XNOR2_X1 U1833 ( .A(n1757), .B(n1443), .ZN(n1377) );
  XNOR2_X1 U1834 ( .A(n1871), .B(n1443), .ZN(n1157) );
  XNOR2_X1 U1835 ( .A(n1861), .B(n1443), .ZN(n1265) );
  XNOR2_X1 U1836 ( .A(n1602), .B(n1866), .ZN(n1152) );
  XNOR2_X1 U1837 ( .A(n1772), .B(n1443), .ZN(n1410) );
  XNOR2_X1 U1838 ( .A(n1864), .B(n1446), .ZN(n1205) );
  XNOR2_X1 U1839 ( .A(n1871), .B(n1446), .ZN(n1160) );
  XNOR2_X1 U1840 ( .A(n1866), .B(n1446), .ZN(n1149) );
  XNOR2_X1 U1841 ( .A(n1921), .B(n1446), .ZN(n1380) );
  XNOR2_X1 U1842 ( .A(n1772), .B(n1446), .ZN(n1413) );
  XNOR2_X1 U1843 ( .A(n1864), .B(n1444), .ZN(n1203) );
  XNOR2_X1 U1844 ( .A(n1871), .B(n1444), .ZN(n1158) );
  XNOR2_X1 U1845 ( .A(n1861), .B(n1444), .ZN(n1266) );
  XNOR2_X1 U1846 ( .A(n1786), .B(n1444), .ZN(n1378) );
  XNOR2_X1 U1847 ( .A(n1444), .B(n1866), .ZN(n1147) );
  XNOR2_X1 U1848 ( .A(n1737), .B(n1437), .ZN(n1311) );
  XNOR2_X1 U1849 ( .A(n1786), .B(n1447), .ZN(n1381) );
  XNOR2_X1 U1850 ( .A(n1748), .B(n1444), .ZN(n1411) );
  XNOR2_X1 U1851 ( .A(n1603), .B(n113), .ZN(n1131) );
  XNOR2_X1 U1852 ( .A(n1918), .B(n1436), .ZN(n1403) );
  XNOR2_X1 U1853 ( .A(n1918), .B(n1435), .ZN(n1402) );
  XNOR2_X1 U1854 ( .A(n1772), .B(n1432), .ZN(n1399) );
  XNOR2_X1 U1855 ( .A(n1748), .B(n1434), .ZN(n1401) );
  XNOR2_X1 U1856 ( .A(n1771), .B(n1433), .ZN(n1400) );
  XNOR2_X1 U1857 ( .A(n1748), .B(n1437), .ZN(n1404) );
  XNOR2_X1 U1858 ( .A(n1749), .B(n1439), .ZN(n1406) );
  XNOR2_X1 U1859 ( .A(n1749), .B(n1438), .ZN(n1405) );
  XNOR2_X1 U1860 ( .A(n1861), .B(n1448), .ZN(n1270) );
  XNOR2_X1 U1861 ( .A(n1871), .B(n1448), .ZN(n1162) );
  XNOR2_X1 U1862 ( .A(n1866), .B(n1448), .ZN(n1151) );
  XNOR2_X1 U1863 ( .A(n1447), .B(n1871), .ZN(n1161) );
  XNOR2_X1 U1864 ( .A(n1736), .B(n1438), .ZN(n1312) );
  XNOR2_X1 U1865 ( .A(n1447), .B(n1866), .ZN(n1150) );
  XNOR2_X1 U1866 ( .A(n1864), .B(n1437), .ZN(n1196) );
  XNOR2_X1 U1867 ( .A(n1864), .B(n1438), .ZN(n1197) );
  XNOR2_X1 U1868 ( .A(n1667), .B(a[22]), .ZN(n1847) );
  INV_X1 U1869 ( .A(n95), .ZN(n1848) );
  CLKBUF_X3 U1870 ( .A(n116), .Z(n1915) );
  XNOR2_X1 U1871 ( .A(n1737), .B(n1435), .ZN(n1309) );
  XNOR2_X1 U1872 ( .A(n1737), .B(n1436), .ZN(n1310) );
  XNOR2_X1 U1873 ( .A(n1792), .B(n1434), .ZN(n1308) );
  XNOR2_X1 U1874 ( .A(n1736), .B(n1431), .ZN(n1305) );
  XNOR2_X1 U1875 ( .A(n1447), .B(n109), .ZN(n1134) );
  XNOR2_X1 U1876 ( .A(n1923), .B(n1433), .ZN(n1367) );
  XNOR2_X1 U1877 ( .A(n1929), .B(n1433), .ZN(n1307) );
  XNOR2_X1 U1878 ( .A(n1746), .B(n1432), .ZN(n1335) );
  XNOR2_X1 U1879 ( .A(n1929), .B(n1432), .ZN(n1306) );
  XNOR2_X1 U1880 ( .A(n1736), .B(n1439), .ZN(n1313) );
  OAI22_X1 U1881 ( .A1(n112), .A2(n1137), .B1(n1136), .B2(n1754), .ZN(n864) );
  OAI22_X1 U1882 ( .A1(n112), .A2(n815), .B1(n1138), .B2(n1754), .ZN(n845) );
  XNOR2_X1 U1883 ( .A(n1917), .B(n109), .ZN(n1137) );
  XNOR2_X1 U1884 ( .A(n1925), .B(n1435), .ZN(n1338) );
  XNOR2_X1 U1885 ( .A(n1736), .B(n1442), .ZN(n1316) );
  XNOR2_X1 U1886 ( .A(n1863), .B(n1442), .ZN(n1201) );
  XNOR2_X1 U1887 ( .A(n1871), .B(n1442), .ZN(n1156) );
  XNOR2_X1 U1888 ( .A(n1928), .B(n1441), .ZN(n1315) );
  XNOR2_X1 U1889 ( .A(n1863), .B(n1441), .ZN(n1200) );
  XNOR2_X1 U1890 ( .A(n1932), .B(n1437), .ZN(n1284) );
  XNOR2_X1 U1891 ( .A(n1923), .B(n1437), .ZN(n1371) );
  XNOR2_X1 U1892 ( .A(n1936), .B(n1437), .ZN(n1259) );
  XNOR2_X1 U1893 ( .A(n1863), .B(n1439), .ZN(n1198) );
  XNOR2_X1 U1894 ( .A(n1718), .B(n1439), .ZN(n1286) );
  XNOR2_X1 U1895 ( .A(n1933), .B(n1438), .ZN(n1285) );
  XNOR2_X1 U1896 ( .A(n1937), .B(n1438), .ZN(n1260) );
  XNOR2_X1 U1897 ( .A(n1918), .B(n1430), .ZN(n1397) );
  XNOR2_X1 U1898 ( .A(n1745), .B(n1433), .ZN(n1336) );
  XNOR2_X1 U1899 ( .A(n1923), .B(n1434), .ZN(n1368) );
  XNOR2_X1 U1900 ( .A(n1866), .B(n1443), .ZN(n1146) );
  XNOR2_X1 U1901 ( .A(n992), .B(n1849), .ZN(n382) );
  XNOR2_X1 U1902 ( .A(n1042), .B(n1016), .ZN(n1849) );
  XNOR2_X1 U1903 ( .A(n1933), .B(n1440), .ZN(n1287) );
  XNOR2_X1 U1904 ( .A(n1928), .B(n1440), .ZN(n1314) );
  XNOR2_X1 U1905 ( .A(n1863), .B(n1440), .ZN(n1199) );
  XNOR2_X1 U1906 ( .A(n1933), .B(n1435), .ZN(n1282) );
  XNOR2_X1 U1907 ( .A(n1757), .B(n1435), .ZN(n1369) );
  XNOR2_X1 U1908 ( .A(n1936), .B(n1435), .ZN(n1257) );
  XNOR2_X1 U1909 ( .A(n1933), .B(n1436), .ZN(n1283) );
  XNOR2_X1 U1910 ( .A(n1923), .B(n1436), .ZN(n1370) );
  XNOR2_X1 U1911 ( .A(n1936), .B(n1436), .ZN(n1258) );
  XNOR2_X1 U1912 ( .A(n152), .B(n1850), .ZN(product[31]) );
  AND2_X1 U1913 ( .A1(n1840), .A2(n151), .ZN(n1850) );
  XNOR2_X1 U1914 ( .A(n161), .B(n1851), .ZN(product[30]) );
  AND2_X1 U1915 ( .A1(n1835), .A2(n160), .ZN(n1851) );
  XNOR2_X1 U1916 ( .A(n1923), .B(n1432), .ZN(n1366) );
  XNOR2_X1 U1917 ( .A(n1596), .B(n1430), .ZN(n1364) );
  XNOR2_X1 U1918 ( .A(n1929), .B(n1430), .ZN(n1304) );
  XNOR2_X1 U1919 ( .A(n1925), .B(n1434), .ZN(n1337) );
  XNOR2_X1 U1920 ( .A(n1933), .B(n1434), .ZN(n1281) );
  XNOR2_X1 U1921 ( .A(n1936), .B(n1433), .ZN(n1255) );
  XNOR2_X1 U1922 ( .A(n1937), .B(n1434), .ZN(n1256) );
  XNOR2_X1 U1923 ( .A(n1933), .B(n1433), .ZN(n1280) );
  XNOR2_X1 U1924 ( .A(n1871), .B(n1441), .ZN(n1155) );
  XNOR2_X1 U1925 ( .A(n1748), .B(n1428), .ZN(n1395) );
  XNOR2_X1 U1926 ( .A(n1772), .B(n1427), .ZN(n1394) );
  XNOR2_X1 U1927 ( .A(n1771), .B(n1429), .ZN(n1396) );
  XNOR2_X1 U1928 ( .A(n1748), .B(b[24]), .ZN(n1393) );
  XNOR2_X1 U1929 ( .A(n1933), .B(n1432), .ZN(n1279) );
  XNOR2_X1 U1930 ( .A(n1936), .B(n1432), .ZN(n1254) );
  XNOR2_X1 U1931 ( .A(n1792), .B(n1429), .ZN(n1303) );
  XNOR2_X1 U1932 ( .A(n1792), .B(n1428), .ZN(n1302) );
  XNOR2_X1 U1933 ( .A(n1861), .B(n1431), .ZN(n1253) );
  XNOR2_X1 U1934 ( .A(n1861), .B(n1430), .ZN(n1252) );
  XNOR2_X1 U1935 ( .A(n1757), .B(n1429), .ZN(n1363) );
  XNOR2_X1 U1936 ( .A(n1745), .B(n1427), .ZN(n1330) );
  XNOR2_X1 U1937 ( .A(n1745), .B(b[24]), .ZN(n1329) );
  XNOR2_X1 U1938 ( .A(n1596), .B(n1428), .ZN(n1362) );
  XNOR2_X1 U1939 ( .A(n1929), .B(n1427), .ZN(n1301) );
  XNOR2_X1 U1940 ( .A(n1929), .B(b[24]), .ZN(n1300) );
  XNOR2_X1 U1941 ( .A(n1916), .B(n113), .ZN(n1132) );
  NAND2_X1 U1942 ( .A1(n356), .A2(n307), .ZN(n143) );
  XNOR2_X1 U1943 ( .A(n189), .B(n1852), .ZN(product[26]) );
  AND2_X1 U1944 ( .A1(n1765), .A2(n188), .ZN(n1852) );
  INV_X1 U1945 ( .A(n109), .ZN(n815) );
  NAND2_X1 U1946 ( .A1(n1452), .A2(n110), .ZN(n112) );
  XOR2_X1 U1947 ( .A(n109), .B(a[28]), .Z(n1452) );
  XOR2_X1 U1948 ( .A(n244), .B(n131), .Z(product[19]) );
  NAND2_X1 U1949 ( .A1(n344), .A2(n243), .ZN(n131) );
  XOR2_X1 U1950 ( .A(n277), .B(n136), .Z(product[14]) );
  NAND2_X1 U1951 ( .A1(n1838), .A2(n276), .ZN(n136) );
  XNOR2_X1 U1952 ( .A(n1922), .B(b[29]), .ZN(n1355) );
  NAND2_X1 U1953 ( .A1(n1451), .A2(n114), .ZN(n115) );
  XOR2_X1 U1954 ( .A(n113), .B(a[30]), .Z(n1451) );
  XNOR2_X1 U1955 ( .A(n148), .B(n329), .ZN(product[2]) );
  NAND2_X1 U1956 ( .A1(n1843), .A2(n328), .ZN(n148) );
  INV_X1 U1957 ( .A(n113), .ZN(n813) );
  INV_X1 U1958 ( .A(n842), .ZN(n6) );
  XNOR2_X1 U1959 ( .A(n213), .B(n127), .ZN(product[23]) );
  XOR2_X1 U1960 ( .A(n204), .B(n1853), .Z(product[24]) );
  AND2_X1 U1961 ( .A1(n1832), .A2(n203), .ZN(n1853) );
  XOR2_X1 U1962 ( .A(n239), .B(n130), .Z(product[20]) );
  XNOR2_X1 U1963 ( .A(n249), .B(n132), .ZN(product[18]) );
  XNOR2_X1 U1964 ( .A(n262), .B(n134), .ZN(product[16]) );
  XOR2_X1 U1965 ( .A(n147), .B(n324), .Z(product[3]) );
  XNOR2_X1 U1966 ( .A(n146), .B(n321), .ZN(product[4]) );
  NAND2_X1 U1967 ( .A1(n1844), .A2(n320), .ZN(n146) );
  NAND2_X1 U1968 ( .A1(n358), .A2(n315), .ZN(n145) );
  NAND2_X1 U1969 ( .A1(n1842), .A2(n312), .ZN(n144) );
  XOR2_X1 U1970 ( .A(n282), .B(n137), .Z(product[13]) );
  NAND2_X1 U1971 ( .A1(n350), .A2(n281), .ZN(n137) );
  XOR2_X1 U1972 ( .A(n269), .B(n135), .Z(product[15]) );
  XNOR2_X1 U1973 ( .A(n293), .B(n139), .ZN(product[11]) );
  NAND2_X1 U1974 ( .A1(n352), .A2(n292), .ZN(n139) );
  XNOR2_X1 U1975 ( .A(n287), .B(n138), .ZN(product[12]) );
  NAND2_X1 U1976 ( .A1(n351), .A2(n1635), .ZN(n138) );
  XOR2_X1 U1977 ( .A(n296), .B(n140), .Z(product[10]) );
  NAND2_X1 U1978 ( .A1(n353), .A2(n295), .ZN(n140) );
  NAND2_X1 U1979 ( .A1(n1839), .A2(n304), .ZN(n142) );
  AND2_X1 U1980 ( .A1(n1916), .A2(n842), .ZN(product[0]) );
  NAND2_X1 U1981 ( .A1(n354), .A2(n299), .ZN(n141) );
  INV_X1 U1982 ( .A(n15), .ZN(n1911) );
  OAI22_X1 U1983 ( .A1(n107), .A2(n1140), .B1(n1704), .B2(n1139), .ZN(n866) );
  OAI22_X1 U1984 ( .A1(n107), .A2(n1142), .B1(n1141), .B2(n1705), .ZN(n868) );
  OAI22_X1 U1985 ( .A1(n107), .A2(n1141), .B1(n1704), .B2(n1140), .ZN(n867) );
  OAI22_X1 U1986 ( .A1(n107), .A2(n1144), .B1(n1143), .B2(n1704), .ZN(n870) );
  OAI22_X1 U1987 ( .A1(n107), .A2(n817), .B1(n1145), .B2(n1705), .ZN(n846) );
  OAI22_X1 U1988 ( .A1(n107), .A2(n1143), .B1(n1705), .B2(n1142), .ZN(n869) );
  INV_X1 U1989 ( .A(n1705), .ZN(n816) );
  AND2_X1 U1990 ( .A1(n1915), .A2(n1819), .ZN(n901) );
  XNOR2_X1 U1991 ( .A(n1750), .B(b[27]), .ZN(n1326) );
  XNOR2_X1 U1992 ( .A(n1751), .B(b[26]), .ZN(n1327) );
  XNOR2_X1 U1993 ( .A(n1751), .B(n1443), .ZN(n1346) );
  XNOR2_X1 U1994 ( .A(n1751), .B(n1444), .ZN(n1347) );
  XNOR2_X1 U1995 ( .A(n1751), .B(n1445), .ZN(n1348) );
  XNOR2_X1 U1996 ( .A(n1750), .B(n1756), .ZN(n1349) );
  XNOR2_X1 U1997 ( .A(n1750), .B(b[25]), .ZN(n1328) );
  XNOR2_X1 U1998 ( .A(n1750), .B(n1447), .ZN(n1350) );
  XNOR2_X1 U1999 ( .A(n1751), .B(n1431), .ZN(n1334) );
  XNOR2_X1 U2000 ( .A(n1751), .B(n1428), .ZN(n1331) );
  XNOR2_X1 U2001 ( .A(n1746), .B(n1430), .ZN(n1333) );
  XNOR2_X1 U2002 ( .A(n1750), .B(n1603), .ZN(n1352) );
  XNOR2_X1 U2003 ( .A(n1745), .B(n1448), .ZN(n1351) );
  XNOR2_X1 U2004 ( .A(n1746), .B(n1429), .ZN(n1332) );
  INV_X1 U2005 ( .A(n192), .ZN(n338) );
  NAND2_X1 U2006 ( .A1(n58), .A2(n1460), .ZN(n61) );
  OAI22_X1 U2007 ( .A1(n1733), .A2(n1297), .B1(n1665), .B2(n1296), .ZN(n1014)
         );
  OAI22_X1 U2008 ( .A1(n1891), .A2(n1286), .B1(n1665), .B2(n1285), .ZN(n1003)
         );
  OAI22_X1 U2009 ( .A1(n1733), .A2(n1278), .B1(n1894), .B2(n1277), .ZN(n995)
         );
  OAI22_X1 U2010 ( .A1(n1891), .A2(n1282), .B1(n1664), .B2(n1281), .ZN(n999)
         );
  OAI22_X1 U2011 ( .A1(n1891), .A2(n1279), .B1(n1278), .B2(n1894), .ZN(n996)
         );
  OAI22_X1 U2012 ( .A1(n1892), .A2(n1280), .B1(n1893), .B2(n1279), .ZN(n997)
         );
  OAI22_X1 U2013 ( .A1(n1891), .A2(n1281), .B1(n1664), .B2(n1280), .ZN(n998)
         );
  BUF_X2 U2014 ( .A(n1724), .Z(n1908) );
  INV_X1 U2015 ( .A(n33), .ZN(n1901) );
  OAI22_X1 U2016 ( .A1(n1892), .A2(n1285), .B1(n1893), .B2(n1284), .ZN(n1002)
         );
  OAI22_X1 U2017 ( .A1(n1909), .A2(n1366), .B1(n1910), .B2(n1365), .ZN(n1080)
         );
  OAI22_X1 U2018 ( .A1(n1733), .A2(n1283), .B1(n1664), .B2(n1282), .ZN(n1000)
         );
  XOR2_X1 U2019 ( .A(n21), .B(a[4]), .Z(n1464) );
  INV_X1 U2020 ( .A(n291), .ZN(n352) );
  NOR2_X1 U2021 ( .A1(n291), .A2(n294), .ZN(n289) );
  OAI21_X1 U2022 ( .B1(n291), .B2(n295), .A(n292), .ZN(n290) );
  INV_X2 U2023 ( .A(n1906), .ZN(n1905) );
  OAI22_X1 U2024 ( .A1(n1903), .A2(n1338), .B1(n1905), .B2(n1337), .ZN(n1053)
         );
  INV_X1 U2025 ( .A(n42), .ZN(n1895) );
  INV_X2 U2026 ( .A(n1669), .ZN(n1894) );
  OAI21_X1 U2027 ( .B1(n300), .B2(n298), .A(n299), .ZN(n297) );
  AOI21_X1 U2028 ( .B1(n305), .B2(n1839), .A(n302), .ZN(n300) );
  OAI22_X1 U2029 ( .A1(n1904), .A2(n1352), .B1(n1744), .B2(n1351), .ZN(n1067)
         );
  XOR2_X1 U2030 ( .A(n30), .B(a[6]), .Z(n1463) );
  OAI22_X1 U2031 ( .A1(n1778), .A2(n1147), .B1(n1593), .B2(n1146), .ZN(n872)
         );
  OAI22_X1 U2032 ( .A1(n1608), .A2(n1149), .B1(n1148), .B2(n1593), .ZN(n874)
         );
  OAI22_X1 U2033 ( .A1(n1778), .A2(n1148), .B1(n1739), .B2(n1147), .ZN(n873)
         );
  OAI22_X1 U2034 ( .A1(n1151), .A2(n1608), .B1(n1150), .B2(n1739), .ZN(n876)
         );
  INV_X1 U2035 ( .A(n1739), .ZN(n818) );
  OAI22_X1 U2036 ( .A1(n1608), .A2(n1150), .B1(n1739), .B2(n1149), .ZN(n875)
         );
  OAI22_X1 U2037 ( .A1(n102), .A2(n1153), .B1(n1152), .B2(n1739), .ZN(n878) );
  OAI22_X1 U2038 ( .A1(n102), .A2(n819), .B1(n1154), .B2(n1739), .ZN(n847) );
  OAI22_X1 U2039 ( .A1(n1778), .A2(n1152), .B1(n1151), .B2(n1739), .ZN(n877)
         );
  INV_X1 U2040 ( .A(n1938), .ZN(n1935) );
  XNOR2_X1 U2041 ( .A(n1445), .B(n104), .ZN(n1139) );
  XNOR2_X1 U2042 ( .A(n1916), .B(n104), .ZN(n1144) );
  XNOR2_X1 U2043 ( .A(n1447), .B(n104), .ZN(n1141) );
  XNOR2_X1 U2044 ( .A(n1446), .B(n104), .ZN(n1140) );
  INV_X1 U2045 ( .A(n104), .ZN(n817) );
  XNOR2_X1 U2046 ( .A(n1603), .B(n104), .ZN(n1143) );
  XNOR2_X1 U2047 ( .A(n1448), .B(n104), .ZN(n1142) );
  XOR2_X1 U2048 ( .A(n104), .B(a[26]), .Z(n1453) );
  OAI22_X1 U2049 ( .A1(n1717), .A2(n1387), .B1(n1386), .B2(n1914), .ZN(n1100)
         );
  OAI22_X1 U2050 ( .A1(n1912), .A2(n1415), .B1(n1414), .B2(n1914), .ZN(n1128)
         );
  OAI22_X1 U2051 ( .A1(n1912), .A2(n1388), .B1(n1387), .B2(n1828), .ZN(n1101)
         );
  OAI22_X1 U2052 ( .A1(n1717), .A2(n1413), .B1(n1412), .B2(n1829), .ZN(n1126)
         );
  OAI22_X1 U2053 ( .A1(n1717), .A2(n1412), .B1(n1411), .B2(n1829), .ZN(n1125)
         );
  OAI22_X1 U2054 ( .A1(n1912), .A2(n1410), .B1(n1409), .B2(n1828), .ZN(n1123)
         );
  OAI22_X1 U2055 ( .A1(n1717), .A2(n1390), .B1(n1389), .B2(n1914), .ZN(n1103)
         );
  OAI22_X1 U2056 ( .A1(n1912), .A2(n1395), .B1(n1394), .B2(n1914), .ZN(n1108)
         );
  OAI22_X1 U2057 ( .A1(n1717), .A2(n1411), .B1(n1410), .B2(n1829), .ZN(n1124)
         );
  OAI22_X1 U2058 ( .A1(n1717), .A2(n1389), .B1(n1388), .B2(n1829), .ZN(n1102)
         );
  OAI22_X1 U2059 ( .A1(n1717), .A2(n1394), .B1(n1393), .B2(n1828), .ZN(n1107)
         );
  OAI22_X1 U2060 ( .A1(n1717), .A2(n1392), .B1(n1391), .B2(n1914), .ZN(n1105)
         );
  OAI22_X1 U2061 ( .A1(n1717), .A2(n1409), .B1(n1408), .B2(n1914), .ZN(n1122)
         );
  OAI22_X1 U2062 ( .A1(n1913), .A2(n1391), .B1(n1390), .B2(n1828), .ZN(n1104)
         );
  OAI22_X1 U2063 ( .A1(n1912), .A2(n1393), .B1(n1392), .B2(n1829), .ZN(n1106)
         );
  OAI22_X1 U2064 ( .A1(n1397), .A2(n1913), .B1(n1396), .B2(n1914), .ZN(n1110)
         );
  OAI22_X1 U2065 ( .A1(n1717), .A2(n1414), .B1(n1413), .B2(n1828), .ZN(n1127)
         );
  OAI22_X1 U2066 ( .A1(n1912), .A2(n1396), .B1(n1395), .B2(n1828), .ZN(n1109)
         );
  OAI22_X1 U2067 ( .A1(n1717), .A2(n1920), .B1(n1418), .B2(n1914), .ZN(n859)
         );
  NAND2_X1 U2068 ( .A1(n1466), .A2(n6), .ZN(n9) );
  XNOR2_X1 U2069 ( .A(n79), .B(a[20]), .ZN(n89) );
  INV_X2 U2070 ( .A(n1930), .ZN(n1929) );
  XNOR2_X1 U2071 ( .A(n1921), .B(b[28]), .ZN(n1356) );
  XNOR2_X1 U2072 ( .A(n1921), .B(b[26]), .ZN(n1358) );
  XNOR2_X1 U2073 ( .A(n1786), .B(b[27]), .ZN(n1357) );
  XNOR2_X1 U2074 ( .A(n1757), .B(b[25]), .ZN(n1359) );
  XNOR2_X1 U2075 ( .A(n1921), .B(n1427), .ZN(n1361) );
  XNOR2_X1 U2076 ( .A(n1922), .B(b[24]), .ZN(n1360) );
  XNOR2_X1 U2077 ( .A(n1596), .B(n1431), .ZN(n1365) );
  XNOR2_X1 U2078 ( .A(n1591), .B(n1428), .ZN(n1275) );
  XNOR2_X1 U2079 ( .A(n1591), .B(n1444), .ZN(n1291) );
  XNOR2_X1 U2080 ( .A(n1592), .B(n1445), .ZN(n1292) );
  XNOR2_X1 U2081 ( .A(n1592), .B(n1430), .ZN(n1277) );
  XNOR2_X1 U2082 ( .A(n1860), .B(n1429), .ZN(n1276) );
  XNOR2_X1 U2083 ( .A(n1591), .B(n1443), .ZN(n1290) );
  XNOR2_X1 U2084 ( .A(n1860), .B(n1431), .ZN(n1278) );
  NOR2_X1 U2085 ( .A1(n753), .A2(n762), .ZN(n285) );
  NAND2_X1 U2086 ( .A1(n1768), .A2(n264), .ZN(n135) );
  NAND2_X1 U2087 ( .A1(n1129), .A2(n1099), .ZN(n328) );
  OAI22_X1 U2088 ( .A1(n1912), .A2(n1416), .B1(n1415), .B2(n1828), .ZN(n1129)
         );
  NAND2_X1 U2089 ( .A1(n1461), .A2(n1888), .ZN(n53) );
  NAND2_X1 U2090 ( .A1(n753), .A2(n762), .ZN(n286) );
  OAI21_X1 U2091 ( .B1(n184), .B2(n1742), .A(n1620), .ZN(n175) );
  NOR2_X1 U2092 ( .A1(n1740), .A2(n1742), .ZN(n174) );
  NOR2_X1 U2093 ( .A1(n475), .A2(n500), .ZN(n176) );
  XNOR2_X1 U2094 ( .A(n144), .B(n313), .ZN(product[6]) );
  OAI22_X1 U2095 ( .A1(n1733), .A2(n1284), .B1(n1665), .B2(n1283), .ZN(n1001)
         );
  NAND2_X1 U2096 ( .A1(n651), .A2(n668), .ZN(n243) );
  OAI22_X1 U2097 ( .A1(n1891), .A2(n1288), .B1(n1664), .B2(n1287), .ZN(n1005)
         );
  OAI22_X1 U2098 ( .A1(n1733), .A2(n1292), .B1(n1664), .B2(n1291), .ZN(n1009)
         );
  OAI22_X1 U2099 ( .A1(n1733), .A2(n1293), .B1(n1665), .B2(n1292), .ZN(n1010)
         );
  XNOR2_X1 U2100 ( .A(a[16]), .B(n63), .ZN(n74) );
  INV_X1 U2101 ( .A(n1827), .ZN(n217) );
  AOI21_X1 U2102 ( .B1(n1837), .B2(n228), .A(n1881), .ZN(n215) );
  OAI22_X1 U2103 ( .A1(n1892), .A2(n1287), .B1(n1893), .B2(n1286), .ZN(n1004)
         );
  NOR2_X1 U2104 ( .A1(n811), .A2(n1128), .ZN(n322) );
  OAI22_X1 U2105 ( .A1(n1896), .A2(n1317), .B1(n1729), .B2(n1316), .ZN(n1033)
         );
  OAI22_X1 U2106 ( .A1(n1897), .A2(n1314), .B1(n1900), .B2(n1313), .ZN(n1030)
         );
  OAI22_X1 U2107 ( .A1(n1898), .A2(n1321), .B1(n1728), .B2(n1320), .ZN(n1037)
         );
  OAI21_X1 U2108 ( .B1(n314), .B2(n316), .A(n315), .ZN(n313) );
  OAI22_X1 U2109 ( .A1(n1897), .A2(n1315), .B1(n1899), .B2(n1314), .ZN(n1031)
         );
  INV_X1 U2110 ( .A(n312), .ZN(n310) );
  AOI21_X1 U2111 ( .B1(n287), .B2(n1727), .A(n1732), .ZN(n277) );
  OAI21_X1 U2112 ( .B1(n195), .B2(n167), .A(n168), .ZN(n166) );
  OAI21_X1 U2113 ( .B1(n1597), .B2(n286), .A(n281), .ZN(n279) );
  INV_X1 U2114 ( .A(n1598), .ZN(n350) );
  CLKBUF_X1 U2115 ( .A(n305), .Z(n1872) );
  XNOR2_X1 U2116 ( .A(n1863), .B(a[18]), .ZN(n1874) );
  AOI21_X1 U2117 ( .B1(n1589), .B2(n1698), .A(n1712), .ZN(n1878) );
  INV_X1 U2118 ( .A(n276), .ZN(n274) );
  NAND2_X1 U2119 ( .A1(n1880), .A2(n248), .ZN(n132) );
  OAI21_X1 U2120 ( .B1(n1818), .B2(n248), .A(n243), .ZN(n241) );
  NAND2_X1 U2121 ( .A1(n669), .A2(n684), .ZN(n248) );
  NAND2_X1 U2122 ( .A1(n240), .A2(n1662), .ZN(n233) );
  NOR2_X1 U2123 ( .A1(n242), .A2(n247), .ZN(n240) );
  INV_X1 U2124 ( .A(n1833), .ZN(n1879) );
  OAI22_X1 U2125 ( .A1(n1903), .A2(n1337), .B1(n1905), .B2(n1336), .ZN(n1052)
         );
  AOI21_X1 U2126 ( .B1(n1842), .B2(n313), .A(n310), .ZN(n308) );
  OR2_X1 U2127 ( .A1(n669), .A2(n684), .ZN(n1880) );
  AOI21_X1 U2128 ( .B1(n1882), .B2(n1698), .A(n1752), .ZN(n257) );
  NAND2_X1 U2129 ( .A1(n278), .A2(n1838), .ZN(n271) );
  OAI22_X1 U2130 ( .A1(n1769), .A2(n1377), .B1(n1699), .B2(n1376), .ZN(n1091)
         );
  OAI22_X1 U2131 ( .A1(n1907), .A2(n1361), .B1(n1753), .B2(n1360), .ZN(n1075)
         );
  OAI22_X1 U2132 ( .A1(n1908), .A2(n1375), .B1(n1753), .B2(n1374), .ZN(n1089)
         );
  OAI22_X1 U2133 ( .A1(n1907), .A2(n1374), .B1(n1753), .B2(n1373), .ZN(n1088)
         );
  OR2_X1 U2134 ( .A1(n1915), .A2(n1485), .ZN(n1250) );
  AND2_X1 U2135 ( .A1(n1916), .A2(n1812), .ZN(n949) );
  AOI21_X1 U2136 ( .B1(n1835), .B2(n163), .A(n158), .ZN(n156) );
  NAND2_X1 U2137 ( .A1(n449), .A2(n474), .ZN(n172) );
  OAI21_X1 U2138 ( .B1(n269), .B2(n263), .A(n264), .ZN(n262) );
  NOR2_X1 U2139 ( .A1(n715), .A2(n728), .ZN(n263) );
  OAI21_X1 U2140 ( .B1(n257), .B2(n253), .A(n254), .ZN(n252) );
  NAND2_X1 U2141 ( .A1(n1708), .A2(n223), .ZN(n128) );
  NAND2_X1 U2142 ( .A1(n1837), .A2(n1788), .ZN(n214) );
  INV_X1 U2143 ( .A(n226), .ZN(n228) );
  NAND2_X1 U2144 ( .A1(n613), .A2(n632), .ZN(n226) );
  AND2_X1 U2145 ( .A1(n593), .A2(n612), .ZN(n1881) );
  OAI21_X1 U2146 ( .B1(n250), .B2(n233), .A(n234), .ZN(n232) );
  NAND2_X1 U2147 ( .A1(n1831), .A2(n165), .ZN(n121) );
  NAND2_X1 U2148 ( .A1(n1662), .A2(n238), .ZN(n130) );
  AOI21_X1 U2149 ( .B1(n251), .B2(n270), .A(n252), .ZN(n250) );
  OAI21_X1 U2150 ( .B1(n271), .B2(n288), .A(n272), .ZN(n270) );
  AOI21_X1 U2151 ( .B1(n279), .B2(n1838), .A(n274), .ZN(n272) );
  NOR2_X1 U2152 ( .A1(n669), .A2(n684), .ZN(n247) );
  XNOR2_X1 U2153 ( .A(n1746), .B(n1915), .ZN(n1353) );
  XNOR2_X1 U2154 ( .A(n1925), .B(n1442), .ZN(n1345) );
  XNOR2_X1 U2155 ( .A(n1746), .B(n1438), .ZN(n1341) );
  XNOR2_X1 U2156 ( .A(n1750), .B(n1441), .ZN(n1344) );
  XNOR2_X1 U2157 ( .A(n1751), .B(n1437), .ZN(n1340) );
  XNOR2_X1 U2158 ( .A(n1750), .B(n1436), .ZN(n1339) );
  XNOR2_X1 U2159 ( .A(n1745), .B(n1440), .ZN(n1343) );
  XNOR2_X1 U2160 ( .A(n1925), .B(n1439), .ZN(n1342) );
  NAND2_X1 U2161 ( .A1(n1589), .A2(n261), .ZN(n134) );
  NAND2_X1 U2162 ( .A1(n1697), .A2(n714), .ZN(n261) );
  NOR2_X1 U2163 ( .A1(n214), .A2(n198), .ZN(n196) );
  XNOR2_X1 U2164 ( .A(n1872), .B(n142), .ZN(product[8]) );
  NAND2_X1 U2165 ( .A1(n805), .A2(n808), .ZN(n315) );
  NOR2_X1 U2166 ( .A1(n805), .A2(n808), .ZN(n314) );
  AOI21_X1 U2167 ( .B1(n1832), .B2(n1833), .A(n1650), .ZN(n199) );
  AOI21_X1 U2168 ( .B1(n182), .B2(n1804), .A(n170), .ZN(n168) );
  INV_X1 U2169 ( .A(n1588), .ZN(n184) );
  NOR2_X1 U2170 ( .A1(n525), .A2(n548), .ZN(n192) );
  OAI22_X1 U2171 ( .A1(n1722), .A2(n1156), .B1(n1706), .B2(n1155), .ZN(n880)
         );
  OAI22_X1 U2172 ( .A1(n1722), .A2(n1159), .B1(n1706), .B2(n1158), .ZN(n883)
         );
  OAI22_X1 U2173 ( .A1(n1722), .A2(n1158), .B1(n1706), .B2(n1157), .ZN(n882)
         );
  OAI22_X1 U2174 ( .A1(n1722), .A2(n1157), .B1(n1706), .B2(n1156), .ZN(n881)
         );
  OAI22_X1 U2175 ( .A1(n1722), .A2(n1160), .B1(n1706), .B2(n1159), .ZN(n884)
         );
  XNOR2_X1 U2176 ( .A(n1743), .B(n1439), .ZN(n1166) );
  OAI22_X1 U2177 ( .A1(n97), .A2(n1161), .B1(n1706), .B2(n1160), .ZN(n885) );
  OAI22_X1 U2178 ( .A1(n1722), .A2(n1163), .B1(n1706), .B2(n1162), .ZN(n887)
         );
  OAI22_X1 U2179 ( .A1(n1722), .A2(n1162), .B1(n1706), .B2(n1161), .ZN(n886)
         );
  OAI22_X1 U2180 ( .A1(n97), .A2(n1164), .B1(n1706), .B2(n1163), .ZN(n888) );
  OAI22_X1 U2181 ( .A1(n97), .A2(n1480), .B1(n1165), .B2(n1706), .ZN(n848) );
  XNOR2_X1 U2182 ( .A(n1743), .B(n1442), .ZN(n1169) );
  XNOR2_X1 U2183 ( .A(n1743), .B(n1441), .ZN(n1168) );
  XNOR2_X1 U2184 ( .A(n1743), .B(n1440), .ZN(n1167) );
  XNOR2_X1 U2185 ( .A(n1743), .B(n1443), .ZN(n1170) );
  XNOR2_X1 U2186 ( .A(n1743), .B(n1444), .ZN(n1171) );
  XNOR2_X1 U2187 ( .A(n1743), .B(n1445), .ZN(n1172) );
  XNOR2_X1 U2188 ( .A(n1743), .B(n1447), .ZN(n1174) );
  XNOR2_X1 U2189 ( .A(n1743), .B(n1446), .ZN(n1173) );
  XNOR2_X1 U2190 ( .A(n1917), .B(n1743), .ZN(n1177) );
  XNOR2_X1 U2191 ( .A(n1743), .B(n1603), .ZN(n1176) );
  XNOR2_X1 U2192 ( .A(n1743), .B(n1448), .ZN(n1175) );
  INV_X1 U2193 ( .A(n1743), .ZN(n1481) );
  XOR2_X1 U2194 ( .A(n1856), .B(a[20]), .Z(n1456) );
  OR2_X1 U2195 ( .A1(n1916), .A2(n1762), .ZN(n1273) );
  XOR2_X1 U2196 ( .A(n308), .B(n143), .Z(product[7]) );
  OAI21_X1 U2197 ( .B1(n308), .B2(n306), .A(n307), .ZN(n305) );
  OAI22_X1 U2198 ( .A1(n1907), .A2(n1379), .B1(n1699), .B2(n1378), .ZN(n1093)
         );
  OAI22_X1 U2199 ( .A1(n1769), .A2(n1378), .B1(n1699), .B2(n1377), .ZN(n1092)
         );
  OAI22_X1 U2200 ( .A1(n1908), .A2(n1380), .B1(n1753), .B2(n1379), .ZN(n1094)
         );
  OAI22_X1 U2201 ( .A1(n1769), .A2(n1382), .B1(n1699), .B2(n1381), .ZN(n1096)
         );
  OAI22_X1 U2202 ( .A1(n1769), .A2(n1370), .B1(n1753), .B2(n1369), .ZN(n1084)
         );
  OAI22_X1 U2203 ( .A1(n1769), .A2(n1371), .B1(n1678), .B2(n1370), .ZN(n1085)
         );
  OAI22_X1 U2204 ( .A1(n1769), .A2(n1373), .B1(n1753), .B2(n1372), .ZN(n1087)
         );
  OAI22_X1 U2205 ( .A1(n1909), .A2(n1369), .B1(n1910), .B2(n1368), .ZN(n1083)
         );
  OAI22_X1 U2206 ( .A1(n1769), .A2(n1372), .B1(n1678), .B2(n1371), .ZN(n1086)
         );
  OAI22_X1 U2207 ( .A1(n1907), .A2(n1384), .B1(n1753), .B2(n1383), .ZN(n1098)
         );
  OAI22_X1 U2208 ( .A1(n1908), .A2(n1381), .B1(n1753), .B2(n1380), .ZN(n1095)
         );
  OAI22_X1 U2209 ( .A1(n1769), .A2(n1383), .B1(n1753), .B2(n1382), .ZN(n1097)
         );
  XNOR2_X1 U2210 ( .A(n880), .B(n1883), .ZN(n386) );
  XNOR2_X1 U2211 ( .A(n950), .B(n916), .ZN(n1883) );
  XNOR2_X1 U2212 ( .A(n1884), .B(n390), .ZN(n380) );
  XNOR2_X1 U2213 ( .A(n388), .B(n386), .ZN(n1884) );
  XNOR2_X1 U2214 ( .A(n412), .B(n1885), .ZN(n374) );
  XNOR2_X1 U2215 ( .A(n380), .B(n410), .ZN(n1885) );
  XNOR2_X1 U2216 ( .A(n224), .B(n128), .ZN(product[22]) );
  OAI21_X1 U2217 ( .B1(n1600), .B2(n225), .A(n226), .ZN(n224) );
  OAI21_X1 U2218 ( .B1(n231), .B2(n1668), .A(n1599), .ZN(n213) );
  OAI21_X1 U2219 ( .B1(n231), .B2(n205), .A(n206), .ZN(n204) );
  INV_X1 U2220 ( .A(n1766), .ZN(n231) );
  NAND2_X1 U2221 ( .A1(n1723), .A2(n1768), .ZN(n256) );
  NAND2_X1 U2222 ( .A1(n169), .A2(n181), .ZN(n167) );
  NOR2_X1 U2223 ( .A1(n176), .A2(n171), .ZN(n169) );
  XNOR2_X1 U2224 ( .A(n1860), .B(n1427), .ZN(n1274) );
  OAI22_X1 U2225 ( .A1(n1867), .A2(n1252), .B1(n1889), .B2(n1251), .ZN(n970)
         );
  OAI22_X1 U2226 ( .A1(n1693), .A2(n1253), .B1(n1889), .B2(n1252), .ZN(n971)
         );
  OAI22_X1 U2227 ( .A1(n1868), .A2(n1266), .B1(n1889), .B2(n1265), .ZN(n984)
         );
  OAI22_X1 U2228 ( .A1(n1693), .A2(n1259), .B1(n1889), .B2(n1258), .ZN(n977)
         );
  OAI22_X1 U2229 ( .A1(n1868), .A2(n1254), .B1(n1889), .B2(n1253), .ZN(n972)
         );
  OAI22_X1 U2230 ( .A1(n1868), .A2(n1255), .B1(n1889), .B2(n1254), .ZN(n973)
         );
  OAI22_X1 U2231 ( .A1(n1693), .A2(n1260), .B1(n1889), .B2(n1259), .ZN(n978)
         );
  OAI22_X1 U2232 ( .A1(n1693), .A2(n1262), .B1(n1889), .B2(n1261), .ZN(n980)
         );
  XNOR2_X1 U2233 ( .A(n1860), .B(n1915), .ZN(n1297) );
  XNOR2_X1 U2234 ( .A(n1933), .B(n1441), .ZN(n1288) );
  OAI22_X1 U2235 ( .A1(n1693), .A2(n1256), .B1(n1889), .B2(n1255), .ZN(n974)
         );
  OAI22_X1 U2236 ( .A1(n1868), .A2(n1264), .B1(n1889), .B2(n1263), .ZN(n982)
         );
  OAI22_X1 U2237 ( .A1(n1868), .A2(n1263), .B1(n1889), .B2(n1262), .ZN(n981)
         );
  OAI22_X1 U2238 ( .A1(n1693), .A2(n1267), .B1(n1889), .B2(n1266), .ZN(n985)
         );
  OAI22_X1 U2239 ( .A1(n1693), .A2(n1257), .B1(n1889), .B2(n1256), .ZN(n975)
         );
  OAI22_X1 U2240 ( .A1(n1868), .A2(n1270), .B1(n1889), .B2(n1269), .ZN(n988)
         );
  OAI22_X1 U2241 ( .A1(n1693), .A2(n1271), .B1(n1889), .B2(n1270), .ZN(n989)
         );
  OAI22_X1 U2242 ( .A1(n1693), .A2(n1261), .B1(n1889), .B2(n1260), .ZN(n979)
         );
  OAI22_X1 U2243 ( .A1(n1868), .A2(n1258), .B1(n1889), .B2(n1257), .ZN(n976)
         );
  OAI22_X1 U2244 ( .A1(n1868), .A2(n1265), .B1(n1889), .B2(n1264), .ZN(n983)
         );
  OAI22_X1 U2245 ( .A1(n1868), .A2(n1272), .B1(n1889), .B2(n1271), .ZN(n990)
         );
  OAI22_X1 U2246 ( .A1(n1693), .A2(n1762), .B1(n1273), .B2(n1889), .ZN(n854)
         );
  OAI22_X1 U2247 ( .A1(n1867), .A2(n1269), .B1(n1798), .B2(n1889), .ZN(n987)
         );
  OAI22_X1 U2248 ( .A1(n1867), .A2(n1798), .B1(n1267), .B2(n1889), .ZN(n986)
         );
  XNOR2_X1 U2249 ( .A(n1933), .B(n1603), .ZN(n1296) );
  XNOR2_X1 U2250 ( .A(n1718), .B(n1442), .ZN(n1289) );
  XNOR2_X1 U2251 ( .A(n1933), .B(n1756), .ZN(n1293) );
  XNOR2_X1 U2252 ( .A(n1933), .B(n1448), .ZN(n1295) );
  XNOR2_X1 U2253 ( .A(n1933), .B(n1447), .ZN(n1294) );
  XNOR2_X1 U2254 ( .A(n39), .B(a[10]), .ZN(n50) );
  XNOR2_X1 U2255 ( .A(n1886), .B(n402), .ZN(n367) );
  XNOR2_X1 U2256 ( .A(n374), .B(n369), .ZN(n1886) );
  XNOR2_X1 U2257 ( .A(n1887), .B(n398), .ZN(n365) );
  XNOR2_X1 U2258 ( .A(n367), .B(n372), .ZN(n1887) );
  INV_X1 U2259 ( .A(n297), .ZN(n296) );
  AOI21_X1 U2260 ( .B1(n289), .B2(n297), .A(n290), .ZN(n288) );
  OR2_X1 U2261 ( .A1(n1916), .A2(n1713), .ZN(n1385) );
  INV_X1 U2262 ( .A(n24), .ZN(n1906) );
  OAI21_X1 U2263 ( .B1(n1716), .B2(n179), .A(n172), .ZN(n170) );
  NOR2_X1 U2264 ( .A1(n1680), .A2(n474), .ZN(n171) );
  XNOR2_X1 U2265 ( .A(n1936), .B(n1429), .ZN(n1251) );
  XNOR2_X1 U2266 ( .A(n1936), .B(n1441), .ZN(n1263) );
  XNOR2_X1 U2267 ( .A(n1937), .B(n1440), .ZN(n1262) );
  XNOR2_X1 U2268 ( .A(n1936), .B(n1915), .ZN(n1272) );
  XNOR2_X1 U2269 ( .A(n1937), .B(n1439), .ZN(n1261) );
  XNOR2_X1 U2270 ( .A(n1936), .B(n1442), .ZN(n1264) );
  XNOR2_X1 U2271 ( .A(n1937), .B(n1603), .ZN(n1271) );
  XNOR2_X1 U2272 ( .A(n1937), .B(n1447), .ZN(n1269) );
  AOI21_X1 U2273 ( .B1(n249), .B2(n1755), .A(n1741), .ZN(n239) );
  AOI21_X1 U2274 ( .B1(n232), .B2(n196), .A(n197), .ZN(n195) );
  AOI21_X1 U2275 ( .B1(n241), .B2(n1662), .A(n1701), .ZN(n234) );
  OAI22_X1 U2276 ( .A1(n1898), .A2(n1300), .B1(n1785), .B2(n1299), .ZN(n1016)
         );
  OAI22_X1 U2277 ( .A1(n1896), .A2(n1301), .B1(n1785), .B2(n1300), .ZN(n1017)
         );
  OAI22_X1 U2278 ( .A1(n1896), .A2(n1302), .B1(n1900), .B2(n1301), .ZN(n1018)
         );
  OAI22_X1 U2279 ( .A1(n1898), .A2(n1303), .B1(n1729), .B2(n1302), .ZN(n1019)
         );
  OAI22_X1 U2280 ( .A1(n1896), .A2(n1304), .B1(n1728), .B2(n1303), .ZN(n1020)
         );
  OAI22_X1 U2281 ( .A1(n1896), .A2(n1320), .B1(n1900), .B2(n1319), .ZN(n1036)
         );
  OAI22_X1 U2282 ( .A1(n1896), .A2(n1319), .B1(n1729), .B2(n1318), .ZN(n1035)
         );
  OAI22_X1 U2283 ( .A1(n1898), .A2(n1318), .B1(n1728), .B2(n1317), .ZN(n1034)
         );
  OAI22_X1 U2284 ( .A1(n1896), .A2(n1930), .B1(n1325), .B2(n1900), .ZN(n856)
         );
  OAI22_X1 U2285 ( .A1(n1897), .A2(n1316), .B1(n1899), .B2(n1315), .ZN(n1032)
         );
  NAND2_X1 U2286 ( .A1(n1463), .A2(n33), .ZN(n36) );
  OAI22_X1 U2287 ( .A1(n1891), .A2(n1275), .B1(n1726), .B2(n1274), .ZN(n992)
         );
  XNOR2_X1 U2288 ( .A(n1792), .B(b[25]), .ZN(n1299) );
  OAI22_X1 U2289 ( .A1(n1733), .A2(n1276), .B1(n1275), .B2(n1894), .ZN(n993)
         );
  OAI22_X1 U2290 ( .A1(n1891), .A2(n1289), .B1(n1894), .B2(n1288), .ZN(n1006)
         );
  OAI22_X1 U2291 ( .A1(n1733), .A2(n1291), .B1(n1894), .B2(n1770), .ZN(n1008)
         );
  OAI22_X1 U2292 ( .A1(n1891), .A2(n1277), .B1(n1894), .B2(n1276), .ZN(n994)
         );
  OAI22_X1 U2293 ( .A1(n1891), .A2(n1725), .B1(n1298), .B2(n1894), .ZN(n855)
         );
  OAI22_X1 U2294 ( .A1(n1891), .A2(n1294), .B1(n1894), .B2(n1293), .ZN(n1011)
         );
  OAI22_X1 U2295 ( .A1(n1733), .A2(n1296), .B1(n1894), .B2(n1295), .ZN(n1013)
         );
  OAI22_X1 U2296 ( .A1(n1891), .A2(n1290), .B1(n1894), .B2(n1289), .ZN(n1007)
         );
  OAI22_X1 U2297 ( .A1(n1733), .A2(n1295), .B1(n1894), .B2(n1294), .ZN(n1012)
         );
  XNOR2_X1 U2298 ( .A(n1929), .B(n1447), .ZN(n1321) );
  XNOR2_X1 U2299 ( .A(n1929), .B(n1448), .ZN(n1322) );
  XNOR2_X1 U2300 ( .A(n1929), .B(n1756), .ZN(n1320) );
  XNOR2_X1 U2301 ( .A(n1929), .B(n1445), .ZN(n1319) );
  XNOR2_X1 U2302 ( .A(n1792), .B(n1916), .ZN(n1324) );
  XNOR2_X1 U2303 ( .A(n1929), .B(n1444), .ZN(n1318) );
  XNOR2_X1 U2304 ( .A(n1929), .B(n1603), .ZN(n1323) );
  NAND2_X1 U2305 ( .A1(n1462), .A2(n1726), .ZN(n44) );
  XNOR2_X1 U2306 ( .A(n30), .B(a[8]), .ZN(n42) );
  INV_X1 U2307 ( .A(n1730), .ZN(n344) );
  NOR2_X1 U2308 ( .A1(n668), .A2(n651), .ZN(n242) );
  XNOR2_X1 U2309 ( .A(n1863), .B(n1447), .ZN(n1206) );
  XNOR2_X1 U2310 ( .A(n1863), .B(n1448), .ZN(n1207) );
  XNOR2_X1 U2311 ( .A(n1864), .B(n1435), .ZN(n1194) );
  XNOR2_X1 U2312 ( .A(n1864), .B(n1436), .ZN(n1195) );
  XOR2_X1 U2313 ( .A(n145), .B(n316), .Z(product[5]) );
  AOI21_X1 U2314 ( .B1(n1844), .B2(n321), .A(n318), .ZN(n316) );
  OAI22_X1 U2315 ( .A1(n1787), .A2(n1170), .B1(n1711), .B2(n1169), .ZN(n893)
         );
  OAI22_X1 U2316 ( .A1(n1787), .A2(n1169), .B1(n1711), .B2(n1168), .ZN(n892)
         );
  OAI22_X1 U2317 ( .A1(n1787), .A2(n1168), .B1(n1711), .B2(n1167), .ZN(n891)
         );
  OAI22_X1 U2318 ( .A1(n1787), .A2(n1167), .B1(n1711), .B2(n1166), .ZN(n890)
         );
  OAI22_X1 U2319 ( .A1(n1787), .A2(n1175), .B1(n1711), .B2(n1174), .ZN(n898)
         );
  OAI22_X1 U2320 ( .A1(n1787), .A2(n1171), .B1(n1711), .B2(n1170), .ZN(n894)
         );
  OAI22_X1 U2321 ( .A1(n1627), .A2(n1174), .B1(n1711), .B2(n1173), .ZN(n897)
         );
  OAI22_X1 U2322 ( .A1(n1627), .A2(n1173), .B1(n1865), .B2(n1172), .ZN(n896)
         );
  OAI22_X1 U2323 ( .A1(n1787), .A2(n1176), .B1(n1711), .B2(n1175), .ZN(n899)
         );
  XNOR2_X1 U2324 ( .A(n1799), .B(n1440), .ZN(n1182) );
  OAI22_X1 U2325 ( .A1(n1627), .A2(n1172), .B1(n1865), .B2(n1171), .ZN(n895)
         );
  XNOR2_X1 U2326 ( .A(n1799), .B(n1439), .ZN(n1181) );
  OAI22_X1 U2327 ( .A1(n91), .A2(n1177), .B1(n1865), .B2(n1176), .ZN(n900) );
  OAI22_X1 U2328 ( .A1(n91), .A2(n1481), .B1(n1178), .B2(n1865), .ZN(n849) );
  XNOR2_X1 U2329 ( .A(n1780), .B(n1445), .ZN(n1187) );
  XNOR2_X1 U2330 ( .A(n1780), .B(n1446), .ZN(n1188) );
  INV_X1 U2331 ( .A(n79), .ZN(n1482) );
  XNOR2_X1 U2332 ( .A(n1780), .B(n1441), .ZN(n1183) );
  XNOR2_X1 U2333 ( .A(n1649), .B(n1447), .ZN(n1189) );
  XNOR2_X1 U2334 ( .A(n1799), .B(n1438), .ZN(n1180) );
  XNOR2_X1 U2335 ( .A(n1784), .B(n1437), .ZN(n1179) );
  XNOR2_X1 U2336 ( .A(n1784), .B(n1444), .ZN(n1186) );
  XNOR2_X1 U2337 ( .A(n1603), .B(n1715), .ZN(n1191) );
  XNOR2_X1 U2338 ( .A(n1715), .B(n1443), .ZN(n1185) );
  XNOR2_X1 U2339 ( .A(n1649), .B(n1448), .ZN(n1190) );
  XNOR2_X1 U2340 ( .A(n1748), .B(b[30]), .ZN(n1387) );
  XNOR2_X1 U2341 ( .A(n1748), .B(b[28]), .ZN(n1389) );
  XNOR2_X1 U2342 ( .A(n1748), .B(b[29]), .ZN(n1388) );
  NAND2_X1 U2343 ( .A1(n1130), .A2(n859), .ZN(n331) );
  XNOR2_X1 U2344 ( .A(n1771), .B(b[27]), .ZN(n1390) );
  XNOR2_X1 U2345 ( .A(n1771), .B(b[26]), .ZN(n1391) );
  XNOR2_X1 U2346 ( .A(n1748), .B(b[25]), .ZN(n1392) );
  XNOR2_X1 U2347 ( .A(n1918), .B(n1431), .ZN(n1398) );
  XOR2_X1 U2348 ( .A(n3), .B(n842), .Z(n1466) );
  NAND2_X1 U2349 ( .A1(n360), .A2(n323), .ZN(n147) );
  INV_X1 U2350 ( .A(n195), .ZN(n194) );
  INV_X1 U2351 ( .A(n1805), .ZN(n249) );
  XNOR2_X1 U2352 ( .A(n1748), .B(b[31]), .ZN(n1386) );
  XNOR2_X1 U2353 ( .A(n1748), .B(n1441), .ZN(n1408) );
  XNOR2_X1 U2354 ( .A(n1749), .B(n1442), .ZN(n1409) );
  XNOR2_X1 U2355 ( .A(n1749), .B(n1440), .ZN(n1407) );
  XNOR2_X1 U2356 ( .A(n1772), .B(n1447), .ZN(n1414) );
  XNOR2_X1 U2357 ( .A(n1772), .B(n1915), .ZN(n1417) );
  XNOR2_X1 U2358 ( .A(n1749), .B(n1448), .ZN(n1415) );
  XNOR2_X1 U2359 ( .A(n1749), .B(n1603), .ZN(n1416) );
  XNOR2_X1 U2360 ( .A(n3), .B(a[2]), .ZN(n15) );
  XNOR2_X1 U2361 ( .A(n1777), .B(n1436), .ZN(n1214) );
  XNOR2_X1 U2362 ( .A(n1777), .B(n1435), .ZN(n1213) );
  XNOR2_X1 U2363 ( .A(n1776), .B(n1441), .ZN(n1219) );
  XNOR2_X1 U2364 ( .A(n1777), .B(n1440), .ZN(n1218) );
  XNOR2_X1 U2365 ( .A(n1776), .B(n1438), .ZN(n1216) );
  XNOR2_X1 U2366 ( .A(n1777), .B(n1439), .ZN(n1217) );
  XNOR2_X1 U2367 ( .A(n1777), .B(n1437), .ZN(n1215) );
  XNOR2_X1 U2368 ( .A(n1776), .B(n1442), .ZN(n1220) );
  XNOR2_X1 U2369 ( .A(n1776), .B(n1443), .ZN(n1221) );
  INV_X1 U2370 ( .A(n1777), .ZN(n1484) );
  XNOR2_X1 U2371 ( .A(n1915), .B(n1776), .ZN(n1228) );
  XNOR2_X1 U2372 ( .A(n1777), .B(n1434), .ZN(n1212) );
  XNOR2_X1 U2373 ( .A(n1776), .B(n1447), .ZN(n1225) );
  XNOR2_X1 U2374 ( .A(n1776), .B(n1433), .ZN(n1211) );
  XNOR2_X1 U2375 ( .A(n1776), .B(n1445), .ZN(n1223) );
  XNOR2_X1 U2376 ( .A(n1776), .B(n1448), .ZN(n1226) );
  XNOR2_X1 U2377 ( .A(n1776), .B(n1603), .ZN(n1227) );
  XNOR2_X1 U2378 ( .A(n1776), .B(n1446), .ZN(n1224) );
  XNOR2_X1 U2379 ( .A(n1777), .B(n1444), .ZN(n1222) );
  OAI21_X1 U2380 ( .B1(n215), .B2(n198), .A(n199), .ZN(n197) );
  NOR2_X1 U2381 ( .A1(n256), .A2(n253), .ZN(n251) );
  XOR2_X1 U2382 ( .A(n300), .B(n141), .Z(product[9]) );
  INV_X1 U2383 ( .A(n1670), .ZN(n269) );
  OAI22_X1 U2384 ( .A1(n1904), .A2(n1327), .B1(n1905), .B2(n1326), .ZN(n1042)
         );
  OAI22_X1 U2385 ( .A1(n1904), .A2(n1328), .B1(n1744), .B2(n1327), .ZN(n1043)
         );
  OAI22_X1 U2386 ( .A1(n1904), .A2(n1330), .B1(n1905), .B2(n1329), .ZN(n1045)
         );
  OAI22_X1 U2387 ( .A1(n1902), .A2(n1329), .B1(n1905), .B2(n1328), .ZN(n1044)
         );
  OAI22_X1 U2388 ( .A1(n1904), .A2(n1346), .B1(n1744), .B2(n1345), .ZN(n1061)
         );
  OAI22_X1 U2389 ( .A1(n1904), .A2(n1331), .B1(n1905), .B2(n1330), .ZN(n1046)
         );
  OAI22_X1 U2390 ( .A1(n1902), .A2(n1347), .B1(n1744), .B2(n1346), .ZN(n1062)
         );
  OAI22_X1 U2391 ( .A1(n1903), .A2(n1333), .B1(n1905), .B2(n1332), .ZN(n1048)
         );
  OAI22_X1 U2392 ( .A1(n1902), .A2(n1345), .B1(n1744), .B2(n1344), .ZN(n1060)
         );
  XNOR2_X1 U2393 ( .A(n1786), .B(n1442), .ZN(n1376) );
  XNOR2_X1 U2394 ( .A(n1596), .B(n1441), .ZN(n1375) );
  XNOR2_X1 U2395 ( .A(n1757), .B(n1440), .ZN(n1374) );
  XNOR2_X1 U2396 ( .A(n1921), .B(n1439), .ZN(n1373) );
  OAI22_X1 U2397 ( .A1(n1902), .A2(n1926), .B1(n1354), .B2(n1905), .ZN(n857)
         );
  XNOR2_X1 U2398 ( .A(n1786), .B(n1438), .ZN(n1372) );
  XNOR2_X1 U2399 ( .A(n1922), .B(n1916), .ZN(n1384) );
  XNOR2_X1 U2400 ( .A(n1922), .B(n1448), .ZN(n1382) );
  XNOR2_X1 U2401 ( .A(n1922), .B(n1603), .ZN(n1383) );
  NAND2_X1 U2402 ( .A1(n1464), .A2(n24), .ZN(n27) );
  OAI22_X1 U2403 ( .A1(n1817), .A2(n1183), .B1(n1873), .B2(n1182), .ZN(n905)
         );
  OAI22_X1 U2404 ( .A1(n1817), .A2(n1182), .B1(n1874), .B2(n1181), .ZN(n904)
         );
  OAI22_X1 U2405 ( .A1(n1817), .A2(n1181), .B1(n1702), .B2(n1180), .ZN(n903)
         );
  OAI22_X1 U2406 ( .A1(n1817), .A2(n1188), .B1(n1874), .B2(n1187), .ZN(n910)
         );
  OAI22_X1 U2407 ( .A1(n1817), .A2(n1185), .B1(n1702), .B2(n1184), .ZN(n907)
         );
  OAI22_X1 U2408 ( .A1(n1187), .A2(n1817), .B1(n1873), .B2(n1186), .ZN(n909)
         );
  OAI22_X1 U2409 ( .A1(n1817), .A2(n1184), .B1(n1702), .B2(n1183), .ZN(n906)
         );
  OAI22_X1 U2410 ( .A1(n84), .A2(n1192), .B1(n1702), .B2(n1191), .ZN(n914) );
  OAI22_X1 U2411 ( .A1(n1817), .A2(n1180), .B1(n1874), .B2(n1179), .ZN(n902)
         );
  OAI22_X1 U2412 ( .A1(n1482), .A2(n84), .B1(n1193), .B2(n1874), .ZN(n850) );
  OAI22_X1 U2413 ( .A1(n1186), .A2(n84), .B1(n1873), .B2(n1185), .ZN(n908) );
  OAI22_X1 U2414 ( .A1(n84), .A2(n1190), .B1(n1764), .B2(n1189), .ZN(n912) );
  INV_X1 U2415 ( .A(n1764), .ZN(n824) );
  OAI22_X1 U2416 ( .A1(n1817), .A2(n1189), .B1(n1873), .B2(n1188), .ZN(n911)
         );
  OAI22_X1 U2417 ( .A1(n84), .A2(n1191), .B1(n1764), .B2(n1190), .ZN(n913) );
  OAI21_X1 U2418 ( .B1(n269), .B2(n256), .A(n1878), .ZN(n255) );
  OAI22_X1 U2419 ( .A1(n1854), .A2(n1233), .B1(n1694), .B2(n1232), .ZN(n952)
         );
  OAI22_X1 U2420 ( .A1(n1855), .A2(n1234), .B1(n1618), .B2(n1233), .ZN(n953)
         );
  OAI22_X1 U2421 ( .A1(n1854), .A2(n1232), .B1(n1695), .B2(n1231), .ZN(n951)
         );
  OAI22_X1 U2422 ( .A1(n1854), .A2(n1239), .B1(n1618), .B2(n1238), .ZN(n958)
         );
  OAI22_X1 U2423 ( .A1(n1854), .A2(n1235), .B1(n1619), .B2(n1234), .ZN(n954)
         );
  OAI22_X1 U2424 ( .A1(n1854), .A2(n1236), .B1(n1694), .B2(n1235), .ZN(n955)
         );
  OAI22_X1 U2425 ( .A1(n1854), .A2(n1238), .B1(n1694), .B2(n1237), .ZN(n957)
         );
  OAI22_X1 U2426 ( .A1(n1854), .A2(n1245), .B1(n1618), .B2(n1244), .ZN(n964)
         );
  OAI22_X1 U2427 ( .A1(n1854), .A2(n1241), .B1(n1695), .B2(n1240), .ZN(n960)
         );
  OAI22_X1 U2428 ( .A1(n1609), .A2(n1237), .B1(n1694), .B2(n1236), .ZN(n956)
         );
  OAI22_X1 U2429 ( .A1(n1854), .A2(n1231), .B1(n1695), .B2(n1230), .ZN(n950)
         );
  OAI22_X1 U2430 ( .A1(n1609), .A2(n1243), .B1(n1619), .B2(n1242), .ZN(n962)
         );
  OAI22_X1 U2431 ( .A1(n1609), .A2(n1240), .B1(n1619), .B2(n1239), .ZN(n959)
         );
  OAI22_X1 U2432 ( .A1(n1854), .A2(n1244), .B1(n1619), .B2(n1243), .ZN(n963)
         );
  OAI22_X1 U2433 ( .A1(n1609), .A2(n1242), .B1(n1618), .B2(n1241), .ZN(n961)
         );
  OAI22_X1 U2434 ( .A1(n1609), .A2(n1246), .B1(n1618), .B2(n1245), .ZN(n965)
         );
  OAI22_X1 U2435 ( .A1(n1854), .A2(n1248), .B1(n1695), .B2(n1247), .ZN(n967)
         );
  OAI22_X1 U2436 ( .A1(n1855), .A2(n1247), .B1(n1694), .B2(n1246), .ZN(n966)
         );
  OAI22_X1 U2437 ( .A1(n1249), .A2(n1855), .B1(n1617), .B2(n1248), .ZN(n968)
         );
  OAI22_X1 U2438 ( .A1(n1609), .A2(n1485), .B1(n1250), .B2(n1695), .ZN(n853)
         );
  NAND2_X1 U2439 ( .A1(n392), .A2(n364), .ZN(n151) );
  OAI22_X1 U2440 ( .A1(n1758), .A2(n1196), .B1(n1869), .B2(n1195), .ZN(n917)
         );
  OAI22_X1 U2441 ( .A1(n1758), .A2(n1198), .B1(n1869), .B2(n1197), .ZN(n919)
         );
  OAI22_X1 U2442 ( .A1(n1758), .A2(n1197), .B1(n1869), .B2(n1196), .ZN(n918)
         );
  OAI22_X1 U2443 ( .A1(n1709), .A2(n1199), .B1(n1869), .B2(n1198), .ZN(n920)
         );
  OAI22_X1 U2444 ( .A1(n1709), .A2(n1202), .B1(n1869), .B2(n1201), .ZN(n923)
         );
  OAI22_X1 U2445 ( .A1(n1710), .A2(n1200), .B1(n1869), .B2(n1199), .ZN(n921)
         );
  OAI22_X1 U2446 ( .A1(n1710), .A2(n1201), .B1(n1869), .B2(n1200), .ZN(n922)
         );
  OAI22_X1 U2447 ( .A1(n1710), .A2(n1205), .B1(n1869), .B2(n1204), .ZN(n926)
         );
  OAI22_X1 U2448 ( .A1(n1709), .A2(n1209), .B1(n1869), .B2(n1208), .ZN(n930)
         );
  OAI22_X1 U2449 ( .A1(n1710), .A2(n1203), .B1(n1869), .B2(n1202), .ZN(n924)
         );
  OAI22_X1 U2450 ( .A1(n1709), .A2(n1204), .B1(n1869), .B2(n1203), .ZN(n925)
         );
  AOI21_X1 U2451 ( .B1(n194), .B2(n338), .A(n191), .ZN(n189) );
  AOI21_X1 U2452 ( .B1(n194), .B2(n174), .A(n175), .ZN(n173) );
  AOI21_X1 U2453 ( .B1(n194), .B2(n1761), .A(n1759), .ZN(n180) );
  INV_X1 U2454 ( .A(n288), .ZN(n287) );
  OAI22_X1 U2455 ( .A1(n1769), .A2(n1356), .B1(n1699), .B2(n1355), .ZN(n1070)
         );
  OAI22_X1 U2456 ( .A1(n1908), .A2(n1357), .B1(n1699), .B2(n1356), .ZN(n1071)
         );
  OAI22_X1 U2457 ( .A1(n1908), .A2(n1358), .B1(n1753), .B2(n1357), .ZN(n1072)
         );
  OAI22_X1 U2458 ( .A1(n1907), .A2(n1359), .B1(n1699), .B2(n1358), .ZN(n1073)
         );
  OAI22_X1 U2459 ( .A1(n1908), .A2(n1360), .B1(n1753), .B2(n1359), .ZN(n1074)
         );
  OAI22_X1 U2460 ( .A1(n1769), .A2(n1362), .B1(n1910), .B2(n1361), .ZN(n1076)
         );
  OAI22_X1 U2461 ( .A1(n1907), .A2(n1364), .B1(n1753), .B2(n1363), .ZN(n1078)
         );
  OAI22_X1 U2462 ( .A1(n1907), .A2(n1363), .B1(n1753), .B2(n1362), .ZN(n1077)
         );
  NAND2_X1 U2463 ( .A1(n811), .A2(n1128), .ZN(n323) );
  OAI22_X1 U2464 ( .A1(n1907), .A2(n1376), .B1(n1678), .B2(n1375), .ZN(n1090)
         );
  OAI22_X1 U2465 ( .A1(n1908), .A2(n1713), .B1(n1385), .B2(n1753), .ZN(n858)
         );
  NAND2_X1 U2466 ( .A1(n15), .A2(n1465), .ZN(n18) );
  OAI22_X1 U2467 ( .A1(n1709), .A2(n1195), .B1(n1869), .B2(n1194), .ZN(n916)
         );
  OAI22_X1 U2468 ( .A1(n77), .A2(n1206), .B1(n1869), .B2(n1205), .ZN(n927) );
  OAI22_X1 U2469 ( .A1(n77), .A2(n1208), .B1(n1869), .B2(n1207), .ZN(n929) );
  OAI22_X1 U2470 ( .A1(n1709), .A2(n1207), .B1(n1869), .B2(n1206), .ZN(n928)
         );
  OAI22_X1 U2471 ( .A1(n1709), .A2(n1483), .B1(n1210), .B2(n1869), .ZN(n851)
         );
  XNOR2_X1 U2472 ( .A(n166), .B(n121), .ZN(product[29]) );
  NAND2_X1 U2473 ( .A1(n1700), .A2(n1879), .ZN(n127) );
  AOI21_X1 U2474 ( .B1(n166), .B2(n1831), .A(n163), .ZN(n161) );
  AOI21_X1 U2475 ( .B1(n166), .B2(n1830), .A(n154), .ZN(n152) );
  NAND2_X1 U2476 ( .A1(n216), .A2(n1700), .ZN(n205) );
  AOI21_X1 U2477 ( .B1(n217), .B2(n1700), .A(n1833), .ZN(n206) );
  NAND2_X1 U2478 ( .A1(n1834), .A2(n1832), .ZN(n198) );
  OAI22_X1 U2479 ( .A1(n1738), .A2(n1215), .B1(n1719), .B2(n1214), .ZN(n935)
         );
  OAI22_X1 U2480 ( .A1(n1814), .A2(n1214), .B1(n1719), .B2(n1213), .ZN(n934)
         );
  OAI22_X1 U2481 ( .A1(n1814), .A2(n1213), .B1(n1875), .B2(n1212), .ZN(n933)
         );
  XNOR2_X1 U2482 ( .A(n1859), .B(n1433), .ZN(n1232) );
  OAI22_X1 U2483 ( .A1(n1814), .A2(n1217), .B1(n1720), .B2(n1216), .ZN(n937)
         );
  XNOR2_X1 U2484 ( .A(n1858), .B(n1434), .ZN(n1233) );
  OAI22_X1 U2485 ( .A1(n1813), .A2(n1218), .B1(n1719), .B2(n1217), .ZN(n938)
         );
  OAI22_X1 U2486 ( .A1(n1738), .A2(n1216), .B1(n1719), .B2(n1215), .ZN(n936)
         );
  OAI22_X1 U2487 ( .A1(n1813), .A2(n1219), .B1(n1720), .B2(n1218), .ZN(n939)
         );
  OAI22_X1 U2488 ( .A1(n1814), .A2(n1220), .B1(n1719), .B2(n1219), .ZN(n940)
         );
  OAI22_X1 U2489 ( .A1(n1814), .A2(n1226), .B1(n1875), .B2(n1225), .ZN(n946)
         );
  OAI22_X1 U2490 ( .A1(n1813), .A2(n1227), .B1(n1719), .B2(n1226), .ZN(n947)
         );
  OAI22_X1 U2491 ( .A1(n1738), .A2(n1224), .B1(n1719), .B2(n1223), .ZN(n944)
         );
  OAI22_X1 U2492 ( .A1(n1738), .A2(n1212), .B1(n1719), .B2(n1211), .ZN(n932)
         );
  OAI22_X1 U2493 ( .A1(n1814), .A2(n1225), .B1(n1720), .B2(n1224), .ZN(n945)
         );
  OAI22_X1 U2494 ( .A1(n1813), .A2(n1221), .B1(n1719), .B2(n1220), .ZN(n941)
         );
  XNOR2_X1 U2495 ( .A(n1859), .B(n1435), .ZN(n1234) );
  OAI22_X1 U2496 ( .A1(n1738), .A2(n1484), .B1(n1229), .B2(n1720), .ZN(n852)
         );
  OAI22_X1 U2497 ( .A1(n1813), .A2(n1223), .B1(n1720), .B2(n1222), .ZN(n943)
         );
  OAI22_X1 U2498 ( .A1(n1813), .A2(n1228), .B1(n1719), .B2(n1227), .ZN(n948)
         );
  XNOR2_X1 U2499 ( .A(n1858), .B(n1436), .ZN(n1235) );
  OAI22_X1 U2500 ( .A1(n1738), .A2(n1222), .B1(n1720), .B2(n1221), .ZN(n942)
         );
  XNOR2_X1 U2501 ( .A(n1858), .B(n1439), .ZN(n1238) );
  XNOR2_X1 U2502 ( .A(n1859), .B(n1438), .ZN(n1237) );
  XNOR2_X1 U2503 ( .A(n1858), .B(n1437), .ZN(n1236) );
  XNOR2_X1 U2504 ( .A(n1858), .B(n1445), .ZN(n1244) );
  XNOR2_X1 U2505 ( .A(n1858), .B(n1431), .ZN(n1230) );
  XNOR2_X1 U2506 ( .A(n1858), .B(n1444), .ZN(n1243) );
  XNOR2_X1 U2507 ( .A(n1858), .B(n1432), .ZN(n1231) );
  XNOR2_X1 U2508 ( .A(n1858), .B(n1443), .ZN(n1242) );
  XNOR2_X1 U2509 ( .A(n1858), .B(n1442), .ZN(n1241) );
  XNOR2_X1 U2510 ( .A(n1859), .B(n1446), .ZN(n1245) );
  XNOR2_X1 U2511 ( .A(n1859), .B(n1440), .ZN(n1239) );
  XNOR2_X1 U2512 ( .A(n1859), .B(n1441), .ZN(n1240) );
  XNOR2_X1 U2513 ( .A(n1859), .B(n1917), .ZN(n1249) );
  XNOR2_X1 U2514 ( .A(n1859), .B(n1448), .ZN(n1247) );
  XNOR2_X1 U2515 ( .A(n1858), .B(n1447), .ZN(n1246) );
  XNOR2_X1 U2516 ( .A(n1859), .B(n1602), .ZN(n1248) );
  INV_X1 U2517 ( .A(n1858), .ZN(n1485) );
  XOR2_X1 U2518 ( .A(n55), .B(a[12]), .Z(n1460) );
  INV_X2 U2519 ( .A(n1934), .ZN(n1933) );
  INV_X1 U2520 ( .A(n50), .ZN(n1890) );
  CLKBUF_X3 U2521 ( .A(n116), .Z(n1917) );
  INV_X1 U2522 ( .A(n1919), .ZN(n1918) );
  INV_X1 U2523 ( .A(n3), .ZN(n1919) );
  INV_X1 U2524 ( .A(n3), .ZN(n1920) );
  INV_X1 U2525 ( .A(n1924), .ZN(n1921) );
  INV_X1 U2526 ( .A(n1924), .ZN(n1923) );
  INV_X1 U2527 ( .A(n21), .ZN(n1926) );
  INV_X1 U2528 ( .A(n21), .ZN(n1927) );
  INV_X1 U2529 ( .A(n30), .ZN(n1930) );
  INV_X1 U2530 ( .A(n30), .ZN(n1931) );
  INV_X1 U2531 ( .A(n1934), .ZN(n1932) );
  INV_X1 U2532 ( .A(n39), .ZN(n1934) );
  XOR2_X1 U2533 ( .A(n890), .B(n866), .Z(n389) );
  XOR2_X1 U2534 ( .A(n902), .B(n932), .Z(n387) );
  XOR2_X1 U2535 ( .A(n1100), .B(n1070), .Z(n383) );
  XOR2_X1 U2536 ( .A(n418), .B(n391), .Z(n377) );
  XOR2_X1 U2537 ( .A(n416), .B(n414), .Z(n375) );
  XOR2_X1 U2538 ( .A(n406), .B(n404), .Z(n369) );
  XOR2_X1 U2539 ( .A(n396), .B(n394), .Z(n363) );
endmodule


module datapath_M13_N16_T32_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n31,
         n32, n33, n35, n37, n38, n39, n40, n41, n43, n45, n46, n47, n48, n49,
         n51, n53, n54, n55, n56, n57, n59, n61, n62, n63, n64, n66, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n181, n182, n184, n186, n188, n191, n192, n193, n194, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n315, n316, n317, n318, n319, n320;

  FA_X1 U3 ( .A(B[30]), .B(A[30]), .CI(n32), .CO(n31), .S(SUM[30]) );
  FA_X1 U4 ( .A(B[29]), .B(A[29]), .CI(n182), .CO(n32), .S(SUM[29]) );
  NOR2_X1 U245 ( .A1(B[13]), .A2(A[13]), .ZN(n116) );
  NOR2_X1 U246 ( .A1(B[3]), .A2(A[3]), .ZN(n171) );
  AND2_X1 U247 ( .A1(n315), .A2(n181), .ZN(SUM[0]) );
  OR2_X1 U248 ( .A1(B[0]), .A2(A[0]), .ZN(n315) );
  NAND2_X1 U249 ( .A1(n139), .A2(n127), .ZN(n125) );
  AOI21_X1 U250 ( .B1(n79), .B2(n88), .A(n80), .ZN(n78) );
  AOI21_X1 U251 ( .B1(n127), .B2(n140), .A(n128), .ZN(n126) );
  NOR2_X1 U252 ( .A1(B[19]), .A2(A[19]), .ZN(n81) );
  NOR2_X1 U253 ( .A1(B[2]), .A2(A[2]), .ZN(n174) );
  NOR2_X1 U254 ( .A1(B[18]), .A2(A[18]), .ZN(n84) );
  NOR2_X1 U255 ( .A1(B[8]), .A2(A[8]), .ZN(n144) );
  NOR2_X1 U256 ( .A1(B[20]), .A2(A[20]), .ZN(n72) );
  NOR2_X1 U257 ( .A1(B[14]), .A2(A[14]), .ZN(n109) );
  NOR2_X1 U258 ( .A1(B[12]), .A2(A[12]), .ZN(n121) );
  NOR2_X1 U259 ( .A1(B[1]), .A2(A[1]), .ZN(n178) );
  NAND2_X1 U260 ( .A1(B[14]), .A2(A[14]), .ZN(n110) );
  NAND2_X1 U261 ( .A1(B[2]), .A2(A[2]), .ZN(n175) );
  NAND2_X1 U262 ( .A1(B[18]), .A2(A[18]), .ZN(n85) );
  NAND2_X1 U263 ( .A1(B[16]), .A2(A[16]), .ZN(n95) );
  NAND2_X1 U264 ( .A1(B[19]), .A2(A[19]), .ZN(n82) );
  OR2_X1 U265 ( .A1(B[21]), .A2(A[21]), .ZN(n316) );
  OR2_X1 U266 ( .A1(B[22]), .A2(A[22]), .ZN(n319) );
  INV_X1 U267 ( .A(n97), .ZN(n96) );
  INV_X1 U268 ( .A(n124), .ZN(n123) );
  INV_X1 U269 ( .A(n147), .ZN(n146) );
  AOI21_X1 U270 ( .B1(n96), .B2(n87), .A(n88), .ZN(n86) );
  AOI21_X1 U271 ( .B1(n167), .B2(n158), .A(n159), .ZN(n157) );
  AOI21_X1 U272 ( .B1(n147), .B2(n98), .A(n99), .ZN(n97) );
  NOR2_X1 U273 ( .A1(n125), .A2(n100), .ZN(n98) );
  OAI21_X1 U274 ( .B1(n126), .B2(n100), .A(n101), .ZN(n99) );
  NAND2_X1 U275 ( .A1(n114), .A2(n102), .ZN(n100) );
  OAI21_X1 U276 ( .B1(n123), .B2(n112), .A(n113), .ZN(n111) );
  INV_X1 U277 ( .A(n114), .ZN(n112) );
  INV_X1 U278 ( .A(n115), .ZN(n113) );
  OAI21_X1 U279 ( .B1(n146), .B2(n137), .A(n138), .ZN(n136) );
  INV_X1 U280 ( .A(n140), .ZN(n138) );
  INV_X1 U281 ( .A(n139), .ZN(n137) );
  INV_X1 U282 ( .A(n168), .ZN(n167) );
  OAI21_X1 U283 ( .B1(n146), .B2(n125), .A(n126), .ZN(n124) );
  AOI21_X1 U284 ( .B1(n96), .B2(n70), .A(n71), .ZN(n69) );
  AOI21_X1 U285 ( .B1(n96), .B2(n75), .A(n76), .ZN(n74) );
  INV_X1 U286 ( .A(n77), .ZN(n75) );
  INV_X1 U287 ( .A(n78), .ZN(n76) );
  INV_X1 U288 ( .A(n177), .ZN(n176) );
  NAND2_X1 U289 ( .A1(n87), .A2(n79), .ZN(n77) );
  AOI21_X1 U290 ( .B1(n46), .B2(n317), .A(n43), .ZN(n41) );
  INV_X1 U291 ( .A(n45), .ZN(n43) );
  AOI21_X1 U292 ( .B1(n62), .B2(n319), .A(n59), .ZN(n57) );
  INV_X1 U293 ( .A(n61), .ZN(n59) );
  AOI21_X1 U294 ( .B1(n54), .B2(n318), .A(n51), .ZN(n49) );
  INV_X1 U295 ( .A(n53), .ZN(n51) );
  OAI21_X1 U296 ( .B1(n89), .B2(n95), .A(n90), .ZN(n88) );
  OAI21_X1 U297 ( .B1(n160), .B2(n166), .A(n161), .ZN(n159) );
  OAI21_X1 U298 ( .B1(n78), .B2(n72), .A(n73), .ZN(n71) );
  OAI21_X1 U299 ( .B1(n81), .B2(n85), .A(n82), .ZN(n80) );
  AOI21_X1 U300 ( .B1(n169), .B2(n177), .A(n170), .ZN(n168) );
  NOR2_X1 U301 ( .A1(n174), .A2(n171), .ZN(n169) );
  OAI21_X1 U302 ( .B1(n171), .B2(n175), .A(n172), .ZN(n170) );
  OAI21_X1 U303 ( .B1(n41), .B2(n39), .A(n40), .ZN(n38) );
  OAI21_X1 U304 ( .B1(n49), .B2(n47), .A(n48), .ZN(n46) );
  OAI21_X1 U305 ( .B1(n57), .B2(n55), .A(n56), .ZN(n54) );
  NOR2_X1 U306 ( .A1(n77), .A2(n72), .ZN(n70) );
  NOR2_X1 U307 ( .A1(n94), .A2(n89), .ZN(n87) );
  NOR2_X1 U308 ( .A1(n165), .A2(n160), .ZN(n158) );
  OAI21_X1 U309 ( .B1(n178), .B2(n181), .A(n179), .ZN(n177) );
  OAI21_X1 U310 ( .B1(n116), .B2(n122), .A(n117), .ZN(n115) );
  NOR2_X1 U311 ( .A1(n84), .A2(n81), .ZN(n79) );
  NOR2_X1 U312 ( .A1(n109), .A2(n104), .ZN(n102) );
  OAI21_X1 U313 ( .B1(n168), .B2(n148), .A(n149), .ZN(n147) );
  NAND2_X1 U314 ( .A1(n158), .A2(n150), .ZN(n148) );
  AOI21_X1 U315 ( .B1(n150), .B2(n159), .A(n151), .ZN(n149) );
  NOR2_X1 U316 ( .A1(n155), .A2(n152), .ZN(n150) );
  AOI21_X1 U317 ( .B1(n102), .B2(n115), .A(n103), .ZN(n101) );
  OAI21_X1 U318 ( .B1(n104), .B2(n110), .A(n105), .ZN(n103) );
  OAI21_X1 U319 ( .B1(n97), .B2(n63), .A(n64), .ZN(n62) );
  NAND2_X1 U320 ( .A1(n70), .A2(n316), .ZN(n63) );
  AOI21_X1 U321 ( .B1(n71), .B2(n316), .A(n66), .ZN(n64) );
  INV_X1 U322 ( .A(n68), .ZN(n66) );
  AOI21_X1 U323 ( .B1(n96), .B2(n92), .A(n93), .ZN(n91) );
  INV_X1 U324 ( .A(n95), .ZN(n93) );
  AOI21_X1 U325 ( .B1(n111), .B2(n197), .A(n108), .ZN(n106) );
  INV_X1 U326 ( .A(n110), .ZN(n108) );
  AOI21_X1 U327 ( .B1(n124), .B2(n199), .A(n120), .ZN(n118) );
  INV_X1 U328 ( .A(n122), .ZN(n120) );
  AOI21_X1 U329 ( .B1(n167), .B2(n207), .A(n164), .ZN(n162) );
  INV_X1 U330 ( .A(n166), .ZN(n164) );
  AOI21_X1 U331 ( .B1(n136), .B2(n201), .A(n133), .ZN(n131) );
  INV_X1 U332 ( .A(n135), .ZN(n133) );
  NOR2_X1 U333 ( .A1(n121), .A2(n116), .ZN(n114) );
  OAI21_X1 U334 ( .B1(n152), .B2(n156), .A(n153), .ZN(n151) );
  INV_X1 U335 ( .A(n94), .ZN(n92) );
  INV_X1 U336 ( .A(n121), .ZN(n199) );
  INV_X1 U337 ( .A(n165), .ZN(n207) );
  INV_X1 U338 ( .A(n109), .ZN(n197) );
  INV_X1 U339 ( .A(n134), .ZN(n201) );
  NAND2_X1 U340 ( .A1(n200), .A2(n130), .ZN(n19) );
  OAI21_X1 U341 ( .B1(n86), .B2(n84), .A(n85), .ZN(n83) );
  OAI21_X1 U342 ( .B1(n146), .B2(n144), .A(n145), .ZN(n143) );
  OAI21_X1 U343 ( .B1(n157), .B2(n155), .A(n156), .ZN(n154) );
  OAI21_X1 U344 ( .B1(n176), .B2(n174), .A(n175), .ZN(n173) );
  NAND2_X1 U345 ( .A1(n208), .A2(n172), .ZN(n27) );
  INV_X1 U346 ( .A(n171), .ZN(n208) );
  NAND2_X1 U347 ( .A1(n196), .A2(n105), .ZN(n15) );
  INV_X1 U348 ( .A(n104), .ZN(n196) );
  NAND2_X1 U349 ( .A1(n198), .A2(n117), .ZN(n17) );
  INV_X1 U350 ( .A(n116), .ZN(n198) );
  NAND2_X1 U351 ( .A1(n191), .A2(n73), .ZN(n10) );
  INV_X1 U352 ( .A(n72), .ZN(n191) );
  NAND2_X1 U353 ( .A1(n193), .A2(n85), .ZN(n12) );
  INV_X1 U354 ( .A(n84), .ZN(n193) );
  NAND2_X1 U355 ( .A1(n205), .A2(n156), .ZN(n24) );
  INV_X1 U356 ( .A(n155), .ZN(n205) );
  NAND2_X1 U357 ( .A1(n192), .A2(n82), .ZN(n11) );
  INV_X1 U358 ( .A(n81), .ZN(n192) );
  NAND2_X1 U359 ( .A1(n194), .A2(n90), .ZN(n13) );
  INV_X1 U360 ( .A(n89), .ZN(n194) );
  NAND2_X1 U361 ( .A1(n206), .A2(n161), .ZN(n25) );
  INV_X1 U362 ( .A(n160), .ZN(n206) );
  NAND2_X1 U363 ( .A1(n203), .A2(n145), .ZN(n22) );
  INV_X1 U364 ( .A(n144), .ZN(n203) );
  NAND2_X1 U365 ( .A1(n210), .A2(n179), .ZN(n29) );
  INV_X1 U366 ( .A(n178), .ZN(n210) );
  NAND2_X1 U367 ( .A1(n320), .A2(n37), .ZN(n2) );
  NAND2_X1 U368 ( .A1(n202), .A2(n142), .ZN(n21) );
  NAND2_X1 U369 ( .A1(n92), .A2(n95), .ZN(n14) );
  NAND2_X1 U370 ( .A1(n207), .A2(n166), .ZN(n26) );
  NAND2_X1 U371 ( .A1(n197), .A2(n110), .ZN(n16) );
  NAND2_X1 U372 ( .A1(n209), .A2(n175), .ZN(n28) );
  INV_X1 U373 ( .A(n174), .ZN(n209) );
  NAND2_X1 U374 ( .A1(n199), .A2(n122), .ZN(n18) );
  NAND2_X1 U375 ( .A1(n204), .A2(n153), .ZN(n23) );
  INV_X1 U376 ( .A(n152), .ZN(n204) );
  NAND2_X1 U377 ( .A1(n201), .A2(n135), .ZN(n20) );
  NAND2_X1 U378 ( .A1(n316), .A2(n68), .ZN(n9) );
  NAND2_X1 U379 ( .A1(n317), .A2(n45), .ZN(n4) );
  NAND2_X1 U380 ( .A1(n318), .A2(n53), .ZN(n6) );
  NAND2_X1 U381 ( .A1(n319), .A2(n61), .ZN(n8) );
  NAND2_X1 U382 ( .A1(n184), .A2(n40), .ZN(n3) );
  INV_X1 U383 ( .A(n39), .ZN(n184) );
  NAND2_X1 U384 ( .A1(n186), .A2(n48), .ZN(n5) );
  INV_X1 U385 ( .A(n47), .ZN(n186) );
  NAND2_X1 U386 ( .A1(n188), .A2(n56), .ZN(n7) );
  INV_X1 U387 ( .A(n55), .ZN(n188) );
  NOR2_X1 U388 ( .A1(B[6]), .A2(A[6]), .ZN(n155) );
  NOR2_X2 U389 ( .A1(B[17]), .A2(A[17]), .ZN(n89) );
  NOR2_X1 U390 ( .A1(B[5]), .A2(A[5]), .ZN(n160) );
  NOR2_X1 U391 ( .A1(B[7]), .A2(A[7]), .ZN(n152) );
  XOR2_X1 U392 ( .A(A[31]), .B(B[31]), .Z(n1) );
  NOR2_X1 U393 ( .A1(B[4]), .A2(A[4]), .ZN(n165) );
  NOR2_X1 U394 ( .A1(B[16]), .A2(A[16]), .ZN(n94) );
  NOR2_X1 U395 ( .A1(B[25]), .A2(A[25]), .ZN(n47) );
  NOR2_X1 U396 ( .A1(B[23]), .A2(A[23]), .ZN(n55) );
  NOR2_X1 U397 ( .A1(B[27]), .A2(A[27]), .ZN(n39) );
  XOR2_X1 U398 ( .A(n41), .B(n3), .Z(SUM[27]) );
  OR2_X1 U399 ( .A1(B[26]), .A2(A[26]), .ZN(n317) );
  OR2_X1 U400 ( .A1(B[24]), .A2(A[24]), .ZN(n318) );
  OR2_X1 U401 ( .A1(B[28]), .A2(A[28]), .ZN(n320) );
  NAND2_X1 U402 ( .A1(B[6]), .A2(A[6]), .ZN(n156) );
  NAND2_X1 U403 ( .A1(B[0]), .A2(A[0]), .ZN(n181) );
  NAND2_X1 U404 ( .A1(B[4]), .A2(A[4]), .ZN(n166) );
  NAND2_X1 U405 ( .A1(B[12]), .A2(A[12]), .ZN(n122) );
  NAND2_X1 U406 ( .A1(B[8]), .A2(A[8]), .ZN(n145) );
  INV_X1 U407 ( .A(n33), .ZN(n182) );
  AOI21_X1 U408 ( .B1(n38), .B2(n320), .A(n35), .ZN(n33) );
  INV_X1 U409 ( .A(n37), .ZN(n35) );
  NAND2_X1 U410 ( .A1(B[7]), .A2(A[7]), .ZN(n153) );
  NAND2_X1 U411 ( .A1(B[17]), .A2(A[17]), .ZN(n90) );
  NAND2_X1 U412 ( .A1(B[25]), .A2(A[25]), .ZN(n48) );
  NAND2_X1 U413 ( .A1(B[20]), .A2(A[20]), .ZN(n73) );
  NAND2_X1 U414 ( .A1(B[5]), .A2(A[5]), .ZN(n161) );
  NAND2_X1 U415 ( .A1(B[23]), .A2(A[23]), .ZN(n56) );
  NAND2_X1 U416 ( .A1(B[27]), .A2(A[27]), .ZN(n40) );
  NAND2_X1 U417 ( .A1(B[1]), .A2(A[1]), .ZN(n179) );
  NOR2_X1 U418 ( .A1(B[10]), .A2(A[10]), .ZN(n134) );
  NAND2_X1 U419 ( .A1(B[10]), .A2(A[10]), .ZN(n135) );
  NAND2_X1 U420 ( .A1(B[26]), .A2(A[26]), .ZN(n45) );
  NAND2_X1 U421 ( .A1(B[24]), .A2(A[24]), .ZN(n53) );
  NAND2_X1 U422 ( .A1(B[21]), .A2(A[21]), .ZN(n68) );
  NAND2_X1 U423 ( .A1(B[22]), .A2(A[22]), .ZN(n61) );
  XNOR2_X1 U424 ( .A(n54), .B(n6), .ZN(SUM[24]) );
  XOR2_X1 U425 ( .A(n57), .B(n7), .Z(SUM[23]) );
  XOR2_X1 U426 ( .A(n69), .B(n9), .Z(SUM[21]) );
  XOR2_X1 U427 ( .A(n74), .B(n10), .Z(SUM[20]) );
  XNOR2_X1 U428 ( .A(n83), .B(n11), .ZN(SUM[19]) );
  XOR2_X1 U429 ( .A(n86), .B(n12), .Z(SUM[18]) );
  XOR2_X1 U430 ( .A(n91), .B(n13), .Z(SUM[17]) );
  XOR2_X1 U431 ( .A(n106), .B(n15), .Z(SUM[15]) );
  XNOR2_X1 U432 ( .A(n111), .B(n16), .ZN(SUM[14]) );
  XOR2_X1 U433 ( .A(n118), .B(n17), .Z(SUM[13]) );
  XOR2_X1 U434 ( .A(n123), .B(n18), .Z(SUM[12]) );
  XOR2_X1 U435 ( .A(n131), .B(n19), .Z(SUM[11]) );
  XNOR2_X1 U436 ( .A(n38), .B(n2), .ZN(SUM[28]) );
  XNOR2_X1 U437 ( .A(n46), .B(n4), .ZN(SUM[26]) );
  XOR2_X1 U438 ( .A(n49), .B(n5), .Z(SUM[25]) );
  XNOR2_X1 U439 ( .A(n62), .B(n8), .ZN(SUM[22]) );
  XNOR2_X1 U440 ( .A(n96), .B(n14), .ZN(SUM[16]) );
  XNOR2_X1 U441 ( .A(n136), .B(n20), .ZN(SUM[10]) );
  XNOR2_X1 U442 ( .A(n143), .B(n21), .ZN(SUM[9]) );
  XOR2_X1 U443 ( .A(n146), .B(n22), .Z(SUM[8]) );
  XNOR2_X1 U444 ( .A(n154), .B(n23), .ZN(SUM[7]) );
  XOR2_X1 U445 ( .A(n157), .B(n24), .Z(SUM[6]) );
  XOR2_X1 U446 ( .A(n162), .B(n25), .Z(SUM[5]) );
  XNOR2_X1 U447 ( .A(n167), .B(n26), .ZN(SUM[4]) );
  XNOR2_X1 U448 ( .A(n173), .B(n27), .ZN(SUM[3]) );
  XOR2_X1 U449 ( .A(n176), .B(n28), .Z(SUM[2]) );
  XOR2_X1 U450 ( .A(n29), .B(n181), .Z(SUM[1]) );
  NAND2_X1 U451 ( .A1(B[28]), .A2(A[28]), .ZN(n37) );
  NAND2_X1 U452 ( .A1(B[13]), .A2(A[13]), .ZN(n117) );
  NAND2_X1 U453 ( .A1(B[15]), .A2(A[15]), .ZN(n105) );
  NOR2_X2 U454 ( .A1(B[15]), .A2(A[15]), .ZN(n104) );
  NAND2_X1 U455 ( .A1(B[3]), .A2(A[3]), .ZN(n172) );
  OAI21_X1 U456 ( .B1(n141), .B2(n145), .A(n142), .ZN(n140) );
  NOR2_X1 U457 ( .A1(n144), .A2(n141), .ZN(n139) );
  INV_X1 U458 ( .A(n141), .ZN(n202) );
  NOR2_X1 U459 ( .A1(B[9]), .A2(A[9]), .ZN(n141) );
  OAI21_X1 U460 ( .B1(n129), .B2(n135), .A(n130), .ZN(n128) );
  NOR2_X1 U461 ( .A1(n134), .A2(n129), .ZN(n127) );
  INV_X1 U462 ( .A(n129), .ZN(n200) );
  NOR2_X1 U463 ( .A1(B[11]), .A2(A[11]), .ZN(n129) );
  NAND2_X1 U464 ( .A1(B[9]), .A2(A[9]), .ZN(n142) );
  NAND2_X1 U465 ( .A1(B[11]), .A2(A[11]), .ZN(n130) );
  XOR2_X1 U466 ( .A(n31), .B(n1), .Z(SUM[31]) );
endmodule


module datapath_M13_N16_T32 ( clk, clear_acc, data_in, data_out, wr_en_x, 
        wr_en_y, addr_x, addr_w, addr_b, m_valid, m_ready );
  input [31:0] data_in;
  output [31:0] data_out;
  input [4:0] addr_x;
  input [7:0] addr_w;
  input [3:0] addr_b;
  input clk, clear_acc, wr_en_x, wr_en_y, m_valid, m_ready;
  wire   delay, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53,
         N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67,
         N68, N69, N70, N71, N72, N73, n111, n112, n113, n114, n117, n118,
         n119, n120, n121, n122, n123, n124, n128, n129, n130, n131, n133,
         n144, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n1, n2, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n115, n116, n125, n126,
         n127, n132, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n145, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289;
  wire   [31:0] data_out_x;
  wire   [31:0] data_out_w;
  wire   [31:0] data_out_b;
  wire   [31:0] f;
  wire   [31:0] adder;
  wire   [31:0] mul_out;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31;

  DFF_X1 more_delay_reg ( .D(delay), .CK(clk), .QN(n111) );
  DFF_X1 \mul_out_reg[31]  ( .D(n177), .CK(clk), .Q(n15) );
  DFF_X1 \mul_out_reg[30]  ( .D(n176), .CK(clk), .Q(n16) );
  DFF_X1 \mul_out_reg[29]  ( .D(n175), .CK(clk), .Q(n17) );
  DFF_X1 \mul_out_reg[26]  ( .D(n172), .CK(clk), .Q(n20) );
  DFF_X1 \mul_out_reg[25]  ( .D(n171), .CK(clk), .Q(n21) );
  DFF_X1 \mul_out_reg[24]  ( .D(n170), .CK(clk), .Q(n22) );
  DFF_X1 \mul_out_reg[23]  ( .D(n169), .CK(clk), .Q(n23) );
  DFF_X1 \mul_out_reg[22]  ( .D(n168), .CK(clk), .Q(mul_out[22]) );
  DFF_X1 \mul_out_reg[21]  ( .D(n167), .CK(clk), .Q(mul_out[21]) );
  DFF_X1 \mul_out_reg[20]  ( .D(n166), .CK(clk), .Q(mul_out[20]), .QN(n133) );
  DFF_X1 \mul_out_reg[19]  ( .D(n165), .CK(clk), .Q(mul_out[19]) );
  DFF_X1 \mul_out_reg[18]  ( .D(n164), .CK(clk), .Q(mul_out[18]), .QN(n131) );
  DFF_X1 \mul_out_reg[17]  ( .D(n163), .CK(clk), .Q(mul_out[17]), .QN(n130) );
  DFF_X1 \mul_out_reg[16]  ( .D(n162), .CK(clk), .Q(mul_out[16]), .QN(n129) );
  DFF_X1 \mul_out_reg[15]  ( .D(n161), .CK(clk), .Q(mul_out[15]), .QN(n128) );
  DFF_X1 \mul_out_reg[12]  ( .D(n158), .CK(clk), .Q(mul_out[12]) );
  DFF_X1 \mul_out_reg[11]  ( .D(n157), .CK(clk), .Q(mul_out[11]), .QN(n124) );
  DFF_X1 \mul_out_reg[10]  ( .D(n156), .CK(clk), .Q(mul_out[10]), .QN(n123) );
  DFF_X1 \mul_out_reg[9]  ( .D(n155), .CK(clk), .Q(mul_out[9]), .QN(n122) );
  DFF_X1 \mul_out_reg[8]  ( .D(n154), .CK(clk), .Q(mul_out[8]), .QN(n121) );
  DFF_X1 \mul_out_reg[7]  ( .D(n153), .CK(clk), .Q(mul_out[7]), .QN(n120) );
  DFF_X1 \mul_out_reg[6]  ( .D(n152), .CK(clk), .Q(mul_out[6]), .QN(n119) );
  DFF_X1 \mul_out_reg[5]  ( .D(n151), .CK(clk), .Q(mul_out[5]), .QN(n118) );
  DFF_X1 \mul_out_reg[4]  ( .D(n150), .CK(clk), .Q(mul_out[4]), .QN(n117) );
  DFF_X1 \mul_out_reg[2]  ( .D(n148), .CK(clk), .Q(mul_out[2]) );
  DFF_X1 \mul_out_reg[1]  ( .D(n147), .CK(clk), .Q(mul_out[1]), .QN(n114) );
  DFF_X1 \mul_out_reg[0]  ( .D(n146), .CK(clk), .Q(mul_out[0]), .QN(n113) );
  DFF_X1 \f_reg[0]  ( .D(n289), .CK(clk), .Q(f[0]), .QN(n209) );
  DFF_X1 \f_reg[1]  ( .D(n288), .CK(clk), .Q(f[1]), .QN(n208) );
  DFF_X1 \f_reg[2]  ( .D(n287), .CK(clk), .Q(f[2]), .QN(n207) );
  DFF_X1 \f_reg[3]  ( .D(n286), .CK(clk), .Q(f[3]), .QN(n206) );
  DFF_X1 \f_reg[4]  ( .D(n285), .CK(clk), .Q(f[4]), .QN(n205) );
  DFF_X1 \f_reg[5]  ( .D(n284), .CK(clk), .Q(f[5]), .QN(n204) );
  DFF_X1 \f_reg[6]  ( .D(n283), .CK(clk), .Q(f[6]), .QN(n203) );
  DFF_X1 \f_reg[7]  ( .D(n282), .CK(clk), .Q(f[7]), .QN(n202) );
  DFF_X1 \f_reg[8]  ( .D(n281), .CK(clk), .Q(f[8]), .QN(n201) );
  DFF_X1 \f_reg[10]  ( .D(n279), .CK(clk), .Q(f[10]), .QN(n199) );
  DFF_X1 \f_reg[11]  ( .D(n278), .CK(clk), .Q(f[11]), .QN(n198) );
  DFF_X1 \f_reg[12]  ( .D(n277), .CK(clk), .Q(f[12]), .QN(n197) );
  DFF_X1 \f_reg[13]  ( .D(n276), .CK(clk), .Q(f[13]), .QN(n196) );
  DFF_X1 \f_reg[14]  ( .D(n275), .CK(clk), .Q(f[14]), .QN(n195) );
  DFF_X1 \f_reg[15]  ( .D(n274), .CK(clk), .Q(f[15]), .QN(n194) );
  DFF_X1 \f_reg[16]  ( .D(n188), .CK(clk), .Q(f[16]), .QN(n193) );
  DFF_X1 \f_reg[17]  ( .D(n187), .CK(clk), .Q(f[17]), .QN(n192) );
  DFF_X1 \f_reg[18]  ( .D(n186), .CK(clk), .Q(f[18]), .QN(n191) );
  DFF_X1 \f_reg[19]  ( .D(n185), .CK(clk), .Q(f[19]), .QN(n190) );
  DFF_X1 \f_reg[20]  ( .D(n184), .CK(clk), .Q(f[20]), .QN(n189) );
  DFF_X1 \f_reg[31]  ( .D(n140), .CK(clk), .Q(f[31]), .QN(n134) );
  memory_WIDTH32_SIZE16_LOGSIZE5 mem_x ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_x), .addr(addr_x), .wr_en(wr_en_x) );
  layer_13_16_1_32_W_rom mem_w ( .clk(clk), .addr(addr_w), .z(data_out_w) );
  layer_13_16_1_32_B_rom mem_b ( .clk(clk), .addr(addr_b), .z(data_out_b) );
  datapath_M13_N16_T32_DW_mult_tc_1 mult_101 ( .a(data_out_x), .b(data_out_w), 
        .product({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, N73, N72, N71, N70, 
        N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, 
        N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42})
         );
  datapath_M13_N16_T32_DW01_add_1 add_105 ( .A({n15, n16, n17, n18, n19, n20, 
        n21, n22, n23, mul_out[22:15], n29, n30, mul_out[12:4], n39, 
        mul_out[2:0]}), .B(f), .CI(1'b0), .SUM(adder) );
  DFF_X1 \mul_out_reg[28]  ( .D(n174), .CK(clk), .Q(n18) );
  DFF_X1 clear_acc_delay_reg ( .D(clear_acc), .CK(clk), .Q(n96), .QN(n112) );
  DFF_X1 delay_reg ( .D(n139), .CK(clk), .Q(delay), .QN(n144) );
  DFF_X1 \data_out_reg[31]  ( .D(n273), .CK(clk), .Q(data_out[31]), .QN(n210)
         );
  DFF_X1 \data_out_reg[30]  ( .D(n272), .CK(clk), .Q(data_out[30]), .QN(n211)
         );
  DFF_X1 \data_out_reg[29]  ( .D(n271), .CK(clk), .Q(data_out[29]), .QN(n212)
         );
  DFF_X1 \data_out_reg[28]  ( .D(n270), .CK(clk), .Q(data_out[28]), .QN(n213)
         );
  DFF_X1 \data_out_reg[27]  ( .D(n269), .CK(clk), .Q(data_out[27]), .QN(n214)
         );
  DFF_X1 \data_out_reg[26]  ( .D(n268), .CK(clk), .Q(data_out[26]), .QN(n215)
         );
  DFF_X1 \data_out_reg[25]  ( .D(n267), .CK(clk), .Q(data_out[25]), .QN(n216)
         );
  DFF_X1 \data_out_reg[24]  ( .D(n266), .CK(clk), .Q(data_out[24]), .QN(n217)
         );
  DFF_X1 \data_out_reg[23]  ( .D(n265), .CK(clk), .Q(data_out[23]), .QN(n218)
         );
  DFF_X1 \data_out_reg[22]  ( .D(n264), .CK(clk), .Q(data_out[22]), .QN(n219)
         );
  DFF_X1 \data_out_reg[21]  ( .D(n263), .CK(clk), .Q(data_out[21]), .QN(n220)
         );
  DFF_X1 \data_out_reg[20]  ( .D(n262), .CK(clk), .Q(data_out[20]), .QN(n221)
         );
  DFF_X1 \data_out_reg[19]  ( .D(n261), .CK(clk), .Q(data_out[19]), .QN(n222)
         );
  DFF_X1 \data_out_reg[18]  ( .D(n260), .CK(clk), .Q(data_out[18]), .QN(n223)
         );
  DFF_X1 \data_out_reg[17]  ( .D(n259), .CK(clk), .Q(data_out[17]), .QN(n224)
         );
  DFF_X1 \data_out_reg[16]  ( .D(n258), .CK(clk), .Q(data_out[16]), .QN(n225)
         );
  DFF_X1 \data_out_reg[15]  ( .D(n257), .CK(clk), .Q(data_out[15]), .QN(n226)
         );
  DFF_X1 \data_out_reg[14]  ( .D(n256), .CK(clk), .Q(data_out[14]), .QN(n227)
         );
  DFF_X1 \data_out_reg[13]  ( .D(n255), .CK(clk), .Q(data_out[13]), .QN(n228)
         );
  DFF_X1 \data_out_reg[12]  ( .D(n254), .CK(clk), .Q(data_out[12]), .QN(n229)
         );
  DFF_X1 \data_out_reg[11]  ( .D(n253), .CK(clk), .Q(data_out[11]), .QN(n230)
         );
  DFF_X1 \data_out_reg[10]  ( .D(n252), .CK(clk), .Q(data_out[10]), .QN(n231)
         );
  DFF_X1 \data_out_reg[9]  ( .D(n251), .CK(clk), .Q(data_out[9]), .QN(n232) );
  DFF_X1 \data_out_reg[8]  ( .D(n250), .CK(clk), .Q(data_out[8]), .QN(n233) );
  DFF_X1 \data_out_reg[7]  ( .D(n249), .CK(clk), .Q(data_out[7]), .QN(n234) );
  DFF_X1 \data_out_reg[6]  ( .D(n248), .CK(clk), .Q(data_out[6]), .QN(n235) );
  DFF_X1 \data_out_reg[5]  ( .D(n247), .CK(clk), .Q(data_out[5]), .QN(n236) );
  DFF_X1 \data_out_reg[4]  ( .D(n246), .CK(clk), .Q(data_out[4]), .QN(n237) );
  DFF_X1 \data_out_reg[3]  ( .D(n245), .CK(clk), .Q(data_out[3]), .QN(n238) );
  DFF_X1 \data_out_reg[2]  ( .D(n244), .CK(clk), .Q(data_out[2]), .QN(n239) );
  DFF_X1 \data_out_reg[1]  ( .D(n243), .CK(clk), .Q(data_out[1]), .QN(n240) );
  DFF_X1 \data_out_reg[0]  ( .D(n242), .CK(clk), .Q(data_out[0]), .QN(n241) );
  DFF_X1 \f_reg[22]  ( .D(n182), .CK(clk), .Q(f[22]), .QN(n100) );
  DFF_X1 \f_reg[23]  ( .D(n181), .CK(clk), .Q(f[23]), .QN(n101) );
  DFF_X1 \f_reg[24]  ( .D(n180), .CK(clk), .Q(f[24]), .QN(n102) );
  DFF_X1 \f_reg[25]  ( .D(n179), .CK(clk), .Q(f[25]), .QN(n103) );
  DFF_X1 \f_reg[26]  ( .D(n178), .CK(clk), .Q(f[26]), .QN(n104) );
  DFF_X1 \f_reg[27]  ( .D(n145), .CK(clk), .Q(f[27]), .QN(n105) );
  DFF_X1 \f_reg[28]  ( .D(n143), .CK(clk), .Q(f[28]), .QN(n106) );
  DFF_X1 \f_reg[21]  ( .D(n183), .CK(clk), .Q(f[21]), .QN(n99) );
  DFF_X1 \f_reg[29]  ( .D(n142), .CK(clk), .Q(f[29]), .QN(n107) );
  DFF_X1 \f_reg[30]  ( .D(n141), .CK(clk), .Q(f[30]), .QN(n108) );
  DFF_X1 \mul_out_reg[14]  ( .D(n160), .CK(clk), .Q(n29) );
  DFF_X1 \mul_out_reg[13]  ( .D(n159), .CK(clk), .Q(n30) );
  DFF_X1 \mul_out_reg[3]  ( .D(n149), .CK(clk), .Q(n39) );
  DFF_X1 \f_reg[9]  ( .D(n280), .CK(clk), .Q(f[9]), .QN(n200) );
  DFF_X1 \mul_out_reg[27]  ( .D(n173), .CK(clk), .Q(n19) );
  NAND2_X1 U3 ( .A1(N66), .A2(n1), .ZN(n2) );
  NAND2_X1 U4 ( .A1(n22), .A2(delay), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n2), .A2(n4), .ZN(n170) );
  INV_X2 U7 ( .A(delay), .ZN(n1) );
  MUX2_X1 U8 ( .A(N67), .B(n21), .S(delay), .Z(n171) );
  MUX2_X1 U9 ( .A(N64), .B(mul_out[22]), .S(delay), .Z(n168) );
  MUX2_X1 U10 ( .A(N65), .B(n23), .S(delay), .Z(n169) );
  MUX2_X1 U11 ( .A(N71), .B(n17), .S(delay), .Z(n175) );
  MUX2_X1 U12 ( .A(N69), .B(n19), .S(delay), .Z(n173) );
  MUX2_X1 U13 ( .A(N70), .B(n18), .S(delay), .Z(n174) );
  MUX2_X1 U14 ( .A(N68), .B(n20), .S(delay), .Z(n172) );
  MUX2_X1 U15 ( .A(N73), .B(n15), .S(delay), .Z(n177) );
  MUX2_X1 U16 ( .A(N72), .B(n16), .S(delay), .Z(n176) );
  AND2_X1 U17 ( .A1(n112), .A2(n44), .ZN(n5) );
  BUF_X1 U18 ( .A(n95), .Z(n6) );
  BUF_X1 U19 ( .A(n5), .Z(n7) );
  BUF_X1 U20 ( .A(n137), .Z(n9) );
  BUF_X1 U21 ( .A(n138), .Z(n10) );
  BUF_X1 U22 ( .A(n96), .Z(n8) );
  BUF_X1 U23 ( .A(n144), .Z(n12) );
  BUF_X1 U24 ( .A(n144), .Z(n11) );
  BUF_X1 U25 ( .A(n144), .Z(n13) );
  INV_X1 U26 ( .A(m_ready), .ZN(n14) );
  NAND2_X1 U27 ( .A1(m_valid), .A2(n14), .ZN(n42) );
  INV_X1 U28 ( .A(n42), .ZN(n139) );
  MUX2_X1 U29 ( .A(mul_out[21]), .B(N63), .S(n11), .Z(n167) );
  INV_X1 U30 ( .A(n133), .ZN(n24) );
  MUX2_X1 U31 ( .A(n24), .B(N62), .S(n11), .Z(n166) );
  MUX2_X1 U32 ( .A(mul_out[19]), .B(N61), .S(n12), .Z(n165) );
  INV_X1 U33 ( .A(n131), .ZN(n25) );
  MUX2_X1 U34 ( .A(n25), .B(N60), .S(n12), .Z(n164) );
  INV_X1 U35 ( .A(n130), .ZN(n26) );
  MUX2_X1 U36 ( .A(n26), .B(N59), .S(n12), .Z(n163) );
  INV_X1 U37 ( .A(n129), .ZN(n27) );
  MUX2_X1 U38 ( .A(n27), .B(N58), .S(n12), .Z(n162) );
  INV_X1 U39 ( .A(n128), .ZN(n28) );
  MUX2_X1 U40 ( .A(n28), .B(N57), .S(n12), .Z(n161) );
  MUX2_X1 U41 ( .A(n29), .B(N56), .S(n12), .Z(n160) );
  MUX2_X1 U42 ( .A(n30), .B(N55), .S(n12), .Z(n159) );
  MUX2_X1 U43 ( .A(mul_out[12]), .B(N54), .S(n12), .Z(n158) );
  INV_X1 U44 ( .A(n124), .ZN(n31) );
  MUX2_X1 U45 ( .A(n31), .B(N53), .S(n12), .Z(n157) );
  INV_X1 U46 ( .A(n123), .ZN(n32) );
  MUX2_X1 U47 ( .A(n32), .B(N52), .S(n12), .Z(n156) );
  INV_X1 U48 ( .A(n122), .ZN(n33) );
  MUX2_X1 U49 ( .A(n33), .B(N51), .S(n12), .Z(n155) );
  INV_X1 U50 ( .A(n121), .ZN(n34) );
  MUX2_X1 U51 ( .A(n34), .B(N50), .S(n12), .Z(n154) );
  INV_X1 U52 ( .A(n120), .ZN(n35) );
  MUX2_X1 U53 ( .A(n35), .B(N49), .S(n13), .Z(n153) );
  INV_X1 U54 ( .A(n119), .ZN(n36) );
  MUX2_X1 U55 ( .A(n36), .B(N48), .S(n13), .Z(n152) );
  INV_X1 U56 ( .A(n118), .ZN(n37) );
  MUX2_X1 U57 ( .A(n37), .B(N47), .S(n13), .Z(n151) );
  INV_X1 U58 ( .A(n117), .ZN(n38) );
  MUX2_X1 U59 ( .A(n38), .B(N46), .S(n13), .Z(n150) );
  MUX2_X1 U60 ( .A(n39), .B(N45), .S(n13), .Z(n149) );
  MUX2_X1 U61 ( .A(mul_out[2]), .B(N44), .S(n13), .Z(n148) );
  INV_X1 U62 ( .A(n114), .ZN(n40) );
  MUX2_X1 U63 ( .A(n40), .B(N43), .S(n13), .Z(n147) );
  INV_X1 U64 ( .A(n113), .ZN(n41) );
  MUX2_X1 U65 ( .A(n41), .B(N42), .S(n13), .Z(n146) );
  NAND3_X1 U66 ( .A1(n111), .A2(n13), .A3(n42), .ZN(n43) );
  NAND2_X1 U67 ( .A1(n112), .A2(n43), .ZN(n44) );
  INV_X1 U68 ( .A(n44), .ZN(n95) );
  AOI222_X1 U69 ( .A1(data_out_b[31]), .A2(n96), .B1(adder[31]), .B2(n5), .C1(
        n6), .C2(f[31]), .ZN(n45) );
  INV_X1 U70 ( .A(n45), .ZN(n140) );
  AOI222_X1 U71 ( .A1(data_out_b[29]), .A2(n96), .B1(adder[29]), .B2(n5), .C1(
        n6), .C2(f[29]), .ZN(n46) );
  INV_X1 U72 ( .A(n46), .ZN(n142) );
  AOI222_X1 U73 ( .A1(data_out_b[28]), .A2(n96), .B1(adder[28]), .B2(n5), .C1(
        n6), .C2(f[28]), .ZN(n47) );
  INV_X1 U74 ( .A(n47), .ZN(n143) );
  AOI222_X1 U75 ( .A1(data_out_b[27]), .A2(n96), .B1(adder[27]), .B2(n5), .C1(
        n6), .C2(f[27]), .ZN(n48) );
  INV_X1 U76 ( .A(n48), .ZN(n145) );
  AOI222_X1 U77 ( .A1(data_out_b[26]), .A2(n96), .B1(adder[26]), .B2(n5), .C1(
        n6), .C2(f[26]), .ZN(n49) );
  INV_X1 U78 ( .A(n49), .ZN(n178) );
  AOI222_X1 U79 ( .A1(data_out_b[25]), .A2(n96), .B1(adder[25]), .B2(n5), .C1(
        n6), .C2(f[25]), .ZN(n50) );
  INV_X1 U80 ( .A(n50), .ZN(n179) );
  AOI222_X1 U81 ( .A1(data_out_b[24]), .A2(n96), .B1(adder[24]), .B2(n5), .C1(
        n6), .C2(f[24]), .ZN(n51) );
  INV_X1 U82 ( .A(n51), .ZN(n180) );
  AOI222_X1 U83 ( .A1(data_out_b[23]), .A2(n96), .B1(adder[23]), .B2(n5), .C1(
        n6), .C2(f[23]), .ZN(n52) );
  INV_X1 U84 ( .A(n52), .ZN(n181) );
  AOI222_X1 U85 ( .A1(data_out_b[22]), .A2(n96), .B1(adder[22]), .B2(n5), .C1(
        n6), .C2(f[22]), .ZN(n53) );
  INV_X1 U86 ( .A(n53), .ZN(n182) );
  AOI222_X1 U87 ( .A1(data_out_b[21]), .A2(n96), .B1(adder[21]), .B2(n5), .C1(
        n6), .C2(f[21]), .ZN(n54) );
  INV_X1 U88 ( .A(n54), .ZN(n183) );
  INV_X1 U89 ( .A(n189), .ZN(n55) );
  AOI222_X1 U90 ( .A1(data_out_b[20]), .A2(n96), .B1(adder[20]), .B2(n5), .C1(
        n6), .C2(n55), .ZN(n56) );
  INV_X1 U91 ( .A(n56), .ZN(n184) );
  INV_X1 U92 ( .A(n190), .ZN(n57) );
  AOI222_X1 U93 ( .A1(data_out_b[19]), .A2(n96), .B1(adder[19]), .B2(n5), .C1(
        n6), .C2(n57), .ZN(n58) );
  INV_X1 U94 ( .A(n58), .ZN(n185) );
  INV_X1 U95 ( .A(n191), .ZN(n59) );
  AOI222_X1 U96 ( .A1(data_out_b[18]), .A2(n96), .B1(adder[18]), .B2(n7), .C1(
        n95), .C2(n59), .ZN(n60) );
  INV_X1 U97 ( .A(n60), .ZN(n186) );
  INV_X1 U98 ( .A(n192), .ZN(n61) );
  AOI222_X1 U99 ( .A1(data_out_b[17]), .A2(n96), .B1(adder[17]), .B2(n7), .C1(
        n95), .C2(n61), .ZN(n62) );
  INV_X1 U100 ( .A(n62), .ZN(n187) );
  INV_X1 U101 ( .A(n193), .ZN(n63) );
  AOI222_X1 U102 ( .A1(data_out_b[16]), .A2(n96), .B1(adder[16]), .B2(n7), 
        .C1(n95), .C2(n63), .ZN(n64) );
  INV_X1 U103 ( .A(n64), .ZN(n188) );
  INV_X1 U104 ( .A(n194), .ZN(n65) );
  AOI222_X1 U105 ( .A1(data_out_b[15]), .A2(n96), .B1(adder[15]), .B2(n7), 
        .C1(n95), .C2(n65), .ZN(n66) );
  INV_X1 U106 ( .A(n66), .ZN(n274) );
  INV_X1 U107 ( .A(n195), .ZN(n67) );
  AOI222_X1 U108 ( .A1(data_out_b[14]), .A2(n96), .B1(adder[14]), .B2(n7), 
        .C1(n95), .C2(n67), .ZN(n68) );
  INV_X1 U109 ( .A(n68), .ZN(n275) );
  INV_X1 U110 ( .A(n196), .ZN(n69) );
  AOI222_X1 U111 ( .A1(data_out_b[13]), .A2(n96), .B1(adder[13]), .B2(n7), 
        .C1(n95), .C2(n69), .ZN(n70) );
  INV_X1 U112 ( .A(n70), .ZN(n276) );
  INV_X1 U113 ( .A(n197), .ZN(n71) );
  AOI222_X1 U114 ( .A1(data_out_b[12]), .A2(n96), .B1(adder[12]), .B2(n7), 
        .C1(n95), .C2(n71), .ZN(n72) );
  INV_X1 U115 ( .A(n72), .ZN(n277) );
  INV_X1 U116 ( .A(n198), .ZN(n73) );
  AOI222_X1 U117 ( .A1(data_out_b[11]), .A2(n96), .B1(adder[11]), .B2(n7), 
        .C1(n95), .C2(n73), .ZN(n74) );
  INV_X1 U118 ( .A(n74), .ZN(n278) );
  INV_X1 U119 ( .A(n199), .ZN(n75) );
  AOI222_X1 U120 ( .A1(data_out_b[10]), .A2(n8), .B1(adder[10]), .B2(n7), .C1(
        n95), .C2(n75), .ZN(n76) );
  INV_X1 U121 ( .A(n76), .ZN(n279) );
  AOI222_X1 U122 ( .A1(data_out_b[9]), .A2(n8), .B1(adder[9]), .B2(n7), .C1(
        n95), .C2(f[9]), .ZN(n77) );
  INV_X1 U123 ( .A(n77), .ZN(n280) );
  INV_X1 U124 ( .A(n201), .ZN(n78) );
  AOI222_X1 U125 ( .A1(data_out_b[8]), .A2(n8), .B1(adder[8]), .B2(n7), .C1(
        n95), .C2(n78), .ZN(n79) );
  INV_X1 U126 ( .A(n79), .ZN(n281) );
  INV_X1 U127 ( .A(n202), .ZN(n80) );
  AOI222_X1 U128 ( .A1(data_out_b[7]), .A2(n8), .B1(adder[7]), .B2(n7), .C1(
        n95), .C2(n80), .ZN(n81) );
  INV_X1 U129 ( .A(n81), .ZN(n282) );
  INV_X1 U130 ( .A(n203), .ZN(n82) );
  AOI222_X1 U131 ( .A1(data_out_b[6]), .A2(n8), .B1(adder[6]), .B2(n5), .C1(
        n95), .C2(n82), .ZN(n83) );
  INV_X1 U132 ( .A(n83), .ZN(n283) );
  INV_X1 U133 ( .A(n204), .ZN(n84) );
  AOI222_X1 U134 ( .A1(data_out_b[5]), .A2(n8), .B1(adder[5]), .B2(n5), .C1(
        n95), .C2(n84), .ZN(n85) );
  INV_X1 U135 ( .A(n85), .ZN(n284) );
  INV_X1 U136 ( .A(n205), .ZN(n86) );
  AOI222_X1 U137 ( .A1(data_out_b[4]), .A2(n8), .B1(adder[4]), .B2(n5), .C1(
        n95), .C2(n86), .ZN(n87) );
  INV_X1 U138 ( .A(n87), .ZN(n285) );
  AOI222_X1 U139 ( .A1(data_out_b[3]), .A2(n8), .B1(adder[3]), .B2(n5), .C1(
        n95), .C2(f[3]), .ZN(n88) );
  INV_X1 U140 ( .A(n88), .ZN(n286) );
  INV_X1 U141 ( .A(n207), .ZN(n89) );
  AOI222_X1 U142 ( .A1(data_out_b[2]), .A2(n8), .B1(adder[2]), .B2(n5), .C1(
        n95), .C2(n89), .ZN(n90) );
  INV_X1 U143 ( .A(n90), .ZN(n287) );
  INV_X1 U144 ( .A(n208), .ZN(n91) );
  AOI222_X1 U145 ( .A1(data_out_b[1]), .A2(n8), .B1(adder[1]), .B2(n5), .C1(
        n95), .C2(n91), .ZN(n92) );
  INV_X1 U146 ( .A(n92), .ZN(n288) );
  INV_X1 U147 ( .A(n209), .ZN(n93) );
  AOI222_X1 U148 ( .A1(data_out_b[0]), .A2(n8), .B1(adder[0]), .B2(n5), .C1(
        n95), .C2(n93), .ZN(n94) );
  INV_X1 U149 ( .A(n94), .ZN(n289) );
  AOI222_X1 U150 ( .A1(data_out_b[30]), .A2(n8), .B1(adder[30]), .B2(n5), .C1(
        n95), .C2(f[30]), .ZN(n97) );
  INV_X1 U151 ( .A(n97), .ZN(n141) );
  NOR4_X1 U152 ( .A1(f[11]), .A2(f[12]), .A3(f[13]), .A4(f[14]), .ZN(n132) );
  NOR4_X1 U153 ( .A1(f[7]), .A2(f[8]), .A3(f[9]), .A4(f[10]), .ZN(n127) );
  NAND4_X1 U154 ( .A1(n203), .A2(n204), .A3(n205), .A4(n206), .ZN(n98) );
  NOR4_X1 U155 ( .A1(n98), .A2(f[0]), .A3(f[1]), .A4(f[2]), .ZN(n126) );
  NAND4_X1 U156 ( .A1(n191), .A2(n192), .A3(n193), .A4(n194), .ZN(n116) );
  NAND4_X1 U157 ( .A1(n100), .A2(n99), .A3(n189), .A4(n190), .ZN(n115) );
  NAND4_X1 U158 ( .A1(n104), .A2(n103), .A3(n102), .A4(n101), .ZN(n110) );
  NAND4_X1 U159 ( .A1(n108), .A2(n107), .A3(n106), .A4(n105), .ZN(n109) );
  NOR4_X1 U160 ( .A1(n116), .A2(n115), .A3(n110), .A4(n109), .ZN(n125) );
  NAND4_X1 U161 ( .A1(n132), .A2(n127), .A3(n126), .A4(n125), .ZN(n135) );
  NAND3_X1 U162 ( .A1(wr_en_y), .A2(n135), .A3(n134), .ZN(n138) );
  INV_X1 U163 ( .A(wr_en_y), .ZN(n136) );
  NAND2_X1 U164 ( .A1(n139), .A2(n136), .ZN(n137) );
  OAI22_X1 U165 ( .A1(n209), .A2(n10), .B1(n241), .B2(n9), .ZN(n242) );
  OAI22_X1 U166 ( .A1(n208), .A2(n10), .B1(n240), .B2(n9), .ZN(n243) );
  OAI22_X1 U167 ( .A1(n207), .A2(n10), .B1(n239), .B2(n9), .ZN(n244) );
  OAI22_X1 U168 ( .A1(n206), .A2(n10), .B1(n238), .B2(n9), .ZN(n245) );
  OAI22_X1 U169 ( .A1(n205), .A2(n10), .B1(n237), .B2(n9), .ZN(n246) );
  OAI22_X1 U170 ( .A1(n204), .A2(n10), .B1(n236), .B2(n9), .ZN(n247) );
  OAI22_X1 U171 ( .A1(n203), .A2(n10), .B1(n235), .B2(n9), .ZN(n248) );
  OAI22_X1 U172 ( .A1(n202), .A2(n10), .B1(n234), .B2(n9), .ZN(n249) );
  OAI22_X1 U173 ( .A1(n201), .A2(n10), .B1(n233), .B2(n9), .ZN(n250) );
  OAI22_X1 U174 ( .A1(n200), .A2(n10), .B1(n232), .B2(n9), .ZN(n251) );
  OAI22_X1 U175 ( .A1(n199), .A2(n10), .B1(n231), .B2(n9), .ZN(n252) );
  OAI22_X1 U176 ( .A1(n198), .A2(n10), .B1(n230), .B2(n9), .ZN(n253) );
  OAI22_X1 U177 ( .A1(n197), .A2(n138), .B1(n229), .B2(n137), .ZN(n254) );
  OAI22_X1 U178 ( .A1(n196), .A2(n138), .B1(n228), .B2(n137), .ZN(n255) );
  OAI22_X1 U179 ( .A1(n195), .A2(n138), .B1(n227), .B2(n137), .ZN(n256) );
  OAI22_X1 U180 ( .A1(n194), .A2(n138), .B1(n226), .B2(n137), .ZN(n257) );
  OAI22_X1 U181 ( .A1(n193), .A2(n138), .B1(n225), .B2(n137), .ZN(n258) );
  OAI22_X1 U182 ( .A1(n192), .A2(n138), .B1(n224), .B2(n137), .ZN(n259) );
  OAI22_X1 U183 ( .A1(n191), .A2(n138), .B1(n223), .B2(n137), .ZN(n260) );
  OAI22_X1 U184 ( .A1(n190), .A2(n138), .B1(n222), .B2(n137), .ZN(n261) );
  OAI22_X1 U185 ( .A1(n189), .A2(n138), .B1(n221), .B2(n137), .ZN(n262) );
  OAI22_X1 U186 ( .A1(n99), .A2(n138), .B1(n220), .B2(n137), .ZN(n263) );
  OAI22_X1 U187 ( .A1(n100), .A2(n138), .B1(n219), .B2(n137), .ZN(n264) );
  OAI22_X1 U188 ( .A1(n101), .A2(n138), .B1(n218), .B2(n137), .ZN(n265) );
  OAI22_X1 U189 ( .A1(n102), .A2(n138), .B1(n217), .B2(n137), .ZN(n266) );
  OAI22_X1 U190 ( .A1(n103), .A2(n138), .B1(n216), .B2(n137), .ZN(n267) );
  OAI22_X1 U191 ( .A1(n104), .A2(n138), .B1(n215), .B2(n137), .ZN(n268) );
  OAI22_X1 U192 ( .A1(n105), .A2(n138), .B1(n214), .B2(n137), .ZN(n269) );
  OAI22_X1 U193 ( .A1(n106), .A2(n138), .B1(n213), .B2(n137), .ZN(n270) );
  OAI22_X1 U194 ( .A1(n107), .A2(n138), .B1(n212), .B2(n137), .ZN(n271) );
  OAI22_X1 U195 ( .A1(n108), .A2(n138), .B1(n211), .B2(n137), .ZN(n272) );
  OAI22_X1 U196 ( .A1(n134), .A2(n138), .B1(n210), .B2(n137), .ZN(n273) );
endmodule


module ctrlpath_M13_N16_T32_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HA_X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HA_X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INV_X1 U1 ( .A(A[0]), .ZN(SUM[0]) );
  XOR2_X1 U2 ( .A(carry[8]), .B(A[8]), .Z(SUM[8]) );
endmodule


module ctrlpath_M13_N16_T32 ( clk, reset, s_valid, s_ready, m_valid, m_ready, 
        clear_acc, wr_en_x, wr_en_y, addr_x, addr_w, addr_b );
  output [4:0] addr_x;
  output [7:0] addr_w;
  output [3:0] addr_b;
  input clk, reset, s_valid, m_ready;
  output s_ready, m_valid, clear_acc, wr_en_x, wr_en_y;
  wire   \addr_w2[8] , N11, N21, N22, N23, N24, clear_acc_delay, N75, N76, N77,
         N78, N79, N80, N81, N82, N83, N100, N103, n31, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, \add_158/carry[4] , \add_158/carry[3] , \add_158/carry[2] , n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n32,
         n43, n44, n45;
  wire   [3:0] state;
  wire   [3:0] out_count;

  DFF_X1 \addr_w2_reg[0]  ( .D(n8), .CK(clk), .Q(addr_w[0]) );
  DFF_X1 \addr_w2_reg[1]  ( .D(n9), .CK(clk), .Q(addr_w[1]) );
  DFF_X1 \addr_w2_reg[2]  ( .D(n10), .CK(clk), .Q(addr_w[2]) );
  DFF_X1 \addr_w2_reg[3]  ( .D(n11), .CK(clk), .Q(addr_w[3]) );
  DFF_X1 \addr_w2_reg[4]  ( .D(n12), .CK(clk), .Q(addr_w[4]) );
  DFF_X1 \addr_w2_reg[5]  ( .D(n13), .CK(clk), .Q(addr_w[5]) );
  DFF_X1 \addr_w2_reg[6]  ( .D(n14), .CK(clk), .Q(addr_w[6]) );
  DFF_X1 \addr_w2_reg[7]  ( .D(n15), .CK(clk), .Q(addr_w[7]) );
  OAI33_X1 U98 ( .A1(n47), .A2(n48), .A3(n49), .B1(n50), .B2(state[2]), .B3(
        reset), .ZN(s_ready) );
  NAND3_X1 U99 ( .A1(n53), .A2(n39), .A3(addr_b[1]), .ZN(n52) );
  NAND3_X1 U100 ( .A1(n62), .A2(n35), .A3(out_count[1]), .ZN(n66) );
  NAND3_X1 U101 ( .A1(n64), .A2(n44), .A3(n70), .ZN(n69) );
  NAND3_X1 U102 ( .A1(n80), .A2(n79), .A3(n48), .ZN(n92) );
  NAND3_X1 U103 ( .A1(state[2]), .A2(n29), .A3(state[1]), .ZN(n102) );
  NAND3_X1 U104 ( .A1(state[1]), .A2(state[2]), .A3(state[0]), .ZN(n70) );
  ctrlpath_M13_N16_T32_DW01_inc_0 add_193_S2 ( .A({\addr_w2[8] , addr_w}), 
        .SUM({N83, N82, N81, N80, N79, N78, N77, N76, N75}) );
  HA_X1 \add_158/U1_1_1  ( .A(addr_x[1]), .B(addr_x[0]), .CO(
        \add_158/carry[2] ), .S(N21) );
  HA_X1 \add_158/U1_1_2  ( .A(addr_x[2]), .B(\add_158/carry[2] ), .CO(
        \add_158/carry[3] ), .S(N22) );
  HA_X1 \add_158/U1_1_3  ( .A(addr_x[3]), .B(\add_158/carry[3] ), .CO(
        \add_158/carry[4] ), .S(N23) );
  DFF_X1 \state_reg[2]  ( .D(n4), .CK(clk), .Q(state[2]), .QN(n31) );
  DFF_X1 clear_acc_reg ( .D(N100), .CK(clk), .Q(clear_acc) );
  DFF_X1 clear_acc_delay_reg ( .D(N103), .CK(clk), .Q(clear_acc_delay) );
  DFF_X1 \state_reg[1]  ( .D(n7), .CK(clk), .Q(state[1]), .QN(n32) );
  DFF_X1 wr_en_y_reg ( .D(n2), .CK(clk), .Q(wr_en_y), .QN(n42) );
  DFF_X1 \addr_b_reg[0]  ( .D(n105), .CK(clk), .Q(addr_b[0]), .QN(n41) );
  DFF_X1 m_valid_reg ( .D(n111), .CK(clk), .Q(m_valid), .QN(n5) );
  DFF_X1 \addr_b_reg[1]  ( .D(n28), .CK(clk), .Q(addr_b[1]), .QN(n40) );
  DFF_X1 \addr_b_reg[2]  ( .D(n104), .CK(clk), .Q(addr_b[2]), .QN(n39) );
  DFF_X1 \out_count_reg[0]  ( .D(n109), .CK(clk), .Q(out_count[0]), .QN(n37)
         );
  DFF_X1 \addr_b_reg[3]  ( .D(n106), .CK(clk), .Q(addr_b[3]), .QN(n38) );
  DFF_X1 \out_count_reg[1]  ( .D(n25), .CK(clk), .Q(out_count[1]), .QN(n36) );
  DFF_X1 \out_count_reg[2]  ( .D(n108), .CK(clk), .Q(out_count[2]), .QN(n35)
         );
  DFF_X1 \out_count_reg[3]  ( .D(n107), .CK(clk), .Q(out_count[3]), .QN(n34)
         );
  DFF_X1 \state_reg[0]  ( .D(N11), .CK(clk), .Q(state[0]), .QN(n29) );
  DFF_X1 \addr_x_reg[4]  ( .D(n110), .CK(clk), .Q(addr_x[4]), .QN(n33) );
  DFF_X1 \addr_w2_reg[8]  ( .D(n16), .CK(clk), .Q(\addr_w2[8] ) );
  DFF_X1 \addr_x_reg[3]  ( .D(n21), .CK(clk), .Q(addr_x[3]) );
  DFF_X1 \addr_x_reg[1]  ( .D(n19), .CK(clk), .Q(addr_x[1]) );
  DFF_X1 \addr_x_reg[0]  ( .D(n18), .CK(clk), .Q(addr_x[0]), .QN(n6) );
  DFF_X1 \addr_x_reg[2]  ( .D(n20), .CK(clk), .Q(addr_x[2]) );
  NOR4_X1 U3 ( .A1(n26), .A2(n30), .A3(n72), .A4(reset), .ZN(n73) );
  AND3_X1 U4 ( .A1(state[2]), .A2(state[0]), .A3(n32), .ZN(n2) );
  NOR2_X1 U5 ( .A1(reset), .A2(n3), .ZN(n4) );
  INV_X1 U6 ( .A(n49), .ZN(n3) );
  INV_X1 U7 ( .A(n47), .ZN(n7) );
  AND3_X1 U8 ( .A1(n92), .A2(n44), .A3(n93), .ZN(n82) );
  AOI21_X1 U9 ( .B1(n48), .B2(n94), .A(n30), .ZN(n93) );
  NAND2_X1 U10 ( .A1(n2), .A2(n44), .ZN(n64) );
  OAI21_X1 U11 ( .B1(n2), .B2(n22), .A(n44), .ZN(n47) );
  INV_X1 U12 ( .A(n70), .ZN(n30) );
  INV_X1 U13 ( .A(n98), .ZN(n26) );
  NAND2_X1 U14 ( .A1(n98), .A2(n44), .ZN(N100) );
  INV_X1 U15 ( .A(n76), .ZN(n18) );
  AOI22_X1 U16 ( .A1(n6), .A2(n72), .B1(addr_x[0]), .B2(n73), .ZN(n76) );
  NOR2_X1 U17 ( .A1(n78), .A2(reset), .ZN(n72) );
  AOI21_X1 U18 ( .B1(n79), .B2(n80), .A(wr_en_x), .ZN(n78) );
  NOR3_X1 U19 ( .A1(n32), .A2(state[2]), .A3(n29), .ZN(n94) );
  AOI21_X1 U20 ( .B1(addr_x[4]), .B2(n80), .A(n22), .ZN(n48) );
  NOR2_X1 U21 ( .A1(n92), .A2(reset), .ZN(n83) );
  NOR2_X1 U22 ( .A1(n31), .A2(n50), .ZN(n80) );
  NOR3_X1 U23 ( .A1(n45), .A2(n48), .A3(n49), .ZN(wr_en_x) );
  INV_X1 U24 ( .A(s_valid), .ZN(n45) );
  NAND2_X1 U25 ( .A1(clear_acc_delay), .A2(n44), .ZN(n57) );
  OAI211_X1 U26 ( .C1(n32), .C2(n29), .A(n57), .B(n44), .ZN(n56) );
  NOR2_X1 U27 ( .A1(n41), .A2(n57), .ZN(n53) );
  AOI21_X1 U28 ( .B1(n40), .B2(n43), .A(n55), .ZN(n51) );
  INV_X1 U29 ( .A(n57), .ZN(n43) );
  AOI21_X1 U30 ( .B1(n36), .B2(n24), .A(n67), .ZN(n65) );
  INV_X1 U31 ( .A(n64), .ZN(n24) );
  NOR2_X1 U32 ( .A1(n37), .A2(n64), .ZN(n62) );
  AOI21_X1 U33 ( .B1(n94), .B2(addr_x[4]), .A(n103), .ZN(n98) );
  NOR3_X1 U34 ( .A1(state[0]), .A2(state[2]), .A3(n32), .ZN(n103) );
  OAI21_X1 U35 ( .B1(addr_b[0]), .B2(n57), .A(n56), .ZN(n55) );
  OAI21_X1 U36 ( .B1(out_count[0]), .B2(n64), .A(n69), .ZN(n67) );
  OAI22_X1 U37 ( .A1(n41), .A2(n56), .B1(addr_b[0]), .B2(n57), .ZN(n105) );
  OAI22_X1 U38 ( .A1(n37), .A2(n69), .B1(out_count[0]), .B2(n64), .ZN(n109) );
  OR4_X1 U39 ( .A1(n26), .A2(n95), .A3(n96), .A4(n80), .ZN(n49) );
  AND4_X1 U40 ( .A1(out_count[3]), .A2(out_count[2]), .A3(n32), .A4(state[2]), 
        .ZN(n96) );
  AOI21_X1 U41 ( .B1(n42), .B2(n79), .A(reset), .ZN(n111) );
  NAND2_X1 U42 ( .A1(n32), .A2(n29), .ZN(n50) );
  OR2_X1 U43 ( .A1(n5), .A2(m_ready), .ZN(n79) );
  OAI21_X1 U44 ( .B1(n33), .B2(n17), .A(n77), .ZN(n110) );
  NAND2_X1 U45 ( .A1(N24), .A2(n72), .ZN(n77) );
  INV_X1 U46 ( .A(n73), .ZN(n17) );
  OAI21_X1 U47 ( .B1(n51), .B2(n39), .A(n52), .ZN(n104) );
  OAI21_X1 U48 ( .B1(n65), .B2(n35), .A(n66), .ZN(n108) );
  OAI21_X1 U49 ( .B1(n23), .B2(n34), .A(n61), .ZN(n107) );
  NAND4_X1 U50 ( .A1(out_count[1]), .A2(n62), .A3(out_count[2]), .A4(n34), 
        .ZN(n61) );
  INV_X1 U51 ( .A(n63), .ZN(n23) );
  OAI21_X1 U52 ( .B1(n64), .B2(out_count[2]), .A(n65), .ZN(n63) );
  INV_X1 U53 ( .A(n99), .ZN(n22) );
  AOI221_X1 U54 ( .B1(s_valid), .B2(n100), .C1(n33), .C2(n94), .A(n95), .ZN(
        n99) );
  NOR2_X1 U55 ( .A1(n50), .A2(state[2]), .ZN(n100) );
  NOR2_X1 U56 ( .A1(reset), .A2(n48), .ZN(N11) );
  OAI21_X1 U57 ( .B1(n27), .B2(n38), .A(n58), .ZN(n106) );
  NAND4_X1 U58 ( .A1(addr_b[2]), .A2(addr_b[1]), .A3(n53), .A4(n38), .ZN(n58)
         );
  INV_X1 U59 ( .A(n59), .ZN(n27) );
  OAI21_X1 U60 ( .B1(n57), .B2(addr_b[2]), .A(n51), .ZN(n59) );
  OAI21_X1 U61 ( .B1(n101), .B2(n70), .A(n102), .ZN(n95) );
  AND2_X1 U62 ( .A1(m_ready), .A2(m_valid), .ZN(n101) );
  INV_X1 U63 ( .A(n74), .ZN(n20) );
  AOI22_X1 U64 ( .A1(N22), .A2(n72), .B1(addr_x[2]), .B2(n73), .ZN(n74) );
  INV_X1 U65 ( .A(n71), .ZN(n21) );
  AOI22_X1 U66 ( .A1(N23), .A2(n72), .B1(addr_x[3]), .B2(n73), .ZN(n71) );
  INV_X1 U67 ( .A(n75), .ZN(n19) );
  AOI22_X1 U68 ( .A1(N21), .A2(n72), .B1(addr_x[1]), .B2(n73), .ZN(n75) );
  INV_X1 U69 ( .A(n91), .ZN(n8) );
  AOI22_X1 U70 ( .A1(addr_w[0]), .A2(n82), .B1(N75), .B2(n83), .ZN(n91) );
  INV_X1 U71 ( .A(n84), .ZN(n15) );
  AOI22_X1 U72 ( .A1(addr_w[7]), .A2(n82), .B1(N82), .B2(n83), .ZN(n84) );
  INV_X1 U73 ( .A(n87), .ZN(n12) );
  AOI22_X1 U74 ( .A1(addr_w[4]), .A2(n82), .B1(N79), .B2(n83), .ZN(n87) );
  INV_X1 U75 ( .A(n89), .ZN(n10) );
  AOI22_X1 U76 ( .A1(addr_w[2]), .A2(n82), .B1(N77), .B2(n83), .ZN(n89) );
  INV_X1 U77 ( .A(n88), .ZN(n11) );
  AOI22_X1 U78 ( .A1(addr_w[3]), .A2(n82), .B1(N78), .B2(n83), .ZN(n88) );
  INV_X1 U79 ( .A(n90), .ZN(n9) );
  AOI22_X1 U80 ( .A1(addr_w[1]), .A2(n82), .B1(N76), .B2(n83), .ZN(n90) );
  INV_X1 U81 ( .A(n85), .ZN(n14) );
  AOI22_X1 U82 ( .A1(addr_w[6]), .A2(n82), .B1(N81), .B2(n83), .ZN(n85) );
  INV_X1 U83 ( .A(n86), .ZN(n13) );
  AOI22_X1 U84 ( .A1(addr_w[5]), .A2(n82), .B1(N80), .B2(n83), .ZN(n86) );
  AND2_X1 U85 ( .A1(clear_acc), .A2(n80), .ZN(N103) );
  INV_X1 U86 ( .A(n81), .ZN(n16) );
  AOI22_X1 U87 ( .A1(\addr_w2[8] ), .A2(n82), .B1(N83), .B2(n83), .ZN(n81) );
  INV_X1 U88 ( .A(n54), .ZN(n28) );
  AOI22_X1 U89 ( .A1(n55), .A2(addr_b[1]), .B1(n40), .B2(n53), .ZN(n54) );
  INV_X1 U90 ( .A(n68), .ZN(n25) );
  AOI22_X1 U91 ( .A1(n67), .A2(out_count[1]), .B1(n36), .B2(n62), .ZN(n68) );
  INV_X1 U92 ( .A(reset), .ZN(n44) );
  XOR2_X1 U93 ( .A(\add_158/carry[4] ), .B(addr_x[4]), .Z(N24) );
endmodule


module layer_13_16_1_32 ( clk, reset, s_valid, m_ready, data_in, m_valid, 
        s_ready, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, s_valid, m_ready;
  output m_valid, s_ready;
  wire   clear_acc, wr_en_x, wr_en_y;
  wire   [4:0] addr_x;
  wire   [7:0] addr_w;
  wire   [3:0] addr_b;

  datapath_M13_N16_T32 d ( .clk(clk), .clear_acc(clear_acc), .data_in(data_in), 
        .data_out(data_out), .wr_en_x(wr_en_x), .wr_en_y(wr_en_y), .addr_x(
        addr_x), .addr_w(addr_w), .addr_b(addr_b), .m_valid(m_valid), 
        .m_ready(m_ready) );
  ctrlpath_M13_N16_T32 c ( .clk(clk), .reset(reset), .s_valid(s_valid), 
        .s_ready(s_ready), .m_valid(m_valid), .m_ready(m_ready), .clear_acc(
        clear_acc), .wr_en_x(wr_en_x), .wr_en_y(wr_en_y), .addr_x(addr_x), 
        .addr_w(addr_w), .addr_b(addr_b) );
endmodule

